// Generator : SpinalHDL v1.8.0    git head : 4e3563a282582b41f4eaafc503787757251d23ea
// Component : CellSARA
// Git hash  : aeab30821bf33dec846c2049cebcf2d24a28afa4

`timescale 1ns/1ps

module CellSARA (
  input      [15:0]   io_in_r_data_0_data,
  input               io_in_r_data_0_load_store,
  input               io_in_r_data_0_df_is_ws,
  input               io_in_r_data_0_stall,
  input      [15:0]   io_in_r_data_1_data,
  input               io_in_r_data_1_load_store,
  input               io_in_r_data_1_df_is_ws,
  input               io_in_r_data_1_stall,
  input      [15:0]   io_in_r_data_2_data,
  input               io_in_r_data_2_load_store,
  input               io_in_r_data_2_df_is_ws,
  input               io_in_r_data_2_stall,
  input      [15:0]   io_in_r_data_3_data,
  input               io_in_r_data_3_load_store,
  input               io_in_r_data_3_df_is_ws,
  input               io_in_r_data_3_stall,
  input      [15:0]   io_in_r_bypass_0_0_data,
  input               io_in_r_bypass_0_0_load_store,
  input               io_in_r_bypass_0_0_df_is_ws,
  input               io_in_r_bypass_0_0_stall,
  input      [15:0]   io_in_r_bypass_0_1_data,
  input               io_in_r_bypass_0_1_load_store,
  input               io_in_r_bypass_0_1_df_is_ws,
  input               io_in_r_bypass_0_1_stall,
  input      [15:0]   io_in_r_bypass_0_2_data,
  input               io_in_r_bypass_0_2_load_store,
  input               io_in_r_bypass_0_2_df_is_ws,
  input               io_in_r_bypass_0_2_stall,
  input      [15:0]   io_in_r_bypass_0_3_data,
  input               io_in_r_bypass_0_3_load_store,
  input               io_in_r_bypass_0_3_df_is_ws,
  input               io_in_r_bypass_0_3_stall,
  input      [15:0]   io_in_r_bypass_1_0_data,
  input               io_in_r_bypass_1_0_load_store,
  input               io_in_r_bypass_1_0_df_is_ws,
  input               io_in_r_bypass_1_0_stall,
  input      [15:0]   io_in_r_bypass_1_1_data,
  input               io_in_r_bypass_1_1_load_store,
  input               io_in_r_bypass_1_1_df_is_ws,
  input               io_in_r_bypass_1_1_stall,
  input      [15:0]   io_in_r_bypass_1_2_data,
  input               io_in_r_bypass_1_2_load_store,
  input               io_in_r_bypass_1_2_df_is_ws,
  input               io_in_r_bypass_1_2_stall,
  input      [15:0]   io_in_r_bypass_1_3_data,
  input               io_in_r_bypass_1_3_load_store,
  input               io_in_r_bypass_1_3_df_is_ws,
  input               io_in_r_bypass_1_3_stall,
  input      [15:0]   io_in_r_bypass_2_0_data,
  input               io_in_r_bypass_2_0_load_store,
  input               io_in_r_bypass_2_0_df_is_ws,
  input               io_in_r_bypass_2_0_stall,
  input      [15:0]   io_in_r_bypass_2_1_data,
  input               io_in_r_bypass_2_1_load_store,
  input               io_in_r_bypass_2_1_df_is_ws,
  input               io_in_r_bypass_2_1_stall,
  input      [15:0]   io_in_r_bypass_2_2_data,
  input               io_in_r_bypass_2_2_load_store,
  input               io_in_r_bypass_2_2_df_is_ws,
  input               io_in_r_bypass_2_2_stall,
  input      [15:0]   io_in_r_bypass_2_3_data,
  input               io_in_r_bypass_2_3_load_store,
  input               io_in_r_bypass_2_3_df_is_ws,
  input               io_in_r_bypass_2_3_stall,
  input      [15:0]   io_in_r_bypass_3_0_data,
  input               io_in_r_bypass_3_0_load_store,
  input               io_in_r_bypass_3_0_df_is_ws,
  input               io_in_r_bypass_3_0_stall,
  input      [15:0]   io_in_r_bypass_3_1_data,
  input               io_in_r_bypass_3_1_load_store,
  input               io_in_r_bypass_3_1_df_is_ws,
  input               io_in_r_bypass_3_1_stall,
  input      [15:0]   io_in_r_bypass_3_2_data,
  input               io_in_r_bypass_3_2_load_store,
  input               io_in_r_bypass_3_2_df_is_ws,
  input               io_in_r_bypass_3_2_stall,
  input      [15:0]   io_in_r_bypass_3_3_data,
  input               io_in_r_bypass_3_3_load_store,
  input               io_in_r_bypass_3_3_df_is_ws,
  input               io_in_r_bypass_3_3_stall,
  input      [15:0]   io_in_r_bypass_4_0_data,
  input               io_in_r_bypass_4_0_load_store,
  input               io_in_r_bypass_4_0_df_is_ws,
  input               io_in_r_bypass_4_0_stall,
  input      [15:0]   io_in_r_bypass_4_1_data,
  input               io_in_r_bypass_4_1_load_store,
  input               io_in_r_bypass_4_1_df_is_ws,
  input               io_in_r_bypass_4_1_stall,
  input      [15:0]   io_in_r_bypass_4_2_data,
  input               io_in_r_bypass_4_2_load_store,
  input               io_in_r_bypass_4_2_df_is_ws,
  input               io_in_r_bypass_4_2_stall,
  input      [15:0]   io_in_r_bypass_4_3_data,
  input               io_in_r_bypass_4_3_load_store,
  input               io_in_r_bypass_4_3_df_is_ws,
  input               io_in_r_bypass_4_3_stall,
  input      [15:0]   io_in_r_bypass_5_0_data,
  input               io_in_r_bypass_5_0_load_store,
  input               io_in_r_bypass_5_0_df_is_ws,
  input               io_in_r_bypass_5_0_stall,
  input      [15:0]   io_in_r_bypass_5_1_data,
  input               io_in_r_bypass_5_1_load_store,
  input               io_in_r_bypass_5_1_df_is_ws,
  input               io_in_r_bypass_5_1_stall,
  input      [15:0]   io_in_r_bypass_5_2_data,
  input               io_in_r_bypass_5_2_load_store,
  input               io_in_r_bypass_5_2_df_is_ws,
  input               io_in_r_bypass_5_2_stall,
  input      [15:0]   io_in_r_bypass_5_3_data,
  input               io_in_r_bypass_5_3_load_store,
  input               io_in_r_bypass_5_3_df_is_ws,
  input               io_in_r_bypass_5_3_stall,
  input      [15:0]   io_in_r_bypass_6_0_data,
  input               io_in_r_bypass_6_0_load_store,
  input               io_in_r_bypass_6_0_df_is_ws,
  input               io_in_r_bypass_6_0_stall,
  input      [15:0]   io_in_r_bypass_6_1_data,
  input               io_in_r_bypass_6_1_load_store,
  input               io_in_r_bypass_6_1_df_is_ws,
  input               io_in_r_bypass_6_1_stall,
  input      [15:0]   io_in_r_bypass_6_2_data,
  input               io_in_r_bypass_6_2_load_store,
  input               io_in_r_bypass_6_2_df_is_ws,
  input               io_in_r_bypass_6_2_stall,
  input      [15:0]   io_in_r_bypass_6_3_data,
  input               io_in_r_bypass_6_3_load_store,
  input               io_in_r_bypass_6_3_df_is_ws,
  input               io_in_r_bypass_6_3_stall,
  input      [15:0]   io_in_r_bypass_7_0_data,
  input               io_in_r_bypass_7_0_load_store,
  input               io_in_r_bypass_7_0_df_is_ws,
  input               io_in_r_bypass_7_0_stall,
  input      [15:0]   io_in_r_bypass_7_1_data,
  input               io_in_r_bypass_7_1_load_store,
  input               io_in_r_bypass_7_1_df_is_ws,
  input               io_in_r_bypass_7_1_stall,
  input      [15:0]   io_in_r_bypass_7_2_data,
  input               io_in_r_bypass_7_2_load_store,
  input               io_in_r_bypass_7_2_df_is_ws,
  input               io_in_r_bypass_7_2_stall,
  input      [15:0]   io_in_r_bypass_7_3_data,
  input               io_in_r_bypass_7_3_load_store,
  input               io_in_r_bypass_7_3_df_is_ws,
  input               io_in_r_bypass_7_3_stall,
  input      [15:0]   io_in_r_bypass_8_0_data,
  input               io_in_r_bypass_8_0_load_store,
  input               io_in_r_bypass_8_0_df_is_ws,
  input               io_in_r_bypass_8_0_stall,
  input      [15:0]   io_in_r_bypass_8_1_data,
  input               io_in_r_bypass_8_1_load_store,
  input               io_in_r_bypass_8_1_df_is_ws,
  input               io_in_r_bypass_8_1_stall,
  input      [15:0]   io_in_r_bypass_8_2_data,
  input               io_in_r_bypass_8_2_load_store,
  input               io_in_r_bypass_8_2_df_is_ws,
  input               io_in_r_bypass_8_2_stall,
  input      [15:0]   io_in_r_bypass_8_3_data,
  input               io_in_r_bypass_8_3_load_store,
  input               io_in_r_bypass_8_3_df_is_ws,
  input               io_in_r_bypass_8_3_stall,
  input      [15:0]   io_in_r_bypass_9_0_data,
  input               io_in_r_bypass_9_0_load_store,
  input               io_in_r_bypass_9_0_df_is_ws,
  input               io_in_r_bypass_9_0_stall,
  input      [15:0]   io_in_r_bypass_9_1_data,
  input               io_in_r_bypass_9_1_load_store,
  input               io_in_r_bypass_9_1_df_is_ws,
  input               io_in_r_bypass_9_1_stall,
  input      [15:0]   io_in_r_bypass_9_2_data,
  input               io_in_r_bypass_9_2_load_store,
  input               io_in_r_bypass_9_2_df_is_ws,
  input               io_in_r_bypass_9_2_stall,
  input      [15:0]   io_in_r_bypass_9_3_data,
  input               io_in_r_bypass_9_3_load_store,
  input               io_in_r_bypass_9_3_df_is_ws,
  input               io_in_r_bypass_9_3_stall,
  input      [15:0]   io_in_r_bypass_10_0_data,
  input               io_in_r_bypass_10_0_load_store,
  input               io_in_r_bypass_10_0_df_is_ws,
  input               io_in_r_bypass_10_0_stall,
  input      [15:0]   io_in_r_bypass_10_1_data,
  input               io_in_r_bypass_10_1_load_store,
  input               io_in_r_bypass_10_1_df_is_ws,
  input               io_in_r_bypass_10_1_stall,
  input      [15:0]   io_in_r_bypass_10_2_data,
  input               io_in_r_bypass_10_2_load_store,
  input               io_in_r_bypass_10_2_df_is_ws,
  input               io_in_r_bypass_10_2_stall,
  input      [15:0]   io_in_r_bypass_10_3_data,
  input               io_in_r_bypass_10_3_load_store,
  input               io_in_r_bypass_10_3_df_is_ws,
  input               io_in_r_bypass_10_3_stall,
  input      [15:0]   io_in_r_bypass_11_0_data,
  input               io_in_r_bypass_11_0_load_store,
  input               io_in_r_bypass_11_0_df_is_ws,
  input               io_in_r_bypass_11_0_stall,
  input      [15:0]   io_in_r_bypass_11_1_data,
  input               io_in_r_bypass_11_1_load_store,
  input               io_in_r_bypass_11_1_df_is_ws,
  input               io_in_r_bypass_11_1_stall,
  input      [15:0]   io_in_r_bypass_11_2_data,
  input               io_in_r_bypass_11_2_load_store,
  input               io_in_r_bypass_11_2_df_is_ws,
  input               io_in_r_bypass_11_2_stall,
  input      [15:0]   io_in_r_bypass_11_3_data,
  input               io_in_r_bypass_11_3_load_store,
  input               io_in_r_bypass_11_3_df_is_ws,
  input               io_in_r_bypass_11_3_stall,
  input      [15:0]   io_in_r_bypass_12_0_data,
  input               io_in_r_bypass_12_0_load_store,
  input               io_in_r_bypass_12_0_df_is_ws,
  input               io_in_r_bypass_12_0_stall,
  input      [15:0]   io_in_r_bypass_12_1_data,
  input               io_in_r_bypass_12_1_load_store,
  input               io_in_r_bypass_12_1_df_is_ws,
  input               io_in_r_bypass_12_1_stall,
  input      [15:0]   io_in_r_bypass_12_2_data,
  input               io_in_r_bypass_12_2_load_store,
  input               io_in_r_bypass_12_2_df_is_ws,
  input               io_in_r_bypass_12_2_stall,
  input      [15:0]   io_in_r_bypass_12_3_data,
  input               io_in_r_bypass_12_3_load_store,
  input               io_in_r_bypass_12_3_df_is_ws,
  input               io_in_r_bypass_12_3_stall,
  input      [15:0]   io_in_r_bypass_13_0_data,
  input               io_in_r_bypass_13_0_load_store,
  input               io_in_r_bypass_13_0_df_is_ws,
  input               io_in_r_bypass_13_0_stall,
  input      [15:0]   io_in_r_bypass_13_1_data,
  input               io_in_r_bypass_13_1_load_store,
  input               io_in_r_bypass_13_1_df_is_ws,
  input               io_in_r_bypass_13_1_stall,
  input      [15:0]   io_in_r_bypass_13_2_data,
  input               io_in_r_bypass_13_2_load_store,
  input               io_in_r_bypass_13_2_df_is_ws,
  input               io_in_r_bypass_13_2_stall,
  input      [15:0]   io_in_r_bypass_13_3_data,
  input               io_in_r_bypass_13_3_load_store,
  input               io_in_r_bypass_13_3_df_is_ws,
  input               io_in_r_bypass_13_3_stall,
  input      [15:0]   io_in_r_bypass_14_0_data,
  input               io_in_r_bypass_14_0_load_store,
  input               io_in_r_bypass_14_0_df_is_ws,
  input               io_in_r_bypass_14_0_stall,
  input      [15:0]   io_in_r_bypass_14_1_data,
  input               io_in_r_bypass_14_1_load_store,
  input               io_in_r_bypass_14_1_df_is_ws,
  input               io_in_r_bypass_14_1_stall,
  input      [15:0]   io_in_r_bypass_14_2_data,
  input               io_in_r_bypass_14_2_load_store,
  input               io_in_r_bypass_14_2_df_is_ws,
  input               io_in_r_bypass_14_2_stall,
  input      [15:0]   io_in_r_bypass_14_3_data,
  input               io_in_r_bypass_14_3_load_store,
  input               io_in_r_bypass_14_3_df_is_ws,
  input               io_in_r_bypass_14_3_stall,
  input      [15:0]   io_in_r_bypass_15_0_data,
  input               io_in_r_bypass_15_0_load_store,
  input               io_in_r_bypass_15_0_df_is_ws,
  input               io_in_r_bypass_15_0_stall,
  input      [15:0]   io_in_r_bypass_15_1_data,
  input               io_in_r_bypass_15_1_load_store,
  input               io_in_r_bypass_15_1_df_is_ws,
  input               io_in_r_bypass_15_1_stall,
  input      [15:0]   io_in_r_bypass_15_2_data,
  input               io_in_r_bypass_15_2_load_store,
  input               io_in_r_bypass_15_2_df_is_ws,
  input               io_in_r_bypass_15_2_stall,
  input      [15:0]   io_in_r_bypass_15_3_data,
  input               io_in_r_bypass_15_3_load_store,
  input               io_in_r_bypass_15_3_df_is_ws,
  input               io_in_r_bypass_15_3_stall,
  input      [15:0]   io_in_r_bypass_16_0_data,
  input               io_in_r_bypass_16_0_load_store,
  input               io_in_r_bypass_16_0_df_is_ws,
  input               io_in_r_bypass_16_0_stall,
  input      [15:0]   io_in_r_bypass_16_1_data,
  input               io_in_r_bypass_16_1_load_store,
  input               io_in_r_bypass_16_1_df_is_ws,
  input               io_in_r_bypass_16_1_stall,
  input      [15:0]   io_in_r_bypass_16_2_data,
  input               io_in_r_bypass_16_2_load_store,
  input               io_in_r_bypass_16_2_df_is_ws,
  input               io_in_r_bypass_16_2_stall,
  input      [15:0]   io_in_r_bypass_16_3_data,
  input               io_in_r_bypass_16_3_load_store,
  input               io_in_r_bypass_16_3_df_is_ws,
  input               io_in_r_bypass_16_3_stall,
  input      [15:0]   io_in_r_bypass_17_0_data,
  input               io_in_r_bypass_17_0_load_store,
  input               io_in_r_bypass_17_0_df_is_ws,
  input               io_in_r_bypass_17_0_stall,
  input      [15:0]   io_in_r_bypass_17_1_data,
  input               io_in_r_bypass_17_1_load_store,
  input               io_in_r_bypass_17_1_df_is_ws,
  input               io_in_r_bypass_17_1_stall,
  input      [15:0]   io_in_r_bypass_17_2_data,
  input               io_in_r_bypass_17_2_load_store,
  input               io_in_r_bypass_17_2_df_is_ws,
  input               io_in_r_bypass_17_2_stall,
  input      [15:0]   io_in_r_bypass_17_3_data,
  input               io_in_r_bypass_17_3_load_store,
  input               io_in_r_bypass_17_3_df_is_ws,
  input               io_in_r_bypass_17_3_stall,
  input      [15:0]   io_in_r_bypass_18_0_data,
  input               io_in_r_bypass_18_0_load_store,
  input               io_in_r_bypass_18_0_df_is_ws,
  input               io_in_r_bypass_18_0_stall,
  input      [15:0]   io_in_r_bypass_18_1_data,
  input               io_in_r_bypass_18_1_load_store,
  input               io_in_r_bypass_18_1_df_is_ws,
  input               io_in_r_bypass_18_1_stall,
  input      [15:0]   io_in_r_bypass_18_2_data,
  input               io_in_r_bypass_18_2_load_store,
  input               io_in_r_bypass_18_2_df_is_ws,
  input               io_in_r_bypass_18_2_stall,
  input      [15:0]   io_in_r_bypass_18_3_data,
  input               io_in_r_bypass_18_3_load_store,
  input               io_in_r_bypass_18_3_df_is_ws,
  input               io_in_r_bypass_18_3_stall,
  input      [15:0]   io_in_r_bypass_19_0_data,
  input               io_in_r_bypass_19_0_load_store,
  input               io_in_r_bypass_19_0_df_is_ws,
  input               io_in_r_bypass_19_0_stall,
  input      [15:0]   io_in_r_bypass_19_1_data,
  input               io_in_r_bypass_19_1_load_store,
  input               io_in_r_bypass_19_1_df_is_ws,
  input               io_in_r_bypass_19_1_stall,
  input      [15:0]   io_in_r_bypass_19_2_data,
  input               io_in_r_bypass_19_2_load_store,
  input               io_in_r_bypass_19_2_df_is_ws,
  input               io_in_r_bypass_19_2_stall,
  input      [15:0]   io_in_r_bypass_19_3_data,
  input               io_in_r_bypass_19_3_load_store,
  input               io_in_r_bypass_19_3_df_is_ws,
  input               io_in_r_bypass_19_3_stall,
  input      [15:0]   io_in_r_bypass_20_0_data,
  input               io_in_r_bypass_20_0_load_store,
  input               io_in_r_bypass_20_0_df_is_ws,
  input               io_in_r_bypass_20_0_stall,
  input      [15:0]   io_in_r_bypass_20_1_data,
  input               io_in_r_bypass_20_1_load_store,
  input               io_in_r_bypass_20_1_df_is_ws,
  input               io_in_r_bypass_20_1_stall,
  input      [15:0]   io_in_r_bypass_20_2_data,
  input               io_in_r_bypass_20_2_load_store,
  input               io_in_r_bypass_20_2_df_is_ws,
  input               io_in_r_bypass_20_2_stall,
  input      [15:0]   io_in_r_bypass_20_3_data,
  input               io_in_r_bypass_20_3_load_store,
  input               io_in_r_bypass_20_3_df_is_ws,
  input               io_in_r_bypass_20_3_stall,
  input      [15:0]   io_in_r_bypass_21_0_data,
  input               io_in_r_bypass_21_0_load_store,
  input               io_in_r_bypass_21_0_df_is_ws,
  input               io_in_r_bypass_21_0_stall,
  input      [15:0]   io_in_r_bypass_21_1_data,
  input               io_in_r_bypass_21_1_load_store,
  input               io_in_r_bypass_21_1_df_is_ws,
  input               io_in_r_bypass_21_1_stall,
  input      [15:0]   io_in_r_bypass_21_2_data,
  input               io_in_r_bypass_21_2_load_store,
  input               io_in_r_bypass_21_2_df_is_ws,
  input               io_in_r_bypass_21_2_stall,
  input      [15:0]   io_in_r_bypass_21_3_data,
  input               io_in_r_bypass_21_3_load_store,
  input               io_in_r_bypass_21_3_df_is_ws,
  input               io_in_r_bypass_21_3_stall,
  input      [15:0]   io_in_r_bypass_22_0_data,
  input               io_in_r_bypass_22_0_load_store,
  input               io_in_r_bypass_22_0_df_is_ws,
  input               io_in_r_bypass_22_0_stall,
  input      [15:0]   io_in_r_bypass_22_1_data,
  input               io_in_r_bypass_22_1_load_store,
  input               io_in_r_bypass_22_1_df_is_ws,
  input               io_in_r_bypass_22_1_stall,
  input      [15:0]   io_in_r_bypass_22_2_data,
  input               io_in_r_bypass_22_2_load_store,
  input               io_in_r_bypass_22_2_df_is_ws,
  input               io_in_r_bypass_22_2_stall,
  input      [15:0]   io_in_r_bypass_22_3_data,
  input               io_in_r_bypass_22_3_load_store,
  input               io_in_r_bypass_22_3_df_is_ws,
  input               io_in_r_bypass_22_3_stall,
  input      [15:0]   io_in_r_bypass_23_0_data,
  input               io_in_r_bypass_23_0_load_store,
  input               io_in_r_bypass_23_0_df_is_ws,
  input               io_in_r_bypass_23_0_stall,
  input      [15:0]   io_in_r_bypass_23_1_data,
  input               io_in_r_bypass_23_1_load_store,
  input               io_in_r_bypass_23_1_df_is_ws,
  input               io_in_r_bypass_23_1_stall,
  input      [15:0]   io_in_r_bypass_23_2_data,
  input               io_in_r_bypass_23_2_load_store,
  input               io_in_r_bypass_23_2_df_is_ws,
  input               io_in_r_bypass_23_2_stall,
  input      [15:0]   io_in_r_bypass_23_3_data,
  input               io_in_r_bypass_23_3_load_store,
  input               io_in_r_bypass_23_3_df_is_ws,
  input               io_in_r_bypass_23_3_stall,
  input      [15:0]   io_in_r_bypass_24_0_data,
  input               io_in_r_bypass_24_0_load_store,
  input               io_in_r_bypass_24_0_df_is_ws,
  input               io_in_r_bypass_24_0_stall,
  input      [15:0]   io_in_r_bypass_24_1_data,
  input               io_in_r_bypass_24_1_load_store,
  input               io_in_r_bypass_24_1_df_is_ws,
  input               io_in_r_bypass_24_1_stall,
  input      [15:0]   io_in_r_bypass_24_2_data,
  input               io_in_r_bypass_24_2_load_store,
  input               io_in_r_bypass_24_2_df_is_ws,
  input               io_in_r_bypass_24_2_stall,
  input      [15:0]   io_in_r_bypass_24_3_data,
  input               io_in_r_bypass_24_3_load_store,
  input               io_in_r_bypass_24_3_df_is_ws,
  input               io_in_r_bypass_24_3_stall,
  input      [15:0]   io_in_r_bypass_25_0_data,
  input               io_in_r_bypass_25_0_load_store,
  input               io_in_r_bypass_25_0_df_is_ws,
  input               io_in_r_bypass_25_0_stall,
  input      [15:0]   io_in_r_bypass_25_1_data,
  input               io_in_r_bypass_25_1_load_store,
  input               io_in_r_bypass_25_1_df_is_ws,
  input               io_in_r_bypass_25_1_stall,
  input      [15:0]   io_in_r_bypass_25_2_data,
  input               io_in_r_bypass_25_2_load_store,
  input               io_in_r_bypass_25_2_df_is_ws,
  input               io_in_r_bypass_25_2_stall,
  input      [15:0]   io_in_r_bypass_25_3_data,
  input               io_in_r_bypass_25_3_load_store,
  input               io_in_r_bypass_25_3_df_is_ws,
  input               io_in_r_bypass_25_3_stall,
  input      [15:0]   io_in_r_bypass_26_0_data,
  input               io_in_r_bypass_26_0_load_store,
  input               io_in_r_bypass_26_0_df_is_ws,
  input               io_in_r_bypass_26_0_stall,
  input      [15:0]   io_in_r_bypass_26_1_data,
  input               io_in_r_bypass_26_1_load_store,
  input               io_in_r_bypass_26_1_df_is_ws,
  input               io_in_r_bypass_26_1_stall,
  input      [15:0]   io_in_r_bypass_26_2_data,
  input               io_in_r_bypass_26_2_load_store,
  input               io_in_r_bypass_26_2_df_is_ws,
  input               io_in_r_bypass_26_2_stall,
  input      [15:0]   io_in_r_bypass_26_3_data,
  input               io_in_r_bypass_26_3_load_store,
  input               io_in_r_bypass_26_3_df_is_ws,
  input               io_in_r_bypass_26_3_stall,
  input      [15:0]   io_in_r_bypass_27_0_data,
  input               io_in_r_bypass_27_0_load_store,
  input               io_in_r_bypass_27_0_df_is_ws,
  input               io_in_r_bypass_27_0_stall,
  input      [15:0]   io_in_r_bypass_27_1_data,
  input               io_in_r_bypass_27_1_load_store,
  input               io_in_r_bypass_27_1_df_is_ws,
  input               io_in_r_bypass_27_1_stall,
  input      [15:0]   io_in_r_bypass_27_2_data,
  input               io_in_r_bypass_27_2_load_store,
  input               io_in_r_bypass_27_2_df_is_ws,
  input               io_in_r_bypass_27_2_stall,
  input      [15:0]   io_in_r_bypass_27_3_data,
  input               io_in_r_bypass_27_3_load_store,
  input               io_in_r_bypass_27_3_df_is_ws,
  input               io_in_r_bypass_27_3_stall,
  input      [15:0]   io_in_r_bypass_28_0_data,
  input               io_in_r_bypass_28_0_load_store,
  input               io_in_r_bypass_28_0_df_is_ws,
  input               io_in_r_bypass_28_0_stall,
  input      [15:0]   io_in_r_bypass_28_1_data,
  input               io_in_r_bypass_28_1_load_store,
  input               io_in_r_bypass_28_1_df_is_ws,
  input               io_in_r_bypass_28_1_stall,
  input      [15:0]   io_in_r_bypass_28_2_data,
  input               io_in_r_bypass_28_2_load_store,
  input               io_in_r_bypass_28_2_df_is_ws,
  input               io_in_r_bypass_28_2_stall,
  input      [15:0]   io_in_r_bypass_28_3_data,
  input               io_in_r_bypass_28_3_load_store,
  input               io_in_r_bypass_28_3_df_is_ws,
  input               io_in_r_bypass_28_3_stall,
  input      [15:0]   io_in_r_bypass_29_0_data,
  input               io_in_r_bypass_29_0_load_store,
  input               io_in_r_bypass_29_0_df_is_ws,
  input               io_in_r_bypass_29_0_stall,
  input      [15:0]   io_in_r_bypass_29_1_data,
  input               io_in_r_bypass_29_1_load_store,
  input               io_in_r_bypass_29_1_df_is_ws,
  input               io_in_r_bypass_29_1_stall,
  input      [15:0]   io_in_r_bypass_29_2_data,
  input               io_in_r_bypass_29_2_load_store,
  input               io_in_r_bypass_29_2_df_is_ws,
  input               io_in_r_bypass_29_2_stall,
  input      [15:0]   io_in_r_bypass_29_3_data,
  input               io_in_r_bypass_29_3_load_store,
  input               io_in_r_bypass_29_3_df_is_ws,
  input               io_in_r_bypass_29_3_stall,
  input      [15:0]   io_in_r_bypass_30_0_data,
  input               io_in_r_bypass_30_0_load_store,
  input               io_in_r_bypass_30_0_df_is_ws,
  input               io_in_r_bypass_30_0_stall,
  input      [15:0]   io_in_r_bypass_30_1_data,
  input               io_in_r_bypass_30_1_load_store,
  input               io_in_r_bypass_30_1_df_is_ws,
  input               io_in_r_bypass_30_1_stall,
  input      [15:0]   io_in_r_bypass_30_2_data,
  input               io_in_r_bypass_30_2_load_store,
  input               io_in_r_bypass_30_2_df_is_ws,
  input               io_in_r_bypass_30_2_stall,
  input      [15:0]   io_in_r_bypass_30_3_data,
  input               io_in_r_bypass_30_3_load_store,
  input               io_in_r_bypass_30_3_df_is_ws,
  input               io_in_r_bypass_30_3_stall,
  input      [15:0]   io_in_r_bypass_31_0_data,
  input               io_in_r_bypass_31_0_load_store,
  input               io_in_r_bypass_31_0_df_is_ws,
  input               io_in_r_bypass_31_0_stall,
  input      [15:0]   io_in_r_bypass_31_1_data,
  input               io_in_r_bypass_31_1_load_store,
  input               io_in_r_bypass_31_1_df_is_ws,
  input               io_in_r_bypass_31_1_stall,
  input      [15:0]   io_in_r_bypass_31_2_data,
  input               io_in_r_bypass_31_2_load_store,
  input               io_in_r_bypass_31_2_df_is_ws,
  input               io_in_r_bypass_31_2_stall,
  input      [15:0]   io_in_r_bypass_31_3_data,
  input               io_in_r_bypass_31_3_load_store,
  input               io_in_r_bypass_31_3_df_is_ws,
  input               io_in_r_bypass_31_3_stall,
  input               io_in_r_input_from_bypass_0,
  input               io_in_r_input_from_bypass_1,
  input               io_in_r_input_from_bypass_2,
  input               io_in_r_input_from_bypass_3,
  input               io_in_r_input_from_bypass_4,
  input               io_in_r_input_from_bypass_5,
  input               io_in_r_input_from_bypass_6,
  input               io_in_r_input_from_bypass_7,
  input               io_in_r_input_from_bypass_8,
  input               io_in_r_input_from_bypass_9,
  input               io_in_r_input_from_bypass_10,
  input               io_in_r_input_from_bypass_11,
  input               io_in_r_input_from_bypass_12,
  input               io_in_r_input_from_bypass_13,
  input               io_in_r_input_from_bypass_14,
  input               io_in_r_input_from_bypass_15,
  input               io_in_r_input_from_bypass_16,
  input               io_in_r_input_from_bypass_17,
  input               io_in_r_input_from_bypass_18,
  input               io_in_r_input_from_bypass_19,
  input               io_in_r_input_from_bypass_20,
  input               io_in_r_input_from_bypass_21,
  input               io_in_r_input_from_bypass_22,
  input               io_in_r_input_from_bypass_23,
  input               io_in_r_input_from_bypass_24,
  input               io_in_r_input_from_bypass_25,
  input               io_in_r_input_from_bypass_26,
  input               io_in_r_input_from_bypass_27,
  input               io_in_r_input_from_bypass_28,
  input               io_in_r_input_from_bypass_29,
  input               io_in_r_input_from_bypass_30,
  input               io_in_r_input_from_bypass_31,
  output     [15:0]   io_out_r_data_0_data,
  output              io_out_r_data_0_load_store,
  output              io_out_r_data_0_df_is_ws,
  output              io_out_r_data_0_stall,
  output     [15:0]   io_out_r_data_1_data,
  output              io_out_r_data_1_load_store,
  output              io_out_r_data_1_df_is_ws,
  output              io_out_r_data_1_stall,
  output     [15:0]   io_out_r_data_2_data,
  output              io_out_r_data_2_load_store,
  output              io_out_r_data_2_df_is_ws,
  output              io_out_r_data_2_stall,
  output     [15:0]   io_out_r_data_3_data,
  output              io_out_r_data_3_load_store,
  output              io_out_r_data_3_df_is_ws,
  output              io_out_r_data_3_stall,
  output     [15:0]   io_out_r_bypass_0_0_data,
  output              io_out_r_bypass_0_0_load_store,
  output              io_out_r_bypass_0_0_df_is_ws,
  output              io_out_r_bypass_0_0_stall,
  output     [15:0]   io_out_r_bypass_0_1_data,
  output              io_out_r_bypass_0_1_load_store,
  output              io_out_r_bypass_0_1_df_is_ws,
  output              io_out_r_bypass_0_1_stall,
  output     [15:0]   io_out_r_bypass_0_2_data,
  output              io_out_r_bypass_0_2_load_store,
  output              io_out_r_bypass_0_2_df_is_ws,
  output              io_out_r_bypass_0_2_stall,
  output     [15:0]   io_out_r_bypass_0_3_data,
  output              io_out_r_bypass_0_3_load_store,
  output              io_out_r_bypass_0_3_df_is_ws,
  output              io_out_r_bypass_0_3_stall,
  output     [15:0]   io_out_r_bypass_1_0_data,
  output              io_out_r_bypass_1_0_load_store,
  output              io_out_r_bypass_1_0_df_is_ws,
  output              io_out_r_bypass_1_0_stall,
  output     [15:0]   io_out_r_bypass_1_1_data,
  output              io_out_r_bypass_1_1_load_store,
  output              io_out_r_bypass_1_1_df_is_ws,
  output              io_out_r_bypass_1_1_stall,
  output     [15:0]   io_out_r_bypass_1_2_data,
  output              io_out_r_bypass_1_2_load_store,
  output              io_out_r_bypass_1_2_df_is_ws,
  output              io_out_r_bypass_1_2_stall,
  output     [15:0]   io_out_r_bypass_1_3_data,
  output              io_out_r_bypass_1_3_load_store,
  output              io_out_r_bypass_1_3_df_is_ws,
  output              io_out_r_bypass_1_3_stall,
  output     [15:0]   io_out_r_bypass_2_0_data,
  output              io_out_r_bypass_2_0_load_store,
  output              io_out_r_bypass_2_0_df_is_ws,
  output              io_out_r_bypass_2_0_stall,
  output     [15:0]   io_out_r_bypass_2_1_data,
  output              io_out_r_bypass_2_1_load_store,
  output              io_out_r_bypass_2_1_df_is_ws,
  output              io_out_r_bypass_2_1_stall,
  output     [15:0]   io_out_r_bypass_2_2_data,
  output              io_out_r_bypass_2_2_load_store,
  output              io_out_r_bypass_2_2_df_is_ws,
  output              io_out_r_bypass_2_2_stall,
  output     [15:0]   io_out_r_bypass_2_3_data,
  output              io_out_r_bypass_2_3_load_store,
  output              io_out_r_bypass_2_3_df_is_ws,
  output              io_out_r_bypass_2_3_stall,
  output     [15:0]   io_out_r_bypass_3_0_data,
  output              io_out_r_bypass_3_0_load_store,
  output              io_out_r_bypass_3_0_df_is_ws,
  output              io_out_r_bypass_3_0_stall,
  output     [15:0]   io_out_r_bypass_3_1_data,
  output              io_out_r_bypass_3_1_load_store,
  output              io_out_r_bypass_3_1_df_is_ws,
  output              io_out_r_bypass_3_1_stall,
  output     [15:0]   io_out_r_bypass_3_2_data,
  output              io_out_r_bypass_3_2_load_store,
  output              io_out_r_bypass_3_2_df_is_ws,
  output              io_out_r_bypass_3_2_stall,
  output     [15:0]   io_out_r_bypass_3_3_data,
  output              io_out_r_bypass_3_3_load_store,
  output              io_out_r_bypass_3_3_df_is_ws,
  output              io_out_r_bypass_3_3_stall,
  output     [15:0]   io_out_r_bypass_4_0_data,
  output              io_out_r_bypass_4_0_load_store,
  output              io_out_r_bypass_4_0_df_is_ws,
  output              io_out_r_bypass_4_0_stall,
  output     [15:0]   io_out_r_bypass_4_1_data,
  output              io_out_r_bypass_4_1_load_store,
  output              io_out_r_bypass_4_1_df_is_ws,
  output              io_out_r_bypass_4_1_stall,
  output     [15:0]   io_out_r_bypass_4_2_data,
  output              io_out_r_bypass_4_2_load_store,
  output              io_out_r_bypass_4_2_df_is_ws,
  output              io_out_r_bypass_4_2_stall,
  output     [15:0]   io_out_r_bypass_4_3_data,
  output              io_out_r_bypass_4_3_load_store,
  output              io_out_r_bypass_4_3_df_is_ws,
  output              io_out_r_bypass_4_3_stall,
  output     [15:0]   io_out_r_bypass_5_0_data,
  output              io_out_r_bypass_5_0_load_store,
  output              io_out_r_bypass_5_0_df_is_ws,
  output              io_out_r_bypass_5_0_stall,
  output     [15:0]   io_out_r_bypass_5_1_data,
  output              io_out_r_bypass_5_1_load_store,
  output              io_out_r_bypass_5_1_df_is_ws,
  output              io_out_r_bypass_5_1_stall,
  output     [15:0]   io_out_r_bypass_5_2_data,
  output              io_out_r_bypass_5_2_load_store,
  output              io_out_r_bypass_5_2_df_is_ws,
  output              io_out_r_bypass_5_2_stall,
  output     [15:0]   io_out_r_bypass_5_3_data,
  output              io_out_r_bypass_5_3_load_store,
  output              io_out_r_bypass_5_3_df_is_ws,
  output              io_out_r_bypass_5_3_stall,
  output     [15:0]   io_out_r_bypass_6_0_data,
  output              io_out_r_bypass_6_0_load_store,
  output              io_out_r_bypass_6_0_df_is_ws,
  output              io_out_r_bypass_6_0_stall,
  output     [15:0]   io_out_r_bypass_6_1_data,
  output              io_out_r_bypass_6_1_load_store,
  output              io_out_r_bypass_6_1_df_is_ws,
  output              io_out_r_bypass_6_1_stall,
  output     [15:0]   io_out_r_bypass_6_2_data,
  output              io_out_r_bypass_6_2_load_store,
  output              io_out_r_bypass_6_2_df_is_ws,
  output              io_out_r_bypass_6_2_stall,
  output     [15:0]   io_out_r_bypass_6_3_data,
  output              io_out_r_bypass_6_3_load_store,
  output              io_out_r_bypass_6_3_df_is_ws,
  output              io_out_r_bypass_6_3_stall,
  output     [15:0]   io_out_r_bypass_7_0_data,
  output              io_out_r_bypass_7_0_load_store,
  output              io_out_r_bypass_7_0_df_is_ws,
  output              io_out_r_bypass_7_0_stall,
  output     [15:0]   io_out_r_bypass_7_1_data,
  output              io_out_r_bypass_7_1_load_store,
  output              io_out_r_bypass_7_1_df_is_ws,
  output              io_out_r_bypass_7_1_stall,
  output     [15:0]   io_out_r_bypass_7_2_data,
  output              io_out_r_bypass_7_2_load_store,
  output              io_out_r_bypass_7_2_df_is_ws,
  output              io_out_r_bypass_7_2_stall,
  output     [15:0]   io_out_r_bypass_7_3_data,
  output              io_out_r_bypass_7_3_load_store,
  output              io_out_r_bypass_7_3_df_is_ws,
  output              io_out_r_bypass_7_3_stall,
  output     [15:0]   io_out_r_bypass_8_0_data,
  output              io_out_r_bypass_8_0_load_store,
  output              io_out_r_bypass_8_0_df_is_ws,
  output              io_out_r_bypass_8_0_stall,
  output     [15:0]   io_out_r_bypass_8_1_data,
  output              io_out_r_bypass_8_1_load_store,
  output              io_out_r_bypass_8_1_df_is_ws,
  output              io_out_r_bypass_8_1_stall,
  output     [15:0]   io_out_r_bypass_8_2_data,
  output              io_out_r_bypass_8_2_load_store,
  output              io_out_r_bypass_8_2_df_is_ws,
  output              io_out_r_bypass_8_2_stall,
  output     [15:0]   io_out_r_bypass_8_3_data,
  output              io_out_r_bypass_8_3_load_store,
  output              io_out_r_bypass_8_3_df_is_ws,
  output              io_out_r_bypass_8_3_stall,
  output     [15:0]   io_out_r_bypass_9_0_data,
  output              io_out_r_bypass_9_0_load_store,
  output              io_out_r_bypass_9_0_df_is_ws,
  output              io_out_r_bypass_9_0_stall,
  output     [15:0]   io_out_r_bypass_9_1_data,
  output              io_out_r_bypass_9_1_load_store,
  output              io_out_r_bypass_9_1_df_is_ws,
  output              io_out_r_bypass_9_1_stall,
  output     [15:0]   io_out_r_bypass_9_2_data,
  output              io_out_r_bypass_9_2_load_store,
  output              io_out_r_bypass_9_2_df_is_ws,
  output              io_out_r_bypass_9_2_stall,
  output     [15:0]   io_out_r_bypass_9_3_data,
  output              io_out_r_bypass_9_3_load_store,
  output              io_out_r_bypass_9_3_df_is_ws,
  output              io_out_r_bypass_9_3_stall,
  output     [15:0]   io_out_r_bypass_10_0_data,
  output              io_out_r_bypass_10_0_load_store,
  output              io_out_r_bypass_10_0_df_is_ws,
  output              io_out_r_bypass_10_0_stall,
  output     [15:0]   io_out_r_bypass_10_1_data,
  output              io_out_r_bypass_10_1_load_store,
  output              io_out_r_bypass_10_1_df_is_ws,
  output              io_out_r_bypass_10_1_stall,
  output     [15:0]   io_out_r_bypass_10_2_data,
  output              io_out_r_bypass_10_2_load_store,
  output              io_out_r_bypass_10_2_df_is_ws,
  output              io_out_r_bypass_10_2_stall,
  output     [15:0]   io_out_r_bypass_10_3_data,
  output              io_out_r_bypass_10_3_load_store,
  output              io_out_r_bypass_10_3_df_is_ws,
  output              io_out_r_bypass_10_3_stall,
  output     [15:0]   io_out_r_bypass_11_0_data,
  output              io_out_r_bypass_11_0_load_store,
  output              io_out_r_bypass_11_0_df_is_ws,
  output              io_out_r_bypass_11_0_stall,
  output     [15:0]   io_out_r_bypass_11_1_data,
  output              io_out_r_bypass_11_1_load_store,
  output              io_out_r_bypass_11_1_df_is_ws,
  output              io_out_r_bypass_11_1_stall,
  output     [15:0]   io_out_r_bypass_11_2_data,
  output              io_out_r_bypass_11_2_load_store,
  output              io_out_r_bypass_11_2_df_is_ws,
  output              io_out_r_bypass_11_2_stall,
  output     [15:0]   io_out_r_bypass_11_3_data,
  output              io_out_r_bypass_11_3_load_store,
  output              io_out_r_bypass_11_3_df_is_ws,
  output              io_out_r_bypass_11_3_stall,
  output     [15:0]   io_out_r_bypass_12_0_data,
  output              io_out_r_bypass_12_0_load_store,
  output              io_out_r_bypass_12_0_df_is_ws,
  output              io_out_r_bypass_12_0_stall,
  output     [15:0]   io_out_r_bypass_12_1_data,
  output              io_out_r_bypass_12_1_load_store,
  output              io_out_r_bypass_12_1_df_is_ws,
  output              io_out_r_bypass_12_1_stall,
  output     [15:0]   io_out_r_bypass_12_2_data,
  output              io_out_r_bypass_12_2_load_store,
  output              io_out_r_bypass_12_2_df_is_ws,
  output              io_out_r_bypass_12_2_stall,
  output     [15:0]   io_out_r_bypass_12_3_data,
  output              io_out_r_bypass_12_3_load_store,
  output              io_out_r_bypass_12_3_df_is_ws,
  output              io_out_r_bypass_12_3_stall,
  output     [15:0]   io_out_r_bypass_13_0_data,
  output              io_out_r_bypass_13_0_load_store,
  output              io_out_r_bypass_13_0_df_is_ws,
  output              io_out_r_bypass_13_0_stall,
  output     [15:0]   io_out_r_bypass_13_1_data,
  output              io_out_r_bypass_13_1_load_store,
  output              io_out_r_bypass_13_1_df_is_ws,
  output              io_out_r_bypass_13_1_stall,
  output     [15:0]   io_out_r_bypass_13_2_data,
  output              io_out_r_bypass_13_2_load_store,
  output              io_out_r_bypass_13_2_df_is_ws,
  output              io_out_r_bypass_13_2_stall,
  output     [15:0]   io_out_r_bypass_13_3_data,
  output              io_out_r_bypass_13_3_load_store,
  output              io_out_r_bypass_13_3_df_is_ws,
  output              io_out_r_bypass_13_3_stall,
  output     [15:0]   io_out_r_bypass_14_0_data,
  output              io_out_r_bypass_14_0_load_store,
  output              io_out_r_bypass_14_0_df_is_ws,
  output              io_out_r_bypass_14_0_stall,
  output     [15:0]   io_out_r_bypass_14_1_data,
  output              io_out_r_bypass_14_1_load_store,
  output              io_out_r_bypass_14_1_df_is_ws,
  output              io_out_r_bypass_14_1_stall,
  output     [15:0]   io_out_r_bypass_14_2_data,
  output              io_out_r_bypass_14_2_load_store,
  output              io_out_r_bypass_14_2_df_is_ws,
  output              io_out_r_bypass_14_2_stall,
  output     [15:0]   io_out_r_bypass_14_3_data,
  output              io_out_r_bypass_14_3_load_store,
  output              io_out_r_bypass_14_3_df_is_ws,
  output              io_out_r_bypass_14_3_stall,
  output     [15:0]   io_out_r_bypass_15_0_data,
  output              io_out_r_bypass_15_0_load_store,
  output              io_out_r_bypass_15_0_df_is_ws,
  output              io_out_r_bypass_15_0_stall,
  output     [15:0]   io_out_r_bypass_15_1_data,
  output              io_out_r_bypass_15_1_load_store,
  output              io_out_r_bypass_15_1_df_is_ws,
  output              io_out_r_bypass_15_1_stall,
  output     [15:0]   io_out_r_bypass_15_2_data,
  output              io_out_r_bypass_15_2_load_store,
  output              io_out_r_bypass_15_2_df_is_ws,
  output              io_out_r_bypass_15_2_stall,
  output     [15:0]   io_out_r_bypass_15_3_data,
  output              io_out_r_bypass_15_3_load_store,
  output              io_out_r_bypass_15_3_df_is_ws,
  output              io_out_r_bypass_15_3_stall,
  output     [15:0]   io_out_r_bypass_16_0_data,
  output              io_out_r_bypass_16_0_load_store,
  output              io_out_r_bypass_16_0_df_is_ws,
  output              io_out_r_bypass_16_0_stall,
  output     [15:0]   io_out_r_bypass_16_1_data,
  output              io_out_r_bypass_16_1_load_store,
  output              io_out_r_bypass_16_1_df_is_ws,
  output              io_out_r_bypass_16_1_stall,
  output     [15:0]   io_out_r_bypass_16_2_data,
  output              io_out_r_bypass_16_2_load_store,
  output              io_out_r_bypass_16_2_df_is_ws,
  output              io_out_r_bypass_16_2_stall,
  output     [15:0]   io_out_r_bypass_16_3_data,
  output              io_out_r_bypass_16_3_load_store,
  output              io_out_r_bypass_16_3_df_is_ws,
  output              io_out_r_bypass_16_3_stall,
  output     [15:0]   io_out_r_bypass_17_0_data,
  output              io_out_r_bypass_17_0_load_store,
  output              io_out_r_bypass_17_0_df_is_ws,
  output              io_out_r_bypass_17_0_stall,
  output     [15:0]   io_out_r_bypass_17_1_data,
  output              io_out_r_bypass_17_1_load_store,
  output              io_out_r_bypass_17_1_df_is_ws,
  output              io_out_r_bypass_17_1_stall,
  output     [15:0]   io_out_r_bypass_17_2_data,
  output              io_out_r_bypass_17_2_load_store,
  output              io_out_r_bypass_17_2_df_is_ws,
  output              io_out_r_bypass_17_2_stall,
  output     [15:0]   io_out_r_bypass_17_3_data,
  output              io_out_r_bypass_17_3_load_store,
  output              io_out_r_bypass_17_3_df_is_ws,
  output              io_out_r_bypass_17_3_stall,
  output     [15:0]   io_out_r_bypass_18_0_data,
  output              io_out_r_bypass_18_0_load_store,
  output              io_out_r_bypass_18_0_df_is_ws,
  output              io_out_r_bypass_18_0_stall,
  output     [15:0]   io_out_r_bypass_18_1_data,
  output              io_out_r_bypass_18_1_load_store,
  output              io_out_r_bypass_18_1_df_is_ws,
  output              io_out_r_bypass_18_1_stall,
  output     [15:0]   io_out_r_bypass_18_2_data,
  output              io_out_r_bypass_18_2_load_store,
  output              io_out_r_bypass_18_2_df_is_ws,
  output              io_out_r_bypass_18_2_stall,
  output     [15:0]   io_out_r_bypass_18_3_data,
  output              io_out_r_bypass_18_3_load_store,
  output              io_out_r_bypass_18_3_df_is_ws,
  output              io_out_r_bypass_18_3_stall,
  output     [15:0]   io_out_r_bypass_19_0_data,
  output              io_out_r_bypass_19_0_load_store,
  output              io_out_r_bypass_19_0_df_is_ws,
  output              io_out_r_bypass_19_0_stall,
  output     [15:0]   io_out_r_bypass_19_1_data,
  output              io_out_r_bypass_19_1_load_store,
  output              io_out_r_bypass_19_1_df_is_ws,
  output              io_out_r_bypass_19_1_stall,
  output     [15:0]   io_out_r_bypass_19_2_data,
  output              io_out_r_bypass_19_2_load_store,
  output              io_out_r_bypass_19_2_df_is_ws,
  output              io_out_r_bypass_19_2_stall,
  output     [15:0]   io_out_r_bypass_19_3_data,
  output              io_out_r_bypass_19_3_load_store,
  output              io_out_r_bypass_19_3_df_is_ws,
  output              io_out_r_bypass_19_3_stall,
  output     [15:0]   io_out_r_bypass_20_0_data,
  output              io_out_r_bypass_20_0_load_store,
  output              io_out_r_bypass_20_0_df_is_ws,
  output              io_out_r_bypass_20_0_stall,
  output     [15:0]   io_out_r_bypass_20_1_data,
  output              io_out_r_bypass_20_1_load_store,
  output              io_out_r_bypass_20_1_df_is_ws,
  output              io_out_r_bypass_20_1_stall,
  output     [15:0]   io_out_r_bypass_20_2_data,
  output              io_out_r_bypass_20_2_load_store,
  output              io_out_r_bypass_20_2_df_is_ws,
  output              io_out_r_bypass_20_2_stall,
  output     [15:0]   io_out_r_bypass_20_3_data,
  output              io_out_r_bypass_20_3_load_store,
  output              io_out_r_bypass_20_3_df_is_ws,
  output              io_out_r_bypass_20_3_stall,
  output     [15:0]   io_out_r_bypass_21_0_data,
  output              io_out_r_bypass_21_0_load_store,
  output              io_out_r_bypass_21_0_df_is_ws,
  output              io_out_r_bypass_21_0_stall,
  output     [15:0]   io_out_r_bypass_21_1_data,
  output              io_out_r_bypass_21_1_load_store,
  output              io_out_r_bypass_21_1_df_is_ws,
  output              io_out_r_bypass_21_1_stall,
  output     [15:0]   io_out_r_bypass_21_2_data,
  output              io_out_r_bypass_21_2_load_store,
  output              io_out_r_bypass_21_2_df_is_ws,
  output              io_out_r_bypass_21_2_stall,
  output     [15:0]   io_out_r_bypass_21_3_data,
  output              io_out_r_bypass_21_3_load_store,
  output              io_out_r_bypass_21_3_df_is_ws,
  output              io_out_r_bypass_21_3_stall,
  output     [15:0]   io_out_r_bypass_22_0_data,
  output              io_out_r_bypass_22_0_load_store,
  output              io_out_r_bypass_22_0_df_is_ws,
  output              io_out_r_bypass_22_0_stall,
  output     [15:0]   io_out_r_bypass_22_1_data,
  output              io_out_r_bypass_22_1_load_store,
  output              io_out_r_bypass_22_1_df_is_ws,
  output              io_out_r_bypass_22_1_stall,
  output     [15:0]   io_out_r_bypass_22_2_data,
  output              io_out_r_bypass_22_2_load_store,
  output              io_out_r_bypass_22_2_df_is_ws,
  output              io_out_r_bypass_22_2_stall,
  output     [15:0]   io_out_r_bypass_22_3_data,
  output              io_out_r_bypass_22_3_load_store,
  output              io_out_r_bypass_22_3_df_is_ws,
  output              io_out_r_bypass_22_3_stall,
  output     [15:0]   io_out_r_bypass_23_0_data,
  output              io_out_r_bypass_23_0_load_store,
  output              io_out_r_bypass_23_0_df_is_ws,
  output              io_out_r_bypass_23_0_stall,
  output     [15:0]   io_out_r_bypass_23_1_data,
  output              io_out_r_bypass_23_1_load_store,
  output              io_out_r_bypass_23_1_df_is_ws,
  output              io_out_r_bypass_23_1_stall,
  output     [15:0]   io_out_r_bypass_23_2_data,
  output              io_out_r_bypass_23_2_load_store,
  output              io_out_r_bypass_23_2_df_is_ws,
  output              io_out_r_bypass_23_2_stall,
  output     [15:0]   io_out_r_bypass_23_3_data,
  output              io_out_r_bypass_23_3_load_store,
  output              io_out_r_bypass_23_3_df_is_ws,
  output              io_out_r_bypass_23_3_stall,
  output     [15:0]   io_out_r_bypass_24_0_data,
  output              io_out_r_bypass_24_0_load_store,
  output              io_out_r_bypass_24_0_df_is_ws,
  output              io_out_r_bypass_24_0_stall,
  output     [15:0]   io_out_r_bypass_24_1_data,
  output              io_out_r_bypass_24_1_load_store,
  output              io_out_r_bypass_24_1_df_is_ws,
  output              io_out_r_bypass_24_1_stall,
  output     [15:0]   io_out_r_bypass_24_2_data,
  output              io_out_r_bypass_24_2_load_store,
  output              io_out_r_bypass_24_2_df_is_ws,
  output              io_out_r_bypass_24_2_stall,
  output     [15:0]   io_out_r_bypass_24_3_data,
  output              io_out_r_bypass_24_3_load_store,
  output              io_out_r_bypass_24_3_df_is_ws,
  output              io_out_r_bypass_24_3_stall,
  output     [15:0]   io_out_r_bypass_25_0_data,
  output              io_out_r_bypass_25_0_load_store,
  output              io_out_r_bypass_25_0_df_is_ws,
  output              io_out_r_bypass_25_0_stall,
  output     [15:0]   io_out_r_bypass_25_1_data,
  output              io_out_r_bypass_25_1_load_store,
  output              io_out_r_bypass_25_1_df_is_ws,
  output              io_out_r_bypass_25_1_stall,
  output     [15:0]   io_out_r_bypass_25_2_data,
  output              io_out_r_bypass_25_2_load_store,
  output              io_out_r_bypass_25_2_df_is_ws,
  output              io_out_r_bypass_25_2_stall,
  output     [15:0]   io_out_r_bypass_25_3_data,
  output              io_out_r_bypass_25_3_load_store,
  output              io_out_r_bypass_25_3_df_is_ws,
  output              io_out_r_bypass_25_3_stall,
  output     [15:0]   io_out_r_bypass_26_0_data,
  output              io_out_r_bypass_26_0_load_store,
  output              io_out_r_bypass_26_0_df_is_ws,
  output              io_out_r_bypass_26_0_stall,
  output     [15:0]   io_out_r_bypass_26_1_data,
  output              io_out_r_bypass_26_1_load_store,
  output              io_out_r_bypass_26_1_df_is_ws,
  output              io_out_r_bypass_26_1_stall,
  output     [15:0]   io_out_r_bypass_26_2_data,
  output              io_out_r_bypass_26_2_load_store,
  output              io_out_r_bypass_26_2_df_is_ws,
  output              io_out_r_bypass_26_2_stall,
  output     [15:0]   io_out_r_bypass_26_3_data,
  output              io_out_r_bypass_26_3_load_store,
  output              io_out_r_bypass_26_3_df_is_ws,
  output              io_out_r_bypass_26_3_stall,
  output     [15:0]   io_out_r_bypass_27_0_data,
  output              io_out_r_bypass_27_0_load_store,
  output              io_out_r_bypass_27_0_df_is_ws,
  output              io_out_r_bypass_27_0_stall,
  output     [15:0]   io_out_r_bypass_27_1_data,
  output              io_out_r_bypass_27_1_load_store,
  output              io_out_r_bypass_27_1_df_is_ws,
  output              io_out_r_bypass_27_1_stall,
  output     [15:0]   io_out_r_bypass_27_2_data,
  output              io_out_r_bypass_27_2_load_store,
  output              io_out_r_bypass_27_2_df_is_ws,
  output              io_out_r_bypass_27_2_stall,
  output     [15:0]   io_out_r_bypass_27_3_data,
  output              io_out_r_bypass_27_3_load_store,
  output              io_out_r_bypass_27_3_df_is_ws,
  output              io_out_r_bypass_27_3_stall,
  output     [15:0]   io_out_r_bypass_28_0_data,
  output              io_out_r_bypass_28_0_load_store,
  output              io_out_r_bypass_28_0_df_is_ws,
  output              io_out_r_bypass_28_0_stall,
  output     [15:0]   io_out_r_bypass_28_1_data,
  output              io_out_r_bypass_28_1_load_store,
  output              io_out_r_bypass_28_1_df_is_ws,
  output              io_out_r_bypass_28_1_stall,
  output     [15:0]   io_out_r_bypass_28_2_data,
  output              io_out_r_bypass_28_2_load_store,
  output              io_out_r_bypass_28_2_df_is_ws,
  output              io_out_r_bypass_28_2_stall,
  output     [15:0]   io_out_r_bypass_28_3_data,
  output              io_out_r_bypass_28_3_load_store,
  output              io_out_r_bypass_28_3_df_is_ws,
  output              io_out_r_bypass_28_3_stall,
  output     [15:0]   io_out_r_bypass_29_0_data,
  output              io_out_r_bypass_29_0_load_store,
  output              io_out_r_bypass_29_0_df_is_ws,
  output              io_out_r_bypass_29_0_stall,
  output     [15:0]   io_out_r_bypass_29_1_data,
  output              io_out_r_bypass_29_1_load_store,
  output              io_out_r_bypass_29_1_df_is_ws,
  output              io_out_r_bypass_29_1_stall,
  output     [15:0]   io_out_r_bypass_29_2_data,
  output              io_out_r_bypass_29_2_load_store,
  output              io_out_r_bypass_29_2_df_is_ws,
  output              io_out_r_bypass_29_2_stall,
  output     [15:0]   io_out_r_bypass_29_3_data,
  output              io_out_r_bypass_29_3_load_store,
  output              io_out_r_bypass_29_3_df_is_ws,
  output              io_out_r_bypass_29_3_stall,
  output     [15:0]   io_out_r_bypass_30_0_data,
  output              io_out_r_bypass_30_0_load_store,
  output              io_out_r_bypass_30_0_df_is_ws,
  output              io_out_r_bypass_30_0_stall,
  output     [15:0]   io_out_r_bypass_30_1_data,
  output              io_out_r_bypass_30_1_load_store,
  output              io_out_r_bypass_30_1_df_is_ws,
  output              io_out_r_bypass_30_1_stall,
  output     [15:0]   io_out_r_bypass_30_2_data,
  output              io_out_r_bypass_30_2_load_store,
  output              io_out_r_bypass_30_2_df_is_ws,
  output              io_out_r_bypass_30_2_stall,
  output     [15:0]   io_out_r_bypass_30_3_data,
  output              io_out_r_bypass_30_3_load_store,
  output              io_out_r_bypass_30_3_df_is_ws,
  output              io_out_r_bypass_30_3_stall,
  output     [15:0]   io_out_r_bypass_31_0_data,
  output              io_out_r_bypass_31_0_load_store,
  output              io_out_r_bypass_31_0_df_is_ws,
  output              io_out_r_bypass_31_0_stall,
  output     [15:0]   io_out_r_bypass_31_1_data,
  output              io_out_r_bypass_31_1_load_store,
  output              io_out_r_bypass_31_1_df_is_ws,
  output              io_out_r_bypass_31_1_stall,
  output     [15:0]   io_out_r_bypass_31_2_data,
  output              io_out_r_bypass_31_2_load_store,
  output              io_out_r_bypass_31_2_df_is_ws,
  output              io_out_r_bypass_31_2_stall,
  output     [15:0]   io_out_r_bypass_31_3_data,
  output              io_out_r_bypass_31_3_load_store,
  output              io_out_r_bypass_31_3_df_is_ws,
  output              io_out_r_bypass_31_3_stall,
  output              io_out_r_input_from_bypass_0,
  output              io_out_r_input_from_bypass_1,
  output              io_out_r_input_from_bypass_2,
  output              io_out_r_input_from_bypass_3,
  output              io_out_r_input_from_bypass_4,
  output              io_out_r_input_from_bypass_5,
  output              io_out_r_input_from_bypass_6,
  output              io_out_r_input_from_bypass_7,
  output              io_out_r_input_from_bypass_8,
  output              io_out_r_input_from_bypass_9,
  output              io_out_r_input_from_bypass_10,
  output              io_out_r_input_from_bypass_11,
  output              io_out_r_input_from_bypass_12,
  output              io_out_r_input_from_bypass_13,
  output              io_out_r_input_from_bypass_14,
  output              io_out_r_input_from_bypass_15,
  output              io_out_r_input_from_bypass_16,
  output              io_out_r_input_from_bypass_17,
  output              io_out_r_input_from_bypass_18,
  output              io_out_r_input_from_bypass_19,
  output              io_out_r_input_from_bypass_20,
  output              io_out_r_input_from_bypass_21,
  output              io_out_r_input_from_bypass_22,
  output              io_out_r_input_from_bypass_23,
  output              io_out_r_input_from_bypass_24,
  output              io_out_r_input_from_bypass_25,
  output              io_out_r_input_from_bypass_26,
  output              io_out_r_input_from_bypass_27,
  output              io_out_r_input_from_bypass_28,
  output              io_out_r_input_from_bypass_29,
  output              io_out_r_input_from_bypass_30,
  output              io_out_r_input_from_bypass_31,
  input      [15:0]   io_in_c_data_0_data,
  input               io_in_c_data_0_is_stationary,
  input      [15:0]   io_in_c_data_1_data,
  input               io_in_c_data_1_is_stationary,
  input      [15:0]   io_in_c_data_2_data,
  input               io_in_c_data_2_is_stationary,
  input      [15:0]   io_in_c_data_3_data,
  input               io_in_c_data_3_is_stationary,
  input      [15:0]   io_in_c_bypass_0_0_data,
  input               io_in_c_bypass_0_0_is_stationary,
  input      [15:0]   io_in_c_bypass_0_1_data,
  input               io_in_c_bypass_0_1_is_stationary,
  input      [15:0]   io_in_c_bypass_0_2_data,
  input               io_in_c_bypass_0_2_is_stationary,
  input      [15:0]   io_in_c_bypass_0_3_data,
  input               io_in_c_bypass_0_3_is_stationary,
  input      [15:0]   io_in_c_bypass_1_0_data,
  input               io_in_c_bypass_1_0_is_stationary,
  input      [15:0]   io_in_c_bypass_1_1_data,
  input               io_in_c_bypass_1_1_is_stationary,
  input      [15:0]   io_in_c_bypass_1_2_data,
  input               io_in_c_bypass_1_2_is_stationary,
  input      [15:0]   io_in_c_bypass_1_3_data,
  input               io_in_c_bypass_1_3_is_stationary,
  input      [15:0]   io_in_c_bypass_2_0_data,
  input               io_in_c_bypass_2_0_is_stationary,
  input      [15:0]   io_in_c_bypass_2_1_data,
  input               io_in_c_bypass_2_1_is_stationary,
  input      [15:0]   io_in_c_bypass_2_2_data,
  input               io_in_c_bypass_2_2_is_stationary,
  input      [15:0]   io_in_c_bypass_2_3_data,
  input               io_in_c_bypass_2_3_is_stationary,
  input      [15:0]   io_in_c_bypass_3_0_data,
  input               io_in_c_bypass_3_0_is_stationary,
  input      [15:0]   io_in_c_bypass_3_1_data,
  input               io_in_c_bypass_3_1_is_stationary,
  input      [15:0]   io_in_c_bypass_3_2_data,
  input               io_in_c_bypass_3_2_is_stationary,
  input      [15:0]   io_in_c_bypass_3_3_data,
  input               io_in_c_bypass_3_3_is_stationary,
  input      [15:0]   io_in_c_bypass_4_0_data,
  input               io_in_c_bypass_4_0_is_stationary,
  input      [15:0]   io_in_c_bypass_4_1_data,
  input               io_in_c_bypass_4_1_is_stationary,
  input      [15:0]   io_in_c_bypass_4_2_data,
  input               io_in_c_bypass_4_2_is_stationary,
  input      [15:0]   io_in_c_bypass_4_3_data,
  input               io_in_c_bypass_4_3_is_stationary,
  input      [15:0]   io_in_c_bypass_5_0_data,
  input               io_in_c_bypass_5_0_is_stationary,
  input      [15:0]   io_in_c_bypass_5_1_data,
  input               io_in_c_bypass_5_1_is_stationary,
  input      [15:0]   io_in_c_bypass_5_2_data,
  input               io_in_c_bypass_5_2_is_stationary,
  input      [15:0]   io_in_c_bypass_5_3_data,
  input               io_in_c_bypass_5_3_is_stationary,
  input      [15:0]   io_in_c_bypass_6_0_data,
  input               io_in_c_bypass_6_0_is_stationary,
  input      [15:0]   io_in_c_bypass_6_1_data,
  input               io_in_c_bypass_6_1_is_stationary,
  input      [15:0]   io_in_c_bypass_6_2_data,
  input               io_in_c_bypass_6_2_is_stationary,
  input      [15:0]   io_in_c_bypass_6_3_data,
  input               io_in_c_bypass_6_3_is_stationary,
  input      [15:0]   io_in_c_bypass_7_0_data,
  input               io_in_c_bypass_7_0_is_stationary,
  input      [15:0]   io_in_c_bypass_7_1_data,
  input               io_in_c_bypass_7_1_is_stationary,
  input      [15:0]   io_in_c_bypass_7_2_data,
  input               io_in_c_bypass_7_2_is_stationary,
  input      [15:0]   io_in_c_bypass_7_3_data,
  input               io_in_c_bypass_7_3_is_stationary,
  input      [15:0]   io_in_c_bypass_8_0_data,
  input               io_in_c_bypass_8_0_is_stationary,
  input      [15:0]   io_in_c_bypass_8_1_data,
  input               io_in_c_bypass_8_1_is_stationary,
  input      [15:0]   io_in_c_bypass_8_2_data,
  input               io_in_c_bypass_8_2_is_stationary,
  input      [15:0]   io_in_c_bypass_8_3_data,
  input               io_in_c_bypass_8_3_is_stationary,
  input      [15:0]   io_in_c_bypass_9_0_data,
  input               io_in_c_bypass_9_0_is_stationary,
  input      [15:0]   io_in_c_bypass_9_1_data,
  input               io_in_c_bypass_9_1_is_stationary,
  input      [15:0]   io_in_c_bypass_9_2_data,
  input               io_in_c_bypass_9_2_is_stationary,
  input      [15:0]   io_in_c_bypass_9_3_data,
  input               io_in_c_bypass_9_3_is_stationary,
  input      [15:0]   io_in_c_bypass_10_0_data,
  input               io_in_c_bypass_10_0_is_stationary,
  input      [15:0]   io_in_c_bypass_10_1_data,
  input               io_in_c_bypass_10_1_is_stationary,
  input      [15:0]   io_in_c_bypass_10_2_data,
  input               io_in_c_bypass_10_2_is_stationary,
  input      [15:0]   io_in_c_bypass_10_3_data,
  input               io_in_c_bypass_10_3_is_stationary,
  input      [15:0]   io_in_c_bypass_11_0_data,
  input               io_in_c_bypass_11_0_is_stationary,
  input      [15:0]   io_in_c_bypass_11_1_data,
  input               io_in_c_bypass_11_1_is_stationary,
  input      [15:0]   io_in_c_bypass_11_2_data,
  input               io_in_c_bypass_11_2_is_stationary,
  input      [15:0]   io_in_c_bypass_11_3_data,
  input               io_in_c_bypass_11_3_is_stationary,
  input      [15:0]   io_in_c_bypass_12_0_data,
  input               io_in_c_bypass_12_0_is_stationary,
  input      [15:0]   io_in_c_bypass_12_1_data,
  input               io_in_c_bypass_12_1_is_stationary,
  input      [15:0]   io_in_c_bypass_12_2_data,
  input               io_in_c_bypass_12_2_is_stationary,
  input      [15:0]   io_in_c_bypass_12_3_data,
  input               io_in_c_bypass_12_3_is_stationary,
  input      [15:0]   io_in_c_bypass_13_0_data,
  input               io_in_c_bypass_13_0_is_stationary,
  input      [15:0]   io_in_c_bypass_13_1_data,
  input               io_in_c_bypass_13_1_is_stationary,
  input      [15:0]   io_in_c_bypass_13_2_data,
  input               io_in_c_bypass_13_2_is_stationary,
  input      [15:0]   io_in_c_bypass_13_3_data,
  input               io_in_c_bypass_13_3_is_stationary,
  input      [15:0]   io_in_c_bypass_14_0_data,
  input               io_in_c_bypass_14_0_is_stationary,
  input      [15:0]   io_in_c_bypass_14_1_data,
  input               io_in_c_bypass_14_1_is_stationary,
  input      [15:0]   io_in_c_bypass_14_2_data,
  input               io_in_c_bypass_14_2_is_stationary,
  input      [15:0]   io_in_c_bypass_14_3_data,
  input               io_in_c_bypass_14_3_is_stationary,
  input      [15:0]   io_in_c_bypass_15_0_data,
  input               io_in_c_bypass_15_0_is_stationary,
  input      [15:0]   io_in_c_bypass_15_1_data,
  input               io_in_c_bypass_15_1_is_stationary,
  input      [15:0]   io_in_c_bypass_15_2_data,
  input               io_in_c_bypass_15_2_is_stationary,
  input      [15:0]   io_in_c_bypass_15_3_data,
  input               io_in_c_bypass_15_3_is_stationary,
  input      [15:0]   io_in_c_bypass_16_0_data,
  input               io_in_c_bypass_16_0_is_stationary,
  input      [15:0]   io_in_c_bypass_16_1_data,
  input               io_in_c_bypass_16_1_is_stationary,
  input      [15:0]   io_in_c_bypass_16_2_data,
  input               io_in_c_bypass_16_2_is_stationary,
  input      [15:0]   io_in_c_bypass_16_3_data,
  input               io_in_c_bypass_16_3_is_stationary,
  input      [15:0]   io_in_c_bypass_17_0_data,
  input               io_in_c_bypass_17_0_is_stationary,
  input      [15:0]   io_in_c_bypass_17_1_data,
  input               io_in_c_bypass_17_1_is_stationary,
  input      [15:0]   io_in_c_bypass_17_2_data,
  input               io_in_c_bypass_17_2_is_stationary,
  input      [15:0]   io_in_c_bypass_17_3_data,
  input               io_in_c_bypass_17_3_is_stationary,
  input      [15:0]   io_in_c_bypass_18_0_data,
  input               io_in_c_bypass_18_0_is_stationary,
  input      [15:0]   io_in_c_bypass_18_1_data,
  input               io_in_c_bypass_18_1_is_stationary,
  input      [15:0]   io_in_c_bypass_18_2_data,
  input               io_in_c_bypass_18_2_is_stationary,
  input      [15:0]   io_in_c_bypass_18_3_data,
  input               io_in_c_bypass_18_3_is_stationary,
  input      [15:0]   io_in_c_bypass_19_0_data,
  input               io_in_c_bypass_19_0_is_stationary,
  input      [15:0]   io_in_c_bypass_19_1_data,
  input               io_in_c_bypass_19_1_is_stationary,
  input      [15:0]   io_in_c_bypass_19_2_data,
  input               io_in_c_bypass_19_2_is_stationary,
  input      [15:0]   io_in_c_bypass_19_3_data,
  input               io_in_c_bypass_19_3_is_stationary,
  input      [15:0]   io_in_c_bypass_20_0_data,
  input               io_in_c_bypass_20_0_is_stationary,
  input      [15:0]   io_in_c_bypass_20_1_data,
  input               io_in_c_bypass_20_1_is_stationary,
  input      [15:0]   io_in_c_bypass_20_2_data,
  input               io_in_c_bypass_20_2_is_stationary,
  input      [15:0]   io_in_c_bypass_20_3_data,
  input               io_in_c_bypass_20_3_is_stationary,
  input      [15:0]   io_in_c_bypass_21_0_data,
  input               io_in_c_bypass_21_0_is_stationary,
  input      [15:0]   io_in_c_bypass_21_1_data,
  input               io_in_c_bypass_21_1_is_stationary,
  input      [15:0]   io_in_c_bypass_21_2_data,
  input               io_in_c_bypass_21_2_is_stationary,
  input      [15:0]   io_in_c_bypass_21_3_data,
  input               io_in_c_bypass_21_3_is_stationary,
  input      [15:0]   io_in_c_bypass_22_0_data,
  input               io_in_c_bypass_22_0_is_stationary,
  input      [15:0]   io_in_c_bypass_22_1_data,
  input               io_in_c_bypass_22_1_is_stationary,
  input      [15:0]   io_in_c_bypass_22_2_data,
  input               io_in_c_bypass_22_2_is_stationary,
  input      [15:0]   io_in_c_bypass_22_3_data,
  input               io_in_c_bypass_22_3_is_stationary,
  input      [15:0]   io_in_c_bypass_23_0_data,
  input               io_in_c_bypass_23_0_is_stationary,
  input      [15:0]   io_in_c_bypass_23_1_data,
  input               io_in_c_bypass_23_1_is_stationary,
  input      [15:0]   io_in_c_bypass_23_2_data,
  input               io_in_c_bypass_23_2_is_stationary,
  input      [15:0]   io_in_c_bypass_23_3_data,
  input               io_in_c_bypass_23_3_is_stationary,
  input      [15:0]   io_in_c_bypass_24_0_data,
  input               io_in_c_bypass_24_0_is_stationary,
  input      [15:0]   io_in_c_bypass_24_1_data,
  input               io_in_c_bypass_24_1_is_stationary,
  input      [15:0]   io_in_c_bypass_24_2_data,
  input               io_in_c_bypass_24_2_is_stationary,
  input      [15:0]   io_in_c_bypass_24_3_data,
  input               io_in_c_bypass_24_3_is_stationary,
  input      [15:0]   io_in_c_bypass_25_0_data,
  input               io_in_c_bypass_25_0_is_stationary,
  input      [15:0]   io_in_c_bypass_25_1_data,
  input               io_in_c_bypass_25_1_is_stationary,
  input      [15:0]   io_in_c_bypass_25_2_data,
  input               io_in_c_bypass_25_2_is_stationary,
  input      [15:0]   io_in_c_bypass_25_3_data,
  input               io_in_c_bypass_25_3_is_stationary,
  input      [15:0]   io_in_c_bypass_26_0_data,
  input               io_in_c_bypass_26_0_is_stationary,
  input      [15:0]   io_in_c_bypass_26_1_data,
  input               io_in_c_bypass_26_1_is_stationary,
  input      [15:0]   io_in_c_bypass_26_2_data,
  input               io_in_c_bypass_26_2_is_stationary,
  input      [15:0]   io_in_c_bypass_26_3_data,
  input               io_in_c_bypass_26_3_is_stationary,
  input      [15:0]   io_in_c_bypass_27_0_data,
  input               io_in_c_bypass_27_0_is_stationary,
  input      [15:0]   io_in_c_bypass_27_1_data,
  input               io_in_c_bypass_27_1_is_stationary,
  input      [15:0]   io_in_c_bypass_27_2_data,
  input               io_in_c_bypass_27_2_is_stationary,
  input      [15:0]   io_in_c_bypass_27_3_data,
  input               io_in_c_bypass_27_3_is_stationary,
  input      [15:0]   io_in_c_bypass_28_0_data,
  input               io_in_c_bypass_28_0_is_stationary,
  input      [15:0]   io_in_c_bypass_28_1_data,
  input               io_in_c_bypass_28_1_is_stationary,
  input      [15:0]   io_in_c_bypass_28_2_data,
  input               io_in_c_bypass_28_2_is_stationary,
  input      [15:0]   io_in_c_bypass_28_3_data,
  input               io_in_c_bypass_28_3_is_stationary,
  input      [15:0]   io_in_c_bypass_29_0_data,
  input               io_in_c_bypass_29_0_is_stationary,
  input      [15:0]   io_in_c_bypass_29_1_data,
  input               io_in_c_bypass_29_1_is_stationary,
  input      [15:0]   io_in_c_bypass_29_2_data,
  input               io_in_c_bypass_29_2_is_stationary,
  input      [15:0]   io_in_c_bypass_29_3_data,
  input               io_in_c_bypass_29_3_is_stationary,
  input      [15:0]   io_in_c_bypass_30_0_data,
  input               io_in_c_bypass_30_0_is_stationary,
  input      [15:0]   io_in_c_bypass_30_1_data,
  input               io_in_c_bypass_30_1_is_stationary,
  input      [15:0]   io_in_c_bypass_30_2_data,
  input               io_in_c_bypass_30_2_is_stationary,
  input      [15:0]   io_in_c_bypass_30_3_data,
  input               io_in_c_bypass_30_3_is_stationary,
  input      [15:0]   io_in_c_bypass_31_0_data,
  input               io_in_c_bypass_31_0_is_stationary,
  input      [15:0]   io_in_c_bypass_31_1_data,
  input               io_in_c_bypass_31_1_is_stationary,
  input      [15:0]   io_in_c_bypass_31_2_data,
  input               io_in_c_bypass_31_2_is_stationary,
  input      [15:0]   io_in_c_bypass_31_3_data,
  input               io_in_c_bypass_31_3_is_stationary,
  input               io_in_c_input_from_bypass_0,
  input               io_in_c_input_from_bypass_1,
  input               io_in_c_input_from_bypass_2,
  input               io_in_c_input_from_bypass_3,
  input               io_in_c_input_from_bypass_4,
  input               io_in_c_input_from_bypass_5,
  input               io_in_c_input_from_bypass_6,
  input               io_in_c_input_from_bypass_7,
  input               io_in_c_input_from_bypass_8,
  input               io_in_c_input_from_bypass_9,
  input               io_in_c_input_from_bypass_10,
  input               io_in_c_input_from_bypass_11,
  input               io_in_c_input_from_bypass_12,
  input               io_in_c_input_from_bypass_13,
  input               io_in_c_input_from_bypass_14,
  input               io_in_c_input_from_bypass_15,
  input               io_in_c_input_from_bypass_16,
  input               io_in_c_input_from_bypass_17,
  input               io_in_c_input_from_bypass_18,
  input               io_in_c_input_from_bypass_19,
  input               io_in_c_input_from_bypass_20,
  input               io_in_c_input_from_bypass_21,
  input               io_in_c_input_from_bypass_22,
  input               io_in_c_input_from_bypass_23,
  input               io_in_c_input_from_bypass_24,
  input               io_in_c_input_from_bypass_25,
  input               io_in_c_input_from_bypass_26,
  input               io_in_c_input_from_bypass_27,
  input               io_in_c_input_from_bypass_28,
  input               io_in_c_input_from_bypass_29,
  input               io_in_c_input_from_bypass_30,
  input               io_in_c_input_from_bypass_31,
  output     [15:0]   io_out_c_data_0_data,
  output              io_out_c_data_0_is_stationary,
  output     [15:0]   io_out_c_data_1_data,
  output              io_out_c_data_1_is_stationary,
  output     [15:0]   io_out_c_data_2_data,
  output              io_out_c_data_2_is_stationary,
  output     [15:0]   io_out_c_data_3_data,
  output              io_out_c_data_3_is_stationary,
  output     [15:0]   io_out_c_bypass_0_0_data,
  output              io_out_c_bypass_0_0_is_stationary,
  output     [15:0]   io_out_c_bypass_0_1_data,
  output              io_out_c_bypass_0_1_is_stationary,
  output     [15:0]   io_out_c_bypass_0_2_data,
  output              io_out_c_bypass_0_2_is_stationary,
  output     [15:0]   io_out_c_bypass_0_3_data,
  output              io_out_c_bypass_0_3_is_stationary,
  output     [15:0]   io_out_c_bypass_1_0_data,
  output              io_out_c_bypass_1_0_is_stationary,
  output     [15:0]   io_out_c_bypass_1_1_data,
  output              io_out_c_bypass_1_1_is_stationary,
  output     [15:0]   io_out_c_bypass_1_2_data,
  output              io_out_c_bypass_1_2_is_stationary,
  output     [15:0]   io_out_c_bypass_1_3_data,
  output              io_out_c_bypass_1_3_is_stationary,
  output     [15:0]   io_out_c_bypass_2_0_data,
  output              io_out_c_bypass_2_0_is_stationary,
  output     [15:0]   io_out_c_bypass_2_1_data,
  output              io_out_c_bypass_2_1_is_stationary,
  output     [15:0]   io_out_c_bypass_2_2_data,
  output              io_out_c_bypass_2_2_is_stationary,
  output     [15:0]   io_out_c_bypass_2_3_data,
  output              io_out_c_bypass_2_3_is_stationary,
  output     [15:0]   io_out_c_bypass_3_0_data,
  output              io_out_c_bypass_3_0_is_stationary,
  output     [15:0]   io_out_c_bypass_3_1_data,
  output              io_out_c_bypass_3_1_is_stationary,
  output     [15:0]   io_out_c_bypass_3_2_data,
  output              io_out_c_bypass_3_2_is_stationary,
  output     [15:0]   io_out_c_bypass_3_3_data,
  output              io_out_c_bypass_3_3_is_stationary,
  output     [15:0]   io_out_c_bypass_4_0_data,
  output              io_out_c_bypass_4_0_is_stationary,
  output     [15:0]   io_out_c_bypass_4_1_data,
  output              io_out_c_bypass_4_1_is_stationary,
  output     [15:0]   io_out_c_bypass_4_2_data,
  output              io_out_c_bypass_4_2_is_stationary,
  output     [15:0]   io_out_c_bypass_4_3_data,
  output              io_out_c_bypass_4_3_is_stationary,
  output     [15:0]   io_out_c_bypass_5_0_data,
  output              io_out_c_bypass_5_0_is_stationary,
  output     [15:0]   io_out_c_bypass_5_1_data,
  output              io_out_c_bypass_5_1_is_stationary,
  output     [15:0]   io_out_c_bypass_5_2_data,
  output              io_out_c_bypass_5_2_is_stationary,
  output     [15:0]   io_out_c_bypass_5_3_data,
  output              io_out_c_bypass_5_3_is_stationary,
  output     [15:0]   io_out_c_bypass_6_0_data,
  output              io_out_c_bypass_6_0_is_stationary,
  output     [15:0]   io_out_c_bypass_6_1_data,
  output              io_out_c_bypass_6_1_is_stationary,
  output     [15:0]   io_out_c_bypass_6_2_data,
  output              io_out_c_bypass_6_2_is_stationary,
  output     [15:0]   io_out_c_bypass_6_3_data,
  output              io_out_c_bypass_6_3_is_stationary,
  output     [15:0]   io_out_c_bypass_7_0_data,
  output              io_out_c_bypass_7_0_is_stationary,
  output     [15:0]   io_out_c_bypass_7_1_data,
  output              io_out_c_bypass_7_1_is_stationary,
  output     [15:0]   io_out_c_bypass_7_2_data,
  output              io_out_c_bypass_7_2_is_stationary,
  output     [15:0]   io_out_c_bypass_7_3_data,
  output              io_out_c_bypass_7_3_is_stationary,
  output     [15:0]   io_out_c_bypass_8_0_data,
  output              io_out_c_bypass_8_0_is_stationary,
  output     [15:0]   io_out_c_bypass_8_1_data,
  output              io_out_c_bypass_8_1_is_stationary,
  output     [15:0]   io_out_c_bypass_8_2_data,
  output              io_out_c_bypass_8_2_is_stationary,
  output     [15:0]   io_out_c_bypass_8_3_data,
  output              io_out_c_bypass_8_3_is_stationary,
  output     [15:0]   io_out_c_bypass_9_0_data,
  output              io_out_c_bypass_9_0_is_stationary,
  output     [15:0]   io_out_c_bypass_9_1_data,
  output              io_out_c_bypass_9_1_is_stationary,
  output     [15:0]   io_out_c_bypass_9_2_data,
  output              io_out_c_bypass_9_2_is_stationary,
  output     [15:0]   io_out_c_bypass_9_3_data,
  output              io_out_c_bypass_9_3_is_stationary,
  output     [15:0]   io_out_c_bypass_10_0_data,
  output              io_out_c_bypass_10_0_is_stationary,
  output     [15:0]   io_out_c_bypass_10_1_data,
  output              io_out_c_bypass_10_1_is_stationary,
  output     [15:0]   io_out_c_bypass_10_2_data,
  output              io_out_c_bypass_10_2_is_stationary,
  output     [15:0]   io_out_c_bypass_10_3_data,
  output              io_out_c_bypass_10_3_is_stationary,
  output     [15:0]   io_out_c_bypass_11_0_data,
  output              io_out_c_bypass_11_0_is_stationary,
  output     [15:0]   io_out_c_bypass_11_1_data,
  output              io_out_c_bypass_11_1_is_stationary,
  output     [15:0]   io_out_c_bypass_11_2_data,
  output              io_out_c_bypass_11_2_is_stationary,
  output     [15:0]   io_out_c_bypass_11_3_data,
  output              io_out_c_bypass_11_3_is_stationary,
  output     [15:0]   io_out_c_bypass_12_0_data,
  output              io_out_c_bypass_12_0_is_stationary,
  output     [15:0]   io_out_c_bypass_12_1_data,
  output              io_out_c_bypass_12_1_is_stationary,
  output     [15:0]   io_out_c_bypass_12_2_data,
  output              io_out_c_bypass_12_2_is_stationary,
  output     [15:0]   io_out_c_bypass_12_3_data,
  output              io_out_c_bypass_12_3_is_stationary,
  output     [15:0]   io_out_c_bypass_13_0_data,
  output              io_out_c_bypass_13_0_is_stationary,
  output     [15:0]   io_out_c_bypass_13_1_data,
  output              io_out_c_bypass_13_1_is_stationary,
  output     [15:0]   io_out_c_bypass_13_2_data,
  output              io_out_c_bypass_13_2_is_stationary,
  output     [15:0]   io_out_c_bypass_13_3_data,
  output              io_out_c_bypass_13_3_is_stationary,
  output     [15:0]   io_out_c_bypass_14_0_data,
  output              io_out_c_bypass_14_0_is_stationary,
  output     [15:0]   io_out_c_bypass_14_1_data,
  output              io_out_c_bypass_14_1_is_stationary,
  output     [15:0]   io_out_c_bypass_14_2_data,
  output              io_out_c_bypass_14_2_is_stationary,
  output     [15:0]   io_out_c_bypass_14_3_data,
  output              io_out_c_bypass_14_3_is_stationary,
  output     [15:0]   io_out_c_bypass_15_0_data,
  output              io_out_c_bypass_15_0_is_stationary,
  output     [15:0]   io_out_c_bypass_15_1_data,
  output              io_out_c_bypass_15_1_is_stationary,
  output     [15:0]   io_out_c_bypass_15_2_data,
  output              io_out_c_bypass_15_2_is_stationary,
  output     [15:0]   io_out_c_bypass_15_3_data,
  output              io_out_c_bypass_15_3_is_stationary,
  output     [15:0]   io_out_c_bypass_16_0_data,
  output              io_out_c_bypass_16_0_is_stationary,
  output     [15:0]   io_out_c_bypass_16_1_data,
  output              io_out_c_bypass_16_1_is_stationary,
  output     [15:0]   io_out_c_bypass_16_2_data,
  output              io_out_c_bypass_16_2_is_stationary,
  output     [15:0]   io_out_c_bypass_16_3_data,
  output              io_out_c_bypass_16_3_is_stationary,
  output     [15:0]   io_out_c_bypass_17_0_data,
  output              io_out_c_bypass_17_0_is_stationary,
  output     [15:0]   io_out_c_bypass_17_1_data,
  output              io_out_c_bypass_17_1_is_stationary,
  output     [15:0]   io_out_c_bypass_17_2_data,
  output              io_out_c_bypass_17_2_is_stationary,
  output     [15:0]   io_out_c_bypass_17_3_data,
  output              io_out_c_bypass_17_3_is_stationary,
  output     [15:0]   io_out_c_bypass_18_0_data,
  output              io_out_c_bypass_18_0_is_stationary,
  output     [15:0]   io_out_c_bypass_18_1_data,
  output              io_out_c_bypass_18_1_is_stationary,
  output     [15:0]   io_out_c_bypass_18_2_data,
  output              io_out_c_bypass_18_2_is_stationary,
  output     [15:0]   io_out_c_bypass_18_3_data,
  output              io_out_c_bypass_18_3_is_stationary,
  output     [15:0]   io_out_c_bypass_19_0_data,
  output              io_out_c_bypass_19_0_is_stationary,
  output     [15:0]   io_out_c_bypass_19_1_data,
  output              io_out_c_bypass_19_1_is_stationary,
  output     [15:0]   io_out_c_bypass_19_2_data,
  output              io_out_c_bypass_19_2_is_stationary,
  output     [15:0]   io_out_c_bypass_19_3_data,
  output              io_out_c_bypass_19_3_is_stationary,
  output     [15:0]   io_out_c_bypass_20_0_data,
  output              io_out_c_bypass_20_0_is_stationary,
  output     [15:0]   io_out_c_bypass_20_1_data,
  output              io_out_c_bypass_20_1_is_stationary,
  output     [15:0]   io_out_c_bypass_20_2_data,
  output              io_out_c_bypass_20_2_is_stationary,
  output     [15:0]   io_out_c_bypass_20_3_data,
  output              io_out_c_bypass_20_3_is_stationary,
  output     [15:0]   io_out_c_bypass_21_0_data,
  output              io_out_c_bypass_21_0_is_stationary,
  output     [15:0]   io_out_c_bypass_21_1_data,
  output              io_out_c_bypass_21_1_is_stationary,
  output     [15:0]   io_out_c_bypass_21_2_data,
  output              io_out_c_bypass_21_2_is_stationary,
  output     [15:0]   io_out_c_bypass_21_3_data,
  output              io_out_c_bypass_21_3_is_stationary,
  output     [15:0]   io_out_c_bypass_22_0_data,
  output              io_out_c_bypass_22_0_is_stationary,
  output     [15:0]   io_out_c_bypass_22_1_data,
  output              io_out_c_bypass_22_1_is_stationary,
  output     [15:0]   io_out_c_bypass_22_2_data,
  output              io_out_c_bypass_22_2_is_stationary,
  output     [15:0]   io_out_c_bypass_22_3_data,
  output              io_out_c_bypass_22_3_is_stationary,
  output     [15:0]   io_out_c_bypass_23_0_data,
  output              io_out_c_bypass_23_0_is_stationary,
  output     [15:0]   io_out_c_bypass_23_1_data,
  output              io_out_c_bypass_23_1_is_stationary,
  output     [15:0]   io_out_c_bypass_23_2_data,
  output              io_out_c_bypass_23_2_is_stationary,
  output     [15:0]   io_out_c_bypass_23_3_data,
  output              io_out_c_bypass_23_3_is_stationary,
  output     [15:0]   io_out_c_bypass_24_0_data,
  output              io_out_c_bypass_24_0_is_stationary,
  output     [15:0]   io_out_c_bypass_24_1_data,
  output              io_out_c_bypass_24_1_is_stationary,
  output     [15:0]   io_out_c_bypass_24_2_data,
  output              io_out_c_bypass_24_2_is_stationary,
  output     [15:0]   io_out_c_bypass_24_3_data,
  output              io_out_c_bypass_24_3_is_stationary,
  output     [15:0]   io_out_c_bypass_25_0_data,
  output              io_out_c_bypass_25_0_is_stationary,
  output     [15:0]   io_out_c_bypass_25_1_data,
  output              io_out_c_bypass_25_1_is_stationary,
  output     [15:0]   io_out_c_bypass_25_2_data,
  output              io_out_c_bypass_25_2_is_stationary,
  output     [15:0]   io_out_c_bypass_25_3_data,
  output              io_out_c_bypass_25_3_is_stationary,
  output     [15:0]   io_out_c_bypass_26_0_data,
  output              io_out_c_bypass_26_0_is_stationary,
  output     [15:0]   io_out_c_bypass_26_1_data,
  output              io_out_c_bypass_26_1_is_stationary,
  output     [15:0]   io_out_c_bypass_26_2_data,
  output              io_out_c_bypass_26_2_is_stationary,
  output     [15:0]   io_out_c_bypass_26_3_data,
  output              io_out_c_bypass_26_3_is_stationary,
  output     [15:0]   io_out_c_bypass_27_0_data,
  output              io_out_c_bypass_27_0_is_stationary,
  output     [15:0]   io_out_c_bypass_27_1_data,
  output              io_out_c_bypass_27_1_is_stationary,
  output     [15:0]   io_out_c_bypass_27_2_data,
  output              io_out_c_bypass_27_2_is_stationary,
  output     [15:0]   io_out_c_bypass_27_3_data,
  output              io_out_c_bypass_27_3_is_stationary,
  output     [15:0]   io_out_c_bypass_28_0_data,
  output              io_out_c_bypass_28_0_is_stationary,
  output     [15:0]   io_out_c_bypass_28_1_data,
  output              io_out_c_bypass_28_1_is_stationary,
  output     [15:0]   io_out_c_bypass_28_2_data,
  output              io_out_c_bypass_28_2_is_stationary,
  output     [15:0]   io_out_c_bypass_28_3_data,
  output              io_out_c_bypass_28_3_is_stationary,
  output     [15:0]   io_out_c_bypass_29_0_data,
  output              io_out_c_bypass_29_0_is_stationary,
  output     [15:0]   io_out_c_bypass_29_1_data,
  output              io_out_c_bypass_29_1_is_stationary,
  output     [15:0]   io_out_c_bypass_29_2_data,
  output              io_out_c_bypass_29_2_is_stationary,
  output     [15:0]   io_out_c_bypass_29_3_data,
  output              io_out_c_bypass_29_3_is_stationary,
  output     [15:0]   io_out_c_bypass_30_0_data,
  output              io_out_c_bypass_30_0_is_stationary,
  output     [15:0]   io_out_c_bypass_30_1_data,
  output              io_out_c_bypass_30_1_is_stationary,
  output     [15:0]   io_out_c_bypass_30_2_data,
  output              io_out_c_bypass_30_2_is_stationary,
  output     [15:0]   io_out_c_bypass_30_3_data,
  output              io_out_c_bypass_30_3_is_stationary,
  output     [15:0]   io_out_c_bypass_31_0_data,
  output              io_out_c_bypass_31_0_is_stationary,
  output     [15:0]   io_out_c_bypass_31_1_data,
  output              io_out_c_bypass_31_1_is_stationary,
  output     [15:0]   io_out_c_bypass_31_2_data,
  output              io_out_c_bypass_31_2_is_stationary,
  output     [15:0]   io_out_c_bypass_31_3_data,
  output              io_out_c_bypass_31_3_is_stationary,
  output              io_out_c_input_from_bypass_0,
  output              io_out_c_input_from_bypass_1,
  output              io_out_c_input_from_bypass_2,
  output              io_out_c_input_from_bypass_3,
  output              io_out_c_input_from_bypass_4,
  output              io_out_c_input_from_bypass_5,
  output              io_out_c_input_from_bypass_6,
  output              io_out_c_input_from_bypass_7,
  output              io_out_c_input_from_bypass_8,
  output              io_out_c_input_from_bypass_9,
  output              io_out_c_input_from_bypass_10,
  output              io_out_c_input_from_bypass_11,
  output              io_out_c_input_from_bypass_12,
  output              io_out_c_input_from_bypass_13,
  output              io_out_c_input_from_bypass_14,
  output              io_out_c_input_from_bypass_15,
  output              io_out_c_input_from_bypass_16,
  output              io_out_c_input_from_bypass_17,
  output              io_out_c_input_from_bypass_18,
  output              io_out_c_input_from_bypass_19,
  output              io_out_c_input_from_bypass_20,
  output              io_out_c_input_from_bypass_21,
  output              io_out_c_input_from_bypass_22,
  output              io_out_c_input_from_bypass_23,
  output              io_out_c_input_from_bypass_24,
  output              io_out_c_input_from_bypass_25,
  output              io_out_c_input_from_bypass_26,
  output              io_out_c_input_from_bypass_27,
  output              io_out_c_input_from_bypass_28,
  output              io_out_c_input_from_bypass_29,
  output              io_out_c_input_from_bypass_30,
  output              io_out_c_input_from_bypass_31,
  input               clk,
  input               reset
);

  wire       [15:0]   pes_0_0_io_out_r_data;
  wire                pes_0_0_io_out_r_load_store;
  wire                pes_0_0_io_out_r_df_is_ws;
  wire                pes_0_0_io_out_r_stall;
  wire       [15:0]   pes_0_0_io_out_c_data;
  wire                pes_0_0_io_out_c_is_stationary;
  wire       [15:0]   pes_0_1_io_out_r_data;
  wire                pes_0_1_io_out_r_load_store;
  wire                pes_0_1_io_out_r_df_is_ws;
  wire                pes_0_1_io_out_r_stall;
  wire       [15:0]   pes_0_1_io_out_c_data;
  wire                pes_0_1_io_out_c_is_stationary;
  wire       [15:0]   pes_0_2_io_out_r_data;
  wire                pes_0_2_io_out_r_load_store;
  wire                pes_0_2_io_out_r_df_is_ws;
  wire                pes_0_2_io_out_r_stall;
  wire       [15:0]   pes_0_2_io_out_c_data;
  wire                pes_0_2_io_out_c_is_stationary;
  wire       [15:0]   pes_0_3_io_out_r_data;
  wire                pes_0_3_io_out_r_load_store;
  wire                pes_0_3_io_out_r_df_is_ws;
  wire                pes_0_3_io_out_r_stall;
  wire       [15:0]   pes_0_3_io_out_c_data;
  wire                pes_0_3_io_out_c_is_stationary;
  wire       [15:0]   pes_1_0_io_out_r_data;
  wire                pes_1_0_io_out_r_load_store;
  wire                pes_1_0_io_out_r_df_is_ws;
  wire                pes_1_0_io_out_r_stall;
  wire       [15:0]   pes_1_0_io_out_c_data;
  wire                pes_1_0_io_out_c_is_stationary;
  wire       [15:0]   pes_1_1_io_out_r_data;
  wire                pes_1_1_io_out_r_load_store;
  wire                pes_1_1_io_out_r_df_is_ws;
  wire                pes_1_1_io_out_r_stall;
  wire       [15:0]   pes_1_1_io_out_c_data;
  wire                pes_1_1_io_out_c_is_stationary;
  wire       [15:0]   pes_1_2_io_out_r_data;
  wire                pes_1_2_io_out_r_load_store;
  wire                pes_1_2_io_out_r_df_is_ws;
  wire                pes_1_2_io_out_r_stall;
  wire       [15:0]   pes_1_2_io_out_c_data;
  wire                pes_1_2_io_out_c_is_stationary;
  wire       [15:0]   pes_1_3_io_out_r_data;
  wire                pes_1_3_io_out_r_load_store;
  wire                pes_1_3_io_out_r_df_is_ws;
  wire                pes_1_3_io_out_r_stall;
  wire       [15:0]   pes_1_3_io_out_c_data;
  wire                pes_1_3_io_out_c_is_stationary;
  wire       [15:0]   pes_2_0_io_out_r_data;
  wire                pes_2_0_io_out_r_load_store;
  wire                pes_2_0_io_out_r_df_is_ws;
  wire                pes_2_0_io_out_r_stall;
  wire       [15:0]   pes_2_0_io_out_c_data;
  wire                pes_2_0_io_out_c_is_stationary;
  wire       [15:0]   pes_2_1_io_out_r_data;
  wire                pes_2_1_io_out_r_load_store;
  wire                pes_2_1_io_out_r_df_is_ws;
  wire                pes_2_1_io_out_r_stall;
  wire       [15:0]   pes_2_1_io_out_c_data;
  wire                pes_2_1_io_out_c_is_stationary;
  wire       [15:0]   pes_2_2_io_out_r_data;
  wire                pes_2_2_io_out_r_load_store;
  wire                pes_2_2_io_out_r_df_is_ws;
  wire                pes_2_2_io_out_r_stall;
  wire       [15:0]   pes_2_2_io_out_c_data;
  wire                pes_2_2_io_out_c_is_stationary;
  wire       [15:0]   pes_2_3_io_out_r_data;
  wire                pes_2_3_io_out_r_load_store;
  wire                pes_2_3_io_out_r_df_is_ws;
  wire                pes_2_3_io_out_r_stall;
  wire       [15:0]   pes_2_3_io_out_c_data;
  wire                pes_2_3_io_out_c_is_stationary;
  wire       [15:0]   pes_3_0_io_out_r_data;
  wire                pes_3_0_io_out_r_load_store;
  wire                pes_3_0_io_out_r_df_is_ws;
  wire                pes_3_0_io_out_r_stall;
  wire       [15:0]   pes_3_0_io_out_c_data;
  wire                pes_3_0_io_out_c_is_stationary;
  wire       [15:0]   pes_3_1_io_out_r_data;
  wire                pes_3_1_io_out_r_load_store;
  wire                pes_3_1_io_out_r_df_is_ws;
  wire                pes_3_1_io_out_r_stall;
  wire       [15:0]   pes_3_1_io_out_c_data;
  wire                pes_3_1_io_out_c_is_stationary;
  wire       [15:0]   pes_3_2_io_out_r_data;
  wire                pes_3_2_io_out_r_load_store;
  wire                pes_3_2_io_out_r_df_is_ws;
  wire                pes_3_2_io_out_r_stall;
  wire       [15:0]   pes_3_2_io_out_c_data;
  wire                pes_3_2_io_out_c_is_stationary;
  wire       [15:0]   pes_3_3_io_out_r_data;
  wire                pes_3_3_io_out_r_load_store;
  wire                pes_3_3_io_out_r_df_is_ws;
  wire                pes_3_3_io_out_r_stall;
  wire       [15:0]   pes_3_3_io_out_c_data;
  wire                pes_3_3_io_out_c_is_stationary;
  wire       [15:0]   in_r_0_data;
  wire                in_r_0_load_store;
  wire                in_r_0_df_is_ws;
  wire                in_r_0_stall;
  wire       [15:0]   in_r_1_data;
  wire                in_r_1_load_store;
  wire                in_r_1_df_is_ws;
  wire                in_r_1_stall;
  wire       [15:0]   in_r_2_data;
  wire                in_r_2_load_store;
  wire                in_r_2_df_is_ws;
  wire                in_r_2_stall;
  wire       [15:0]   in_r_3_data;
  wire                in_r_3_load_store;
  wire                in_r_3_df_is_ws;
  wire                in_r_3_stall;
  wire       [15:0]   in_c_0_data;
  wire                in_c_0_is_stationary;
  wire       [15:0]   in_c_1_data;
  wire                in_c_1_is_stationary;
  wire       [15:0]   in_c_2_data;
  wire                in_c_2_is_stationary;
  wire       [15:0]   in_c_3_data;
  wire                in_c_3_is_stationary;
  wire       [15:0]   out_r_0_data;
  wire                out_r_0_load_store;
  wire                out_r_0_df_is_ws;
  wire                out_r_0_stall;
  wire       [15:0]   out_r_1_data;
  wire                out_r_1_load_store;
  wire                out_r_1_df_is_ws;
  wire                out_r_1_stall;
  wire       [15:0]   out_r_2_data;
  wire                out_r_2_load_store;
  wire                out_r_2_df_is_ws;
  wire                out_r_2_stall;
  wire       [15:0]   out_r_3_data;
  wire                out_r_3_load_store;
  wire                out_r_3_df_is_ws;
  wire                out_r_3_stall;
  wire       [15:0]   out_c_0_data;
  wire                out_c_0_is_stationary;
  wire       [15:0]   out_c_1_data;
  wire                out_c_1_is_stationary;
  wire       [15:0]   out_c_2_data;
  wire                out_c_2_is_stationary;
  wire       [15:0]   out_c_3_data;
  wire                out_c_3_is_stationary;
  reg        [15:0]   out_r_regNext_0_data;
  reg                 out_r_regNext_0_load_store;
  reg                 out_r_regNext_0_df_is_ws;
  reg                 out_r_regNext_0_stall;
  reg        [15:0]   out_r_regNext_1_data;
  reg                 out_r_regNext_1_load_store;
  reg                 out_r_regNext_1_df_is_ws;
  reg                 out_r_regNext_1_stall;
  reg        [15:0]   out_r_regNext_2_data;
  reg                 out_r_regNext_2_load_store;
  reg                 out_r_regNext_2_df_is_ws;
  reg                 out_r_regNext_2_stall;
  reg        [15:0]   out_r_regNext_3_data;
  reg                 out_r_regNext_3_load_store;
  reg                 out_r_regNext_3_df_is_ws;
  reg                 out_r_regNext_3_stall;
  reg        [15:0]   out_c_regNext_0_data;
  reg                 out_c_regNext_0_is_stationary;
  reg        [15:0]   out_c_regNext_1_data;
  reg                 out_c_regNext_1_is_stationary;
  reg        [15:0]   out_c_regNext_2_data;
  reg                 out_c_regNext_2_is_stationary;
  reg        [15:0]   out_c_regNext_3_data;
  reg                 out_c_regNext_3_is_stationary;
  reg        [15:0]   io_in_r_bypass_regNext_0_0_data;
  reg                 io_in_r_bypass_regNext_0_0_load_store;
  reg                 io_in_r_bypass_regNext_0_0_df_is_ws;
  reg                 io_in_r_bypass_regNext_0_0_stall;
  reg        [15:0]   io_in_r_bypass_regNext_0_1_data;
  reg                 io_in_r_bypass_regNext_0_1_load_store;
  reg                 io_in_r_bypass_regNext_0_1_df_is_ws;
  reg                 io_in_r_bypass_regNext_0_1_stall;
  reg        [15:0]   io_in_r_bypass_regNext_0_2_data;
  reg                 io_in_r_bypass_regNext_0_2_load_store;
  reg                 io_in_r_bypass_regNext_0_2_df_is_ws;
  reg                 io_in_r_bypass_regNext_0_2_stall;
  reg        [15:0]   io_in_r_bypass_regNext_0_3_data;
  reg                 io_in_r_bypass_regNext_0_3_load_store;
  reg                 io_in_r_bypass_regNext_0_3_df_is_ws;
  reg                 io_in_r_bypass_regNext_0_3_stall;
  reg        [15:0]   io_in_r_bypass_regNext_1_0_data;
  reg                 io_in_r_bypass_regNext_1_0_load_store;
  reg                 io_in_r_bypass_regNext_1_0_df_is_ws;
  reg                 io_in_r_bypass_regNext_1_0_stall;
  reg        [15:0]   io_in_r_bypass_regNext_1_1_data;
  reg                 io_in_r_bypass_regNext_1_1_load_store;
  reg                 io_in_r_bypass_regNext_1_1_df_is_ws;
  reg                 io_in_r_bypass_regNext_1_1_stall;
  reg        [15:0]   io_in_r_bypass_regNext_1_2_data;
  reg                 io_in_r_bypass_regNext_1_2_load_store;
  reg                 io_in_r_bypass_regNext_1_2_df_is_ws;
  reg                 io_in_r_bypass_regNext_1_2_stall;
  reg        [15:0]   io_in_r_bypass_regNext_1_3_data;
  reg                 io_in_r_bypass_regNext_1_3_load_store;
  reg                 io_in_r_bypass_regNext_1_3_df_is_ws;
  reg                 io_in_r_bypass_regNext_1_3_stall;
  reg        [15:0]   io_in_r_bypass_regNext_2_0_data;
  reg                 io_in_r_bypass_regNext_2_0_load_store;
  reg                 io_in_r_bypass_regNext_2_0_df_is_ws;
  reg                 io_in_r_bypass_regNext_2_0_stall;
  reg        [15:0]   io_in_r_bypass_regNext_2_1_data;
  reg                 io_in_r_bypass_regNext_2_1_load_store;
  reg                 io_in_r_bypass_regNext_2_1_df_is_ws;
  reg                 io_in_r_bypass_regNext_2_1_stall;
  reg        [15:0]   io_in_r_bypass_regNext_2_2_data;
  reg                 io_in_r_bypass_regNext_2_2_load_store;
  reg                 io_in_r_bypass_regNext_2_2_df_is_ws;
  reg                 io_in_r_bypass_regNext_2_2_stall;
  reg        [15:0]   io_in_r_bypass_regNext_2_3_data;
  reg                 io_in_r_bypass_regNext_2_3_load_store;
  reg                 io_in_r_bypass_regNext_2_3_df_is_ws;
  reg                 io_in_r_bypass_regNext_2_3_stall;
  reg        [15:0]   io_in_r_bypass_regNext_3_0_data;
  reg                 io_in_r_bypass_regNext_3_0_load_store;
  reg                 io_in_r_bypass_regNext_3_0_df_is_ws;
  reg                 io_in_r_bypass_regNext_3_0_stall;
  reg        [15:0]   io_in_r_bypass_regNext_3_1_data;
  reg                 io_in_r_bypass_regNext_3_1_load_store;
  reg                 io_in_r_bypass_regNext_3_1_df_is_ws;
  reg                 io_in_r_bypass_regNext_3_1_stall;
  reg        [15:0]   io_in_r_bypass_regNext_3_2_data;
  reg                 io_in_r_bypass_regNext_3_2_load_store;
  reg                 io_in_r_bypass_regNext_3_2_df_is_ws;
  reg                 io_in_r_bypass_regNext_3_2_stall;
  reg        [15:0]   io_in_r_bypass_regNext_3_3_data;
  reg                 io_in_r_bypass_regNext_3_3_load_store;
  reg                 io_in_r_bypass_regNext_3_3_df_is_ws;
  reg                 io_in_r_bypass_regNext_3_3_stall;
  reg        [15:0]   io_in_r_bypass_regNext_4_0_data;
  reg                 io_in_r_bypass_regNext_4_0_load_store;
  reg                 io_in_r_bypass_regNext_4_0_df_is_ws;
  reg                 io_in_r_bypass_regNext_4_0_stall;
  reg        [15:0]   io_in_r_bypass_regNext_4_1_data;
  reg                 io_in_r_bypass_regNext_4_1_load_store;
  reg                 io_in_r_bypass_regNext_4_1_df_is_ws;
  reg                 io_in_r_bypass_regNext_4_1_stall;
  reg        [15:0]   io_in_r_bypass_regNext_4_2_data;
  reg                 io_in_r_bypass_regNext_4_2_load_store;
  reg                 io_in_r_bypass_regNext_4_2_df_is_ws;
  reg                 io_in_r_bypass_regNext_4_2_stall;
  reg        [15:0]   io_in_r_bypass_regNext_4_3_data;
  reg                 io_in_r_bypass_regNext_4_3_load_store;
  reg                 io_in_r_bypass_regNext_4_3_df_is_ws;
  reg                 io_in_r_bypass_regNext_4_3_stall;
  reg        [15:0]   io_in_r_bypass_regNext_5_0_data;
  reg                 io_in_r_bypass_regNext_5_0_load_store;
  reg                 io_in_r_bypass_regNext_5_0_df_is_ws;
  reg                 io_in_r_bypass_regNext_5_0_stall;
  reg        [15:0]   io_in_r_bypass_regNext_5_1_data;
  reg                 io_in_r_bypass_regNext_5_1_load_store;
  reg                 io_in_r_bypass_regNext_5_1_df_is_ws;
  reg                 io_in_r_bypass_regNext_5_1_stall;
  reg        [15:0]   io_in_r_bypass_regNext_5_2_data;
  reg                 io_in_r_bypass_regNext_5_2_load_store;
  reg                 io_in_r_bypass_regNext_5_2_df_is_ws;
  reg                 io_in_r_bypass_regNext_5_2_stall;
  reg        [15:0]   io_in_r_bypass_regNext_5_3_data;
  reg                 io_in_r_bypass_regNext_5_3_load_store;
  reg                 io_in_r_bypass_regNext_5_3_df_is_ws;
  reg                 io_in_r_bypass_regNext_5_3_stall;
  reg        [15:0]   io_in_r_bypass_regNext_6_0_data;
  reg                 io_in_r_bypass_regNext_6_0_load_store;
  reg                 io_in_r_bypass_regNext_6_0_df_is_ws;
  reg                 io_in_r_bypass_regNext_6_0_stall;
  reg        [15:0]   io_in_r_bypass_regNext_6_1_data;
  reg                 io_in_r_bypass_regNext_6_1_load_store;
  reg                 io_in_r_bypass_regNext_6_1_df_is_ws;
  reg                 io_in_r_bypass_regNext_6_1_stall;
  reg        [15:0]   io_in_r_bypass_regNext_6_2_data;
  reg                 io_in_r_bypass_regNext_6_2_load_store;
  reg                 io_in_r_bypass_regNext_6_2_df_is_ws;
  reg                 io_in_r_bypass_regNext_6_2_stall;
  reg        [15:0]   io_in_r_bypass_regNext_6_3_data;
  reg                 io_in_r_bypass_regNext_6_3_load_store;
  reg                 io_in_r_bypass_regNext_6_3_df_is_ws;
  reg                 io_in_r_bypass_regNext_6_3_stall;
  reg        [15:0]   io_in_r_bypass_regNext_7_0_data;
  reg                 io_in_r_bypass_regNext_7_0_load_store;
  reg                 io_in_r_bypass_regNext_7_0_df_is_ws;
  reg                 io_in_r_bypass_regNext_7_0_stall;
  reg        [15:0]   io_in_r_bypass_regNext_7_1_data;
  reg                 io_in_r_bypass_regNext_7_1_load_store;
  reg                 io_in_r_bypass_regNext_7_1_df_is_ws;
  reg                 io_in_r_bypass_regNext_7_1_stall;
  reg        [15:0]   io_in_r_bypass_regNext_7_2_data;
  reg                 io_in_r_bypass_regNext_7_2_load_store;
  reg                 io_in_r_bypass_regNext_7_2_df_is_ws;
  reg                 io_in_r_bypass_regNext_7_2_stall;
  reg        [15:0]   io_in_r_bypass_regNext_7_3_data;
  reg                 io_in_r_bypass_regNext_7_3_load_store;
  reg                 io_in_r_bypass_regNext_7_3_df_is_ws;
  reg                 io_in_r_bypass_regNext_7_3_stall;
  reg        [15:0]   io_in_r_bypass_regNext_8_0_data;
  reg                 io_in_r_bypass_regNext_8_0_load_store;
  reg                 io_in_r_bypass_regNext_8_0_df_is_ws;
  reg                 io_in_r_bypass_regNext_8_0_stall;
  reg        [15:0]   io_in_r_bypass_regNext_8_1_data;
  reg                 io_in_r_bypass_regNext_8_1_load_store;
  reg                 io_in_r_bypass_regNext_8_1_df_is_ws;
  reg                 io_in_r_bypass_regNext_8_1_stall;
  reg        [15:0]   io_in_r_bypass_regNext_8_2_data;
  reg                 io_in_r_bypass_regNext_8_2_load_store;
  reg                 io_in_r_bypass_regNext_8_2_df_is_ws;
  reg                 io_in_r_bypass_regNext_8_2_stall;
  reg        [15:0]   io_in_r_bypass_regNext_8_3_data;
  reg                 io_in_r_bypass_regNext_8_3_load_store;
  reg                 io_in_r_bypass_regNext_8_3_df_is_ws;
  reg                 io_in_r_bypass_regNext_8_3_stall;
  reg        [15:0]   io_in_r_bypass_regNext_9_0_data;
  reg                 io_in_r_bypass_regNext_9_0_load_store;
  reg                 io_in_r_bypass_regNext_9_0_df_is_ws;
  reg                 io_in_r_bypass_regNext_9_0_stall;
  reg        [15:0]   io_in_r_bypass_regNext_9_1_data;
  reg                 io_in_r_bypass_regNext_9_1_load_store;
  reg                 io_in_r_bypass_regNext_9_1_df_is_ws;
  reg                 io_in_r_bypass_regNext_9_1_stall;
  reg        [15:0]   io_in_r_bypass_regNext_9_2_data;
  reg                 io_in_r_bypass_regNext_9_2_load_store;
  reg                 io_in_r_bypass_regNext_9_2_df_is_ws;
  reg                 io_in_r_bypass_regNext_9_2_stall;
  reg        [15:0]   io_in_r_bypass_regNext_9_3_data;
  reg                 io_in_r_bypass_regNext_9_3_load_store;
  reg                 io_in_r_bypass_regNext_9_3_df_is_ws;
  reg                 io_in_r_bypass_regNext_9_3_stall;
  reg        [15:0]   io_in_r_bypass_regNext_10_0_data;
  reg                 io_in_r_bypass_regNext_10_0_load_store;
  reg                 io_in_r_bypass_regNext_10_0_df_is_ws;
  reg                 io_in_r_bypass_regNext_10_0_stall;
  reg        [15:0]   io_in_r_bypass_regNext_10_1_data;
  reg                 io_in_r_bypass_regNext_10_1_load_store;
  reg                 io_in_r_bypass_regNext_10_1_df_is_ws;
  reg                 io_in_r_bypass_regNext_10_1_stall;
  reg        [15:0]   io_in_r_bypass_regNext_10_2_data;
  reg                 io_in_r_bypass_regNext_10_2_load_store;
  reg                 io_in_r_bypass_regNext_10_2_df_is_ws;
  reg                 io_in_r_bypass_regNext_10_2_stall;
  reg        [15:0]   io_in_r_bypass_regNext_10_3_data;
  reg                 io_in_r_bypass_regNext_10_3_load_store;
  reg                 io_in_r_bypass_regNext_10_3_df_is_ws;
  reg                 io_in_r_bypass_regNext_10_3_stall;
  reg        [15:0]   io_in_r_bypass_regNext_11_0_data;
  reg                 io_in_r_bypass_regNext_11_0_load_store;
  reg                 io_in_r_bypass_regNext_11_0_df_is_ws;
  reg                 io_in_r_bypass_regNext_11_0_stall;
  reg        [15:0]   io_in_r_bypass_regNext_11_1_data;
  reg                 io_in_r_bypass_regNext_11_1_load_store;
  reg                 io_in_r_bypass_regNext_11_1_df_is_ws;
  reg                 io_in_r_bypass_regNext_11_1_stall;
  reg        [15:0]   io_in_r_bypass_regNext_11_2_data;
  reg                 io_in_r_bypass_regNext_11_2_load_store;
  reg                 io_in_r_bypass_regNext_11_2_df_is_ws;
  reg                 io_in_r_bypass_regNext_11_2_stall;
  reg        [15:0]   io_in_r_bypass_regNext_11_3_data;
  reg                 io_in_r_bypass_regNext_11_3_load_store;
  reg                 io_in_r_bypass_regNext_11_3_df_is_ws;
  reg                 io_in_r_bypass_regNext_11_3_stall;
  reg        [15:0]   io_in_r_bypass_regNext_12_0_data;
  reg                 io_in_r_bypass_regNext_12_0_load_store;
  reg                 io_in_r_bypass_regNext_12_0_df_is_ws;
  reg                 io_in_r_bypass_regNext_12_0_stall;
  reg        [15:0]   io_in_r_bypass_regNext_12_1_data;
  reg                 io_in_r_bypass_regNext_12_1_load_store;
  reg                 io_in_r_bypass_regNext_12_1_df_is_ws;
  reg                 io_in_r_bypass_regNext_12_1_stall;
  reg        [15:0]   io_in_r_bypass_regNext_12_2_data;
  reg                 io_in_r_bypass_regNext_12_2_load_store;
  reg                 io_in_r_bypass_regNext_12_2_df_is_ws;
  reg                 io_in_r_bypass_regNext_12_2_stall;
  reg        [15:0]   io_in_r_bypass_regNext_12_3_data;
  reg                 io_in_r_bypass_regNext_12_3_load_store;
  reg                 io_in_r_bypass_regNext_12_3_df_is_ws;
  reg                 io_in_r_bypass_regNext_12_3_stall;
  reg        [15:0]   io_in_r_bypass_regNext_13_0_data;
  reg                 io_in_r_bypass_regNext_13_0_load_store;
  reg                 io_in_r_bypass_regNext_13_0_df_is_ws;
  reg                 io_in_r_bypass_regNext_13_0_stall;
  reg        [15:0]   io_in_r_bypass_regNext_13_1_data;
  reg                 io_in_r_bypass_regNext_13_1_load_store;
  reg                 io_in_r_bypass_regNext_13_1_df_is_ws;
  reg                 io_in_r_bypass_regNext_13_1_stall;
  reg        [15:0]   io_in_r_bypass_regNext_13_2_data;
  reg                 io_in_r_bypass_regNext_13_2_load_store;
  reg                 io_in_r_bypass_regNext_13_2_df_is_ws;
  reg                 io_in_r_bypass_regNext_13_2_stall;
  reg        [15:0]   io_in_r_bypass_regNext_13_3_data;
  reg                 io_in_r_bypass_regNext_13_3_load_store;
  reg                 io_in_r_bypass_regNext_13_3_df_is_ws;
  reg                 io_in_r_bypass_regNext_13_3_stall;
  reg        [15:0]   io_in_r_bypass_regNext_14_0_data;
  reg                 io_in_r_bypass_regNext_14_0_load_store;
  reg                 io_in_r_bypass_regNext_14_0_df_is_ws;
  reg                 io_in_r_bypass_regNext_14_0_stall;
  reg        [15:0]   io_in_r_bypass_regNext_14_1_data;
  reg                 io_in_r_bypass_regNext_14_1_load_store;
  reg                 io_in_r_bypass_regNext_14_1_df_is_ws;
  reg                 io_in_r_bypass_regNext_14_1_stall;
  reg        [15:0]   io_in_r_bypass_regNext_14_2_data;
  reg                 io_in_r_bypass_regNext_14_2_load_store;
  reg                 io_in_r_bypass_regNext_14_2_df_is_ws;
  reg                 io_in_r_bypass_regNext_14_2_stall;
  reg        [15:0]   io_in_r_bypass_regNext_14_3_data;
  reg                 io_in_r_bypass_regNext_14_3_load_store;
  reg                 io_in_r_bypass_regNext_14_3_df_is_ws;
  reg                 io_in_r_bypass_regNext_14_3_stall;
  reg        [15:0]   io_in_r_bypass_regNext_15_0_data;
  reg                 io_in_r_bypass_regNext_15_0_load_store;
  reg                 io_in_r_bypass_regNext_15_0_df_is_ws;
  reg                 io_in_r_bypass_regNext_15_0_stall;
  reg        [15:0]   io_in_r_bypass_regNext_15_1_data;
  reg                 io_in_r_bypass_regNext_15_1_load_store;
  reg                 io_in_r_bypass_regNext_15_1_df_is_ws;
  reg                 io_in_r_bypass_regNext_15_1_stall;
  reg        [15:0]   io_in_r_bypass_regNext_15_2_data;
  reg                 io_in_r_bypass_regNext_15_2_load_store;
  reg                 io_in_r_bypass_regNext_15_2_df_is_ws;
  reg                 io_in_r_bypass_regNext_15_2_stall;
  reg        [15:0]   io_in_r_bypass_regNext_15_3_data;
  reg                 io_in_r_bypass_regNext_15_3_load_store;
  reg                 io_in_r_bypass_regNext_15_3_df_is_ws;
  reg                 io_in_r_bypass_regNext_15_3_stall;
  reg        [15:0]   io_in_r_bypass_regNext_16_0_data;
  reg                 io_in_r_bypass_regNext_16_0_load_store;
  reg                 io_in_r_bypass_regNext_16_0_df_is_ws;
  reg                 io_in_r_bypass_regNext_16_0_stall;
  reg        [15:0]   io_in_r_bypass_regNext_16_1_data;
  reg                 io_in_r_bypass_regNext_16_1_load_store;
  reg                 io_in_r_bypass_regNext_16_1_df_is_ws;
  reg                 io_in_r_bypass_regNext_16_1_stall;
  reg        [15:0]   io_in_r_bypass_regNext_16_2_data;
  reg                 io_in_r_bypass_regNext_16_2_load_store;
  reg                 io_in_r_bypass_regNext_16_2_df_is_ws;
  reg                 io_in_r_bypass_regNext_16_2_stall;
  reg        [15:0]   io_in_r_bypass_regNext_16_3_data;
  reg                 io_in_r_bypass_regNext_16_3_load_store;
  reg                 io_in_r_bypass_regNext_16_3_df_is_ws;
  reg                 io_in_r_bypass_regNext_16_3_stall;
  reg        [15:0]   io_in_r_bypass_regNext_17_0_data;
  reg                 io_in_r_bypass_regNext_17_0_load_store;
  reg                 io_in_r_bypass_regNext_17_0_df_is_ws;
  reg                 io_in_r_bypass_regNext_17_0_stall;
  reg        [15:0]   io_in_r_bypass_regNext_17_1_data;
  reg                 io_in_r_bypass_regNext_17_1_load_store;
  reg                 io_in_r_bypass_regNext_17_1_df_is_ws;
  reg                 io_in_r_bypass_regNext_17_1_stall;
  reg        [15:0]   io_in_r_bypass_regNext_17_2_data;
  reg                 io_in_r_bypass_regNext_17_2_load_store;
  reg                 io_in_r_bypass_regNext_17_2_df_is_ws;
  reg                 io_in_r_bypass_regNext_17_2_stall;
  reg        [15:0]   io_in_r_bypass_regNext_17_3_data;
  reg                 io_in_r_bypass_regNext_17_3_load_store;
  reg                 io_in_r_bypass_regNext_17_3_df_is_ws;
  reg                 io_in_r_bypass_regNext_17_3_stall;
  reg        [15:0]   io_in_r_bypass_regNext_18_0_data;
  reg                 io_in_r_bypass_regNext_18_0_load_store;
  reg                 io_in_r_bypass_regNext_18_0_df_is_ws;
  reg                 io_in_r_bypass_regNext_18_0_stall;
  reg        [15:0]   io_in_r_bypass_regNext_18_1_data;
  reg                 io_in_r_bypass_regNext_18_1_load_store;
  reg                 io_in_r_bypass_regNext_18_1_df_is_ws;
  reg                 io_in_r_bypass_regNext_18_1_stall;
  reg        [15:0]   io_in_r_bypass_regNext_18_2_data;
  reg                 io_in_r_bypass_regNext_18_2_load_store;
  reg                 io_in_r_bypass_regNext_18_2_df_is_ws;
  reg                 io_in_r_bypass_regNext_18_2_stall;
  reg        [15:0]   io_in_r_bypass_regNext_18_3_data;
  reg                 io_in_r_bypass_regNext_18_3_load_store;
  reg                 io_in_r_bypass_regNext_18_3_df_is_ws;
  reg                 io_in_r_bypass_regNext_18_3_stall;
  reg        [15:0]   io_in_r_bypass_regNext_19_0_data;
  reg                 io_in_r_bypass_regNext_19_0_load_store;
  reg                 io_in_r_bypass_regNext_19_0_df_is_ws;
  reg                 io_in_r_bypass_regNext_19_0_stall;
  reg        [15:0]   io_in_r_bypass_regNext_19_1_data;
  reg                 io_in_r_bypass_regNext_19_1_load_store;
  reg                 io_in_r_bypass_regNext_19_1_df_is_ws;
  reg                 io_in_r_bypass_regNext_19_1_stall;
  reg        [15:0]   io_in_r_bypass_regNext_19_2_data;
  reg                 io_in_r_bypass_regNext_19_2_load_store;
  reg                 io_in_r_bypass_regNext_19_2_df_is_ws;
  reg                 io_in_r_bypass_regNext_19_2_stall;
  reg        [15:0]   io_in_r_bypass_regNext_19_3_data;
  reg                 io_in_r_bypass_regNext_19_3_load_store;
  reg                 io_in_r_bypass_regNext_19_3_df_is_ws;
  reg                 io_in_r_bypass_regNext_19_3_stall;
  reg        [15:0]   io_in_r_bypass_regNext_20_0_data;
  reg                 io_in_r_bypass_regNext_20_0_load_store;
  reg                 io_in_r_bypass_regNext_20_0_df_is_ws;
  reg                 io_in_r_bypass_regNext_20_0_stall;
  reg        [15:0]   io_in_r_bypass_regNext_20_1_data;
  reg                 io_in_r_bypass_regNext_20_1_load_store;
  reg                 io_in_r_bypass_regNext_20_1_df_is_ws;
  reg                 io_in_r_bypass_regNext_20_1_stall;
  reg        [15:0]   io_in_r_bypass_regNext_20_2_data;
  reg                 io_in_r_bypass_regNext_20_2_load_store;
  reg                 io_in_r_bypass_regNext_20_2_df_is_ws;
  reg                 io_in_r_bypass_regNext_20_2_stall;
  reg        [15:0]   io_in_r_bypass_regNext_20_3_data;
  reg                 io_in_r_bypass_regNext_20_3_load_store;
  reg                 io_in_r_bypass_regNext_20_3_df_is_ws;
  reg                 io_in_r_bypass_regNext_20_3_stall;
  reg        [15:0]   io_in_r_bypass_regNext_21_0_data;
  reg                 io_in_r_bypass_regNext_21_0_load_store;
  reg                 io_in_r_bypass_regNext_21_0_df_is_ws;
  reg                 io_in_r_bypass_regNext_21_0_stall;
  reg        [15:0]   io_in_r_bypass_regNext_21_1_data;
  reg                 io_in_r_bypass_regNext_21_1_load_store;
  reg                 io_in_r_bypass_regNext_21_1_df_is_ws;
  reg                 io_in_r_bypass_regNext_21_1_stall;
  reg        [15:0]   io_in_r_bypass_regNext_21_2_data;
  reg                 io_in_r_bypass_regNext_21_2_load_store;
  reg                 io_in_r_bypass_regNext_21_2_df_is_ws;
  reg                 io_in_r_bypass_regNext_21_2_stall;
  reg        [15:0]   io_in_r_bypass_regNext_21_3_data;
  reg                 io_in_r_bypass_regNext_21_3_load_store;
  reg                 io_in_r_bypass_regNext_21_3_df_is_ws;
  reg                 io_in_r_bypass_regNext_21_3_stall;
  reg        [15:0]   io_in_r_bypass_regNext_22_0_data;
  reg                 io_in_r_bypass_regNext_22_0_load_store;
  reg                 io_in_r_bypass_regNext_22_0_df_is_ws;
  reg                 io_in_r_bypass_regNext_22_0_stall;
  reg        [15:0]   io_in_r_bypass_regNext_22_1_data;
  reg                 io_in_r_bypass_regNext_22_1_load_store;
  reg                 io_in_r_bypass_regNext_22_1_df_is_ws;
  reg                 io_in_r_bypass_regNext_22_1_stall;
  reg        [15:0]   io_in_r_bypass_regNext_22_2_data;
  reg                 io_in_r_bypass_regNext_22_2_load_store;
  reg                 io_in_r_bypass_regNext_22_2_df_is_ws;
  reg                 io_in_r_bypass_regNext_22_2_stall;
  reg        [15:0]   io_in_r_bypass_regNext_22_3_data;
  reg                 io_in_r_bypass_regNext_22_3_load_store;
  reg                 io_in_r_bypass_regNext_22_3_df_is_ws;
  reg                 io_in_r_bypass_regNext_22_3_stall;
  reg        [15:0]   io_in_r_bypass_regNext_23_0_data;
  reg                 io_in_r_bypass_regNext_23_0_load_store;
  reg                 io_in_r_bypass_regNext_23_0_df_is_ws;
  reg                 io_in_r_bypass_regNext_23_0_stall;
  reg        [15:0]   io_in_r_bypass_regNext_23_1_data;
  reg                 io_in_r_bypass_regNext_23_1_load_store;
  reg                 io_in_r_bypass_regNext_23_1_df_is_ws;
  reg                 io_in_r_bypass_regNext_23_1_stall;
  reg        [15:0]   io_in_r_bypass_regNext_23_2_data;
  reg                 io_in_r_bypass_regNext_23_2_load_store;
  reg                 io_in_r_bypass_regNext_23_2_df_is_ws;
  reg                 io_in_r_bypass_regNext_23_2_stall;
  reg        [15:0]   io_in_r_bypass_regNext_23_3_data;
  reg                 io_in_r_bypass_regNext_23_3_load_store;
  reg                 io_in_r_bypass_regNext_23_3_df_is_ws;
  reg                 io_in_r_bypass_regNext_23_3_stall;
  reg        [15:0]   io_in_r_bypass_regNext_24_0_data;
  reg                 io_in_r_bypass_regNext_24_0_load_store;
  reg                 io_in_r_bypass_regNext_24_0_df_is_ws;
  reg                 io_in_r_bypass_regNext_24_0_stall;
  reg        [15:0]   io_in_r_bypass_regNext_24_1_data;
  reg                 io_in_r_bypass_regNext_24_1_load_store;
  reg                 io_in_r_bypass_regNext_24_1_df_is_ws;
  reg                 io_in_r_bypass_regNext_24_1_stall;
  reg        [15:0]   io_in_r_bypass_regNext_24_2_data;
  reg                 io_in_r_bypass_regNext_24_2_load_store;
  reg                 io_in_r_bypass_regNext_24_2_df_is_ws;
  reg                 io_in_r_bypass_regNext_24_2_stall;
  reg        [15:0]   io_in_r_bypass_regNext_24_3_data;
  reg                 io_in_r_bypass_regNext_24_3_load_store;
  reg                 io_in_r_bypass_regNext_24_3_df_is_ws;
  reg                 io_in_r_bypass_regNext_24_3_stall;
  reg        [15:0]   io_in_r_bypass_regNext_25_0_data;
  reg                 io_in_r_bypass_regNext_25_0_load_store;
  reg                 io_in_r_bypass_regNext_25_0_df_is_ws;
  reg                 io_in_r_bypass_regNext_25_0_stall;
  reg        [15:0]   io_in_r_bypass_regNext_25_1_data;
  reg                 io_in_r_bypass_regNext_25_1_load_store;
  reg                 io_in_r_bypass_regNext_25_1_df_is_ws;
  reg                 io_in_r_bypass_regNext_25_1_stall;
  reg        [15:0]   io_in_r_bypass_regNext_25_2_data;
  reg                 io_in_r_bypass_regNext_25_2_load_store;
  reg                 io_in_r_bypass_regNext_25_2_df_is_ws;
  reg                 io_in_r_bypass_regNext_25_2_stall;
  reg        [15:0]   io_in_r_bypass_regNext_25_3_data;
  reg                 io_in_r_bypass_regNext_25_3_load_store;
  reg                 io_in_r_bypass_regNext_25_3_df_is_ws;
  reg                 io_in_r_bypass_regNext_25_3_stall;
  reg        [15:0]   io_in_r_bypass_regNext_26_0_data;
  reg                 io_in_r_bypass_regNext_26_0_load_store;
  reg                 io_in_r_bypass_regNext_26_0_df_is_ws;
  reg                 io_in_r_bypass_regNext_26_0_stall;
  reg        [15:0]   io_in_r_bypass_regNext_26_1_data;
  reg                 io_in_r_bypass_regNext_26_1_load_store;
  reg                 io_in_r_bypass_regNext_26_1_df_is_ws;
  reg                 io_in_r_bypass_regNext_26_1_stall;
  reg        [15:0]   io_in_r_bypass_regNext_26_2_data;
  reg                 io_in_r_bypass_regNext_26_2_load_store;
  reg                 io_in_r_bypass_regNext_26_2_df_is_ws;
  reg                 io_in_r_bypass_regNext_26_2_stall;
  reg        [15:0]   io_in_r_bypass_regNext_26_3_data;
  reg                 io_in_r_bypass_regNext_26_3_load_store;
  reg                 io_in_r_bypass_regNext_26_3_df_is_ws;
  reg                 io_in_r_bypass_regNext_26_3_stall;
  reg        [15:0]   io_in_r_bypass_regNext_27_0_data;
  reg                 io_in_r_bypass_regNext_27_0_load_store;
  reg                 io_in_r_bypass_regNext_27_0_df_is_ws;
  reg                 io_in_r_bypass_regNext_27_0_stall;
  reg        [15:0]   io_in_r_bypass_regNext_27_1_data;
  reg                 io_in_r_bypass_regNext_27_1_load_store;
  reg                 io_in_r_bypass_regNext_27_1_df_is_ws;
  reg                 io_in_r_bypass_regNext_27_1_stall;
  reg        [15:0]   io_in_r_bypass_regNext_27_2_data;
  reg                 io_in_r_bypass_regNext_27_2_load_store;
  reg                 io_in_r_bypass_regNext_27_2_df_is_ws;
  reg                 io_in_r_bypass_regNext_27_2_stall;
  reg        [15:0]   io_in_r_bypass_regNext_27_3_data;
  reg                 io_in_r_bypass_regNext_27_3_load_store;
  reg                 io_in_r_bypass_regNext_27_3_df_is_ws;
  reg                 io_in_r_bypass_regNext_27_3_stall;
  reg        [15:0]   io_in_r_bypass_regNext_28_0_data;
  reg                 io_in_r_bypass_regNext_28_0_load_store;
  reg                 io_in_r_bypass_regNext_28_0_df_is_ws;
  reg                 io_in_r_bypass_regNext_28_0_stall;
  reg        [15:0]   io_in_r_bypass_regNext_28_1_data;
  reg                 io_in_r_bypass_regNext_28_1_load_store;
  reg                 io_in_r_bypass_regNext_28_1_df_is_ws;
  reg                 io_in_r_bypass_regNext_28_1_stall;
  reg        [15:0]   io_in_r_bypass_regNext_28_2_data;
  reg                 io_in_r_bypass_regNext_28_2_load_store;
  reg                 io_in_r_bypass_regNext_28_2_df_is_ws;
  reg                 io_in_r_bypass_regNext_28_2_stall;
  reg        [15:0]   io_in_r_bypass_regNext_28_3_data;
  reg                 io_in_r_bypass_regNext_28_3_load_store;
  reg                 io_in_r_bypass_regNext_28_3_df_is_ws;
  reg                 io_in_r_bypass_regNext_28_3_stall;
  reg        [15:0]   io_in_r_bypass_regNext_29_0_data;
  reg                 io_in_r_bypass_regNext_29_0_load_store;
  reg                 io_in_r_bypass_regNext_29_0_df_is_ws;
  reg                 io_in_r_bypass_regNext_29_0_stall;
  reg        [15:0]   io_in_r_bypass_regNext_29_1_data;
  reg                 io_in_r_bypass_regNext_29_1_load_store;
  reg                 io_in_r_bypass_regNext_29_1_df_is_ws;
  reg                 io_in_r_bypass_regNext_29_1_stall;
  reg        [15:0]   io_in_r_bypass_regNext_29_2_data;
  reg                 io_in_r_bypass_regNext_29_2_load_store;
  reg                 io_in_r_bypass_regNext_29_2_df_is_ws;
  reg                 io_in_r_bypass_regNext_29_2_stall;
  reg        [15:0]   io_in_r_bypass_regNext_29_3_data;
  reg                 io_in_r_bypass_regNext_29_3_load_store;
  reg                 io_in_r_bypass_regNext_29_3_df_is_ws;
  reg                 io_in_r_bypass_regNext_29_3_stall;
  reg        [15:0]   io_in_r_bypass_regNext_30_0_data;
  reg                 io_in_r_bypass_regNext_30_0_load_store;
  reg                 io_in_r_bypass_regNext_30_0_df_is_ws;
  reg                 io_in_r_bypass_regNext_30_0_stall;
  reg        [15:0]   io_in_r_bypass_regNext_30_1_data;
  reg                 io_in_r_bypass_regNext_30_1_load_store;
  reg                 io_in_r_bypass_regNext_30_1_df_is_ws;
  reg                 io_in_r_bypass_regNext_30_1_stall;
  reg        [15:0]   io_in_r_bypass_regNext_30_2_data;
  reg                 io_in_r_bypass_regNext_30_2_load_store;
  reg                 io_in_r_bypass_regNext_30_2_df_is_ws;
  reg                 io_in_r_bypass_regNext_30_2_stall;
  reg        [15:0]   io_in_r_bypass_regNext_30_3_data;
  reg                 io_in_r_bypass_regNext_30_3_load_store;
  reg                 io_in_r_bypass_regNext_30_3_df_is_ws;
  reg                 io_in_r_bypass_regNext_30_3_stall;
  reg        [15:0]   io_in_r_bypass_regNext_31_0_data;
  reg                 io_in_r_bypass_regNext_31_0_load_store;
  reg                 io_in_r_bypass_regNext_31_0_df_is_ws;
  reg                 io_in_r_bypass_regNext_31_0_stall;
  reg        [15:0]   io_in_r_bypass_regNext_31_1_data;
  reg                 io_in_r_bypass_regNext_31_1_load_store;
  reg                 io_in_r_bypass_regNext_31_1_df_is_ws;
  reg                 io_in_r_bypass_regNext_31_1_stall;
  reg        [15:0]   io_in_r_bypass_regNext_31_2_data;
  reg                 io_in_r_bypass_regNext_31_2_load_store;
  reg                 io_in_r_bypass_regNext_31_2_df_is_ws;
  reg                 io_in_r_bypass_regNext_31_2_stall;
  reg        [15:0]   io_in_r_bypass_regNext_31_3_data;
  reg                 io_in_r_bypass_regNext_31_3_load_store;
  reg                 io_in_r_bypass_regNext_31_3_df_is_ws;
  reg                 io_in_r_bypass_regNext_31_3_stall;
  reg        [15:0]   io_in_r_bypass_regNext_0_0_data_1;
  reg                 io_in_r_bypass_regNext_0_0_load_store_1;
  reg                 io_in_r_bypass_regNext_0_0_df_is_ws_1;
  reg                 io_in_r_bypass_regNext_0_0_stall_1;
  reg        [15:0]   io_in_r_bypass_regNext_0_1_data_1;
  reg                 io_in_r_bypass_regNext_0_1_load_store_1;
  reg                 io_in_r_bypass_regNext_0_1_df_is_ws_1;
  reg                 io_in_r_bypass_regNext_0_1_stall_1;
  reg        [15:0]   io_in_r_bypass_regNext_0_2_data_1;
  reg                 io_in_r_bypass_regNext_0_2_load_store_1;
  reg                 io_in_r_bypass_regNext_0_2_df_is_ws_1;
  reg                 io_in_r_bypass_regNext_0_2_stall_1;
  reg        [15:0]   io_in_r_bypass_regNext_0_3_data_1;
  reg                 io_in_r_bypass_regNext_0_3_load_store_1;
  reg                 io_in_r_bypass_regNext_0_3_df_is_ws_1;
  reg                 io_in_r_bypass_regNext_0_3_stall_1;
  reg        [15:0]   io_in_r_bypass_regNext_1_0_data_1;
  reg                 io_in_r_bypass_regNext_1_0_load_store_1;
  reg                 io_in_r_bypass_regNext_1_0_df_is_ws_1;
  reg                 io_in_r_bypass_regNext_1_0_stall_1;
  reg        [15:0]   io_in_r_bypass_regNext_1_1_data_1;
  reg                 io_in_r_bypass_regNext_1_1_load_store_1;
  reg                 io_in_r_bypass_regNext_1_1_df_is_ws_1;
  reg                 io_in_r_bypass_regNext_1_1_stall_1;
  reg        [15:0]   io_in_r_bypass_regNext_1_2_data_1;
  reg                 io_in_r_bypass_regNext_1_2_load_store_1;
  reg                 io_in_r_bypass_regNext_1_2_df_is_ws_1;
  reg                 io_in_r_bypass_regNext_1_2_stall_1;
  reg        [15:0]   io_in_r_bypass_regNext_1_3_data_1;
  reg                 io_in_r_bypass_regNext_1_3_load_store_1;
  reg                 io_in_r_bypass_regNext_1_3_df_is_ws_1;
  reg                 io_in_r_bypass_regNext_1_3_stall_1;
  reg        [15:0]   io_in_r_bypass_regNext_2_0_data_1;
  reg                 io_in_r_bypass_regNext_2_0_load_store_1;
  reg                 io_in_r_bypass_regNext_2_0_df_is_ws_1;
  reg                 io_in_r_bypass_regNext_2_0_stall_1;
  reg        [15:0]   io_in_r_bypass_regNext_2_1_data_1;
  reg                 io_in_r_bypass_regNext_2_1_load_store_1;
  reg                 io_in_r_bypass_regNext_2_1_df_is_ws_1;
  reg                 io_in_r_bypass_regNext_2_1_stall_1;
  reg        [15:0]   io_in_r_bypass_regNext_2_2_data_1;
  reg                 io_in_r_bypass_regNext_2_2_load_store_1;
  reg                 io_in_r_bypass_regNext_2_2_df_is_ws_1;
  reg                 io_in_r_bypass_regNext_2_2_stall_1;
  reg        [15:0]   io_in_r_bypass_regNext_2_3_data_1;
  reg                 io_in_r_bypass_regNext_2_3_load_store_1;
  reg                 io_in_r_bypass_regNext_2_3_df_is_ws_1;
  reg                 io_in_r_bypass_regNext_2_3_stall_1;
  reg        [15:0]   io_in_r_bypass_regNext_3_0_data_1;
  reg                 io_in_r_bypass_regNext_3_0_load_store_1;
  reg                 io_in_r_bypass_regNext_3_0_df_is_ws_1;
  reg                 io_in_r_bypass_regNext_3_0_stall_1;
  reg        [15:0]   io_in_r_bypass_regNext_3_1_data_1;
  reg                 io_in_r_bypass_regNext_3_1_load_store_1;
  reg                 io_in_r_bypass_regNext_3_1_df_is_ws_1;
  reg                 io_in_r_bypass_regNext_3_1_stall_1;
  reg        [15:0]   io_in_r_bypass_regNext_3_2_data_1;
  reg                 io_in_r_bypass_regNext_3_2_load_store_1;
  reg                 io_in_r_bypass_regNext_3_2_df_is_ws_1;
  reg                 io_in_r_bypass_regNext_3_2_stall_1;
  reg        [15:0]   io_in_r_bypass_regNext_3_3_data_1;
  reg                 io_in_r_bypass_regNext_3_3_load_store_1;
  reg                 io_in_r_bypass_regNext_3_3_df_is_ws_1;
  reg                 io_in_r_bypass_regNext_3_3_stall_1;
  reg        [15:0]   io_in_r_bypass_regNext_4_0_data_1;
  reg                 io_in_r_bypass_regNext_4_0_load_store_1;
  reg                 io_in_r_bypass_regNext_4_0_df_is_ws_1;
  reg                 io_in_r_bypass_regNext_4_0_stall_1;
  reg        [15:0]   io_in_r_bypass_regNext_4_1_data_1;
  reg                 io_in_r_bypass_regNext_4_1_load_store_1;
  reg                 io_in_r_bypass_regNext_4_1_df_is_ws_1;
  reg                 io_in_r_bypass_regNext_4_1_stall_1;
  reg        [15:0]   io_in_r_bypass_regNext_4_2_data_1;
  reg                 io_in_r_bypass_regNext_4_2_load_store_1;
  reg                 io_in_r_bypass_regNext_4_2_df_is_ws_1;
  reg                 io_in_r_bypass_regNext_4_2_stall_1;
  reg        [15:0]   io_in_r_bypass_regNext_4_3_data_1;
  reg                 io_in_r_bypass_regNext_4_3_load_store_1;
  reg                 io_in_r_bypass_regNext_4_3_df_is_ws_1;
  reg                 io_in_r_bypass_regNext_4_3_stall_1;
  reg        [15:0]   io_in_r_bypass_regNext_5_0_data_1;
  reg                 io_in_r_bypass_regNext_5_0_load_store_1;
  reg                 io_in_r_bypass_regNext_5_0_df_is_ws_1;
  reg                 io_in_r_bypass_regNext_5_0_stall_1;
  reg        [15:0]   io_in_r_bypass_regNext_5_1_data_1;
  reg                 io_in_r_bypass_regNext_5_1_load_store_1;
  reg                 io_in_r_bypass_regNext_5_1_df_is_ws_1;
  reg                 io_in_r_bypass_regNext_5_1_stall_1;
  reg        [15:0]   io_in_r_bypass_regNext_5_2_data_1;
  reg                 io_in_r_bypass_regNext_5_2_load_store_1;
  reg                 io_in_r_bypass_regNext_5_2_df_is_ws_1;
  reg                 io_in_r_bypass_regNext_5_2_stall_1;
  reg        [15:0]   io_in_r_bypass_regNext_5_3_data_1;
  reg                 io_in_r_bypass_regNext_5_3_load_store_1;
  reg                 io_in_r_bypass_regNext_5_3_df_is_ws_1;
  reg                 io_in_r_bypass_regNext_5_3_stall_1;
  reg        [15:0]   io_in_r_bypass_regNext_6_0_data_1;
  reg                 io_in_r_bypass_regNext_6_0_load_store_1;
  reg                 io_in_r_bypass_regNext_6_0_df_is_ws_1;
  reg                 io_in_r_bypass_regNext_6_0_stall_1;
  reg        [15:0]   io_in_r_bypass_regNext_6_1_data_1;
  reg                 io_in_r_bypass_regNext_6_1_load_store_1;
  reg                 io_in_r_bypass_regNext_6_1_df_is_ws_1;
  reg                 io_in_r_bypass_regNext_6_1_stall_1;
  reg        [15:0]   io_in_r_bypass_regNext_6_2_data_1;
  reg                 io_in_r_bypass_regNext_6_2_load_store_1;
  reg                 io_in_r_bypass_regNext_6_2_df_is_ws_1;
  reg                 io_in_r_bypass_regNext_6_2_stall_1;
  reg        [15:0]   io_in_r_bypass_regNext_6_3_data_1;
  reg                 io_in_r_bypass_regNext_6_3_load_store_1;
  reg                 io_in_r_bypass_regNext_6_3_df_is_ws_1;
  reg                 io_in_r_bypass_regNext_6_3_stall_1;
  reg        [15:0]   io_in_r_bypass_regNext_7_0_data_1;
  reg                 io_in_r_bypass_regNext_7_0_load_store_1;
  reg                 io_in_r_bypass_regNext_7_0_df_is_ws_1;
  reg                 io_in_r_bypass_regNext_7_0_stall_1;
  reg        [15:0]   io_in_r_bypass_regNext_7_1_data_1;
  reg                 io_in_r_bypass_regNext_7_1_load_store_1;
  reg                 io_in_r_bypass_regNext_7_1_df_is_ws_1;
  reg                 io_in_r_bypass_regNext_7_1_stall_1;
  reg        [15:0]   io_in_r_bypass_regNext_7_2_data_1;
  reg                 io_in_r_bypass_regNext_7_2_load_store_1;
  reg                 io_in_r_bypass_regNext_7_2_df_is_ws_1;
  reg                 io_in_r_bypass_regNext_7_2_stall_1;
  reg        [15:0]   io_in_r_bypass_regNext_7_3_data_1;
  reg                 io_in_r_bypass_regNext_7_3_load_store_1;
  reg                 io_in_r_bypass_regNext_7_3_df_is_ws_1;
  reg                 io_in_r_bypass_regNext_7_3_stall_1;
  reg        [15:0]   io_in_r_bypass_regNext_8_0_data_1;
  reg                 io_in_r_bypass_regNext_8_0_load_store_1;
  reg                 io_in_r_bypass_regNext_8_0_df_is_ws_1;
  reg                 io_in_r_bypass_regNext_8_0_stall_1;
  reg        [15:0]   io_in_r_bypass_regNext_8_1_data_1;
  reg                 io_in_r_bypass_regNext_8_1_load_store_1;
  reg                 io_in_r_bypass_regNext_8_1_df_is_ws_1;
  reg                 io_in_r_bypass_regNext_8_1_stall_1;
  reg        [15:0]   io_in_r_bypass_regNext_8_2_data_1;
  reg                 io_in_r_bypass_regNext_8_2_load_store_1;
  reg                 io_in_r_bypass_regNext_8_2_df_is_ws_1;
  reg                 io_in_r_bypass_regNext_8_2_stall_1;
  reg        [15:0]   io_in_r_bypass_regNext_8_3_data_1;
  reg                 io_in_r_bypass_regNext_8_3_load_store_1;
  reg                 io_in_r_bypass_regNext_8_3_df_is_ws_1;
  reg                 io_in_r_bypass_regNext_8_3_stall_1;
  reg        [15:0]   io_in_r_bypass_regNext_9_0_data_1;
  reg                 io_in_r_bypass_regNext_9_0_load_store_1;
  reg                 io_in_r_bypass_regNext_9_0_df_is_ws_1;
  reg                 io_in_r_bypass_regNext_9_0_stall_1;
  reg        [15:0]   io_in_r_bypass_regNext_9_1_data_1;
  reg                 io_in_r_bypass_regNext_9_1_load_store_1;
  reg                 io_in_r_bypass_regNext_9_1_df_is_ws_1;
  reg                 io_in_r_bypass_regNext_9_1_stall_1;
  reg        [15:0]   io_in_r_bypass_regNext_9_2_data_1;
  reg                 io_in_r_bypass_regNext_9_2_load_store_1;
  reg                 io_in_r_bypass_regNext_9_2_df_is_ws_1;
  reg                 io_in_r_bypass_regNext_9_2_stall_1;
  reg        [15:0]   io_in_r_bypass_regNext_9_3_data_1;
  reg                 io_in_r_bypass_regNext_9_3_load_store_1;
  reg                 io_in_r_bypass_regNext_9_3_df_is_ws_1;
  reg                 io_in_r_bypass_regNext_9_3_stall_1;
  reg        [15:0]   io_in_r_bypass_regNext_10_0_data_1;
  reg                 io_in_r_bypass_regNext_10_0_load_store_1;
  reg                 io_in_r_bypass_regNext_10_0_df_is_ws_1;
  reg                 io_in_r_bypass_regNext_10_0_stall_1;
  reg        [15:0]   io_in_r_bypass_regNext_10_1_data_1;
  reg                 io_in_r_bypass_regNext_10_1_load_store_1;
  reg                 io_in_r_bypass_regNext_10_1_df_is_ws_1;
  reg                 io_in_r_bypass_regNext_10_1_stall_1;
  reg        [15:0]   io_in_r_bypass_regNext_10_2_data_1;
  reg                 io_in_r_bypass_regNext_10_2_load_store_1;
  reg                 io_in_r_bypass_regNext_10_2_df_is_ws_1;
  reg                 io_in_r_bypass_regNext_10_2_stall_1;
  reg        [15:0]   io_in_r_bypass_regNext_10_3_data_1;
  reg                 io_in_r_bypass_regNext_10_3_load_store_1;
  reg                 io_in_r_bypass_regNext_10_3_df_is_ws_1;
  reg                 io_in_r_bypass_regNext_10_3_stall_1;
  reg        [15:0]   io_in_r_bypass_regNext_11_0_data_1;
  reg                 io_in_r_bypass_regNext_11_0_load_store_1;
  reg                 io_in_r_bypass_regNext_11_0_df_is_ws_1;
  reg                 io_in_r_bypass_regNext_11_0_stall_1;
  reg        [15:0]   io_in_r_bypass_regNext_11_1_data_1;
  reg                 io_in_r_bypass_regNext_11_1_load_store_1;
  reg                 io_in_r_bypass_regNext_11_1_df_is_ws_1;
  reg                 io_in_r_bypass_regNext_11_1_stall_1;
  reg        [15:0]   io_in_r_bypass_regNext_11_2_data_1;
  reg                 io_in_r_bypass_regNext_11_2_load_store_1;
  reg                 io_in_r_bypass_regNext_11_2_df_is_ws_1;
  reg                 io_in_r_bypass_regNext_11_2_stall_1;
  reg        [15:0]   io_in_r_bypass_regNext_11_3_data_1;
  reg                 io_in_r_bypass_regNext_11_3_load_store_1;
  reg                 io_in_r_bypass_regNext_11_3_df_is_ws_1;
  reg                 io_in_r_bypass_regNext_11_3_stall_1;
  reg        [15:0]   io_in_r_bypass_regNext_12_0_data_1;
  reg                 io_in_r_bypass_regNext_12_0_load_store_1;
  reg                 io_in_r_bypass_regNext_12_0_df_is_ws_1;
  reg                 io_in_r_bypass_regNext_12_0_stall_1;
  reg        [15:0]   io_in_r_bypass_regNext_12_1_data_1;
  reg                 io_in_r_bypass_regNext_12_1_load_store_1;
  reg                 io_in_r_bypass_regNext_12_1_df_is_ws_1;
  reg                 io_in_r_bypass_regNext_12_1_stall_1;
  reg        [15:0]   io_in_r_bypass_regNext_12_2_data_1;
  reg                 io_in_r_bypass_regNext_12_2_load_store_1;
  reg                 io_in_r_bypass_regNext_12_2_df_is_ws_1;
  reg                 io_in_r_bypass_regNext_12_2_stall_1;
  reg        [15:0]   io_in_r_bypass_regNext_12_3_data_1;
  reg                 io_in_r_bypass_regNext_12_3_load_store_1;
  reg                 io_in_r_bypass_regNext_12_3_df_is_ws_1;
  reg                 io_in_r_bypass_regNext_12_3_stall_1;
  reg        [15:0]   io_in_r_bypass_regNext_13_0_data_1;
  reg                 io_in_r_bypass_regNext_13_0_load_store_1;
  reg                 io_in_r_bypass_regNext_13_0_df_is_ws_1;
  reg                 io_in_r_bypass_regNext_13_0_stall_1;
  reg        [15:0]   io_in_r_bypass_regNext_13_1_data_1;
  reg                 io_in_r_bypass_regNext_13_1_load_store_1;
  reg                 io_in_r_bypass_regNext_13_1_df_is_ws_1;
  reg                 io_in_r_bypass_regNext_13_1_stall_1;
  reg        [15:0]   io_in_r_bypass_regNext_13_2_data_1;
  reg                 io_in_r_bypass_regNext_13_2_load_store_1;
  reg                 io_in_r_bypass_regNext_13_2_df_is_ws_1;
  reg                 io_in_r_bypass_regNext_13_2_stall_1;
  reg        [15:0]   io_in_r_bypass_regNext_13_3_data_1;
  reg                 io_in_r_bypass_regNext_13_3_load_store_1;
  reg                 io_in_r_bypass_regNext_13_3_df_is_ws_1;
  reg                 io_in_r_bypass_regNext_13_3_stall_1;
  reg        [15:0]   io_in_r_bypass_regNext_14_0_data_1;
  reg                 io_in_r_bypass_regNext_14_0_load_store_1;
  reg                 io_in_r_bypass_regNext_14_0_df_is_ws_1;
  reg                 io_in_r_bypass_regNext_14_0_stall_1;
  reg        [15:0]   io_in_r_bypass_regNext_14_1_data_1;
  reg                 io_in_r_bypass_regNext_14_1_load_store_1;
  reg                 io_in_r_bypass_regNext_14_1_df_is_ws_1;
  reg                 io_in_r_bypass_regNext_14_1_stall_1;
  reg        [15:0]   io_in_r_bypass_regNext_14_2_data_1;
  reg                 io_in_r_bypass_regNext_14_2_load_store_1;
  reg                 io_in_r_bypass_regNext_14_2_df_is_ws_1;
  reg                 io_in_r_bypass_regNext_14_2_stall_1;
  reg        [15:0]   io_in_r_bypass_regNext_14_3_data_1;
  reg                 io_in_r_bypass_regNext_14_3_load_store_1;
  reg                 io_in_r_bypass_regNext_14_3_df_is_ws_1;
  reg                 io_in_r_bypass_regNext_14_3_stall_1;
  reg        [15:0]   io_in_r_bypass_regNext_15_0_data_1;
  reg                 io_in_r_bypass_regNext_15_0_load_store_1;
  reg                 io_in_r_bypass_regNext_15_0_df_is_ws_1;
  reg                 io_in_r_bypass_regNext_15_0_stall_1;
  reg        [15:0]   io_in_r_bypass_regNext_15_1_data_1;
  reg                 io_in_r_bypass_regNext_15_1_load_store_1;
  reg                 io_in_r_bypass_regNext_15_1_df_is_ws_1;
  reg                 io_in_r_bypass_regNext_15_1_stall_1;
  reg        [15:0]   io_in_r_bypass_regNext_15_2_data_1;
  reg                 io_in_r_bypass_regNext_15_2_load_store_1;
  reg                 io_in_r_bypass_regNext_15_2_df_is_ws_1;
  reg                 io_in_r_bypass_regNext_15_2_stall_1;
  reg        [15:0]   io_in_r_bypass_regNext_15_3_data_1;
  reg                 io_in_r_bypass_regNext_15_3_load_store_1;
  reg                 io_in_r_bypass_regNext_15_3_df_is_ws_1;
  reg                 io_in_r_bypass_regNext_15_3_stall_1;
  reg        [15:0]   io_in_r_bypass_regNext_16_0_data_1;
  reg                 io_in_r_bypass_regNext_16_0_load_store_1;
  reg                 io_in_r_bypass_regNext_16_0_df_is_ws_1;
  reg                 io_in_r_bypass_regNext_16_0_stall_1;
  reg        [15:0]   io_in_r_bypass_regNext_16_1_data_1;
  reg                 io_in_r_bypass_regNext_16_1_load_store_1;
  reg                 io_in_r_bypass_regNext_16_1_df_is_ws_1;
  reg                 io_in_r_bypass_regNext_16_1_stall_1;
  reg        [15:0]   io_in_r_bypass_regNext_16_2_data_1;
  reg                 io_in_r_bypass_regNext_16_2_load_store_1;
  reg                 io_in_r_bypass_regNext_16_2_df_is_ws_1;
  reg                 io_in_r_bypass_regNext_16_2_stall_1;
  reg        [15:0]   io_in_r_bypass_regNext_16_3_data_1;
  reg                 io_in_r_bypass_regNext_16_3_load_store_1;
  reg                 io_in_r_bypass_regNext_16_3_df_is_ws_1;
  reg                 io_in_r_bypass_regNext_16_3_stall_1;
  reg        [15:0]   io_in_r_bypass_regNext_17_0_data_1;
  reg                 io_in_r_bypass_regNext_17_0_load_store_1;
  reg                 io_in_r_bypass_regNext_17_0_df_is_ws_1;
  reg                 io_in_r_bypass_regNext_17_0_stall_1;
  reg        [15:0]   io_in_r_bypass_regNext_17_1_data_1;
  reg                 io_in_r_bypass_regNext_17_1_load_store_1;
  reg                 io_in_r_bypass_regNext_17_1_df_is_ws_1;
  reg                 io_in_r_bypass_regNext_17_1_stall_1;
  reg        [15:0]   io_in_r_bypass_regNext_17_2_data_1;
  reg                 io_in_r_bypass_regNext_17_2_load_store_1;
  reg                 io_in_r_bypass_regNext_17_2_df_is_ws_1;
  reg                 io_in_r_bypass_regNext_17_2_stall_1;
  reg        [15:0]   io_in_r_bypass_regNext_17_3_data_1;
  reg                 io_in_r_bypass_regNext_17_3_load_store_1;
  reg                 io_in_r_bypass_regNext_17_3_df_is_ws_1;
  reg                 io_in_r_bypass_regNext_17_3_stall_1;
  reg        [15:0]   io_in_r_bypass_regNext_18_0_data_1;
  reg                 io_in_r_bypass_regNext_18_0_load_store_1;
  reg                 io_in_r_bypass_regNext_18_0_df_is_ws_1;
  reg                 io_in_r_bypass_regNext_18_0_stall_1;
  reg        [15:0]   io_in_r_bypass_regNext_18_1_data_1;
  reg                 io_in_r_bypass_regNext_18_1_load_store_1;
  reg                 io_in_r_bypass_regNext_18_1_df_is_ws_1;
  reg                 io_in_r_bypass_regNext_18_1_stall_1;
  reg        [15:0]   io_in_r_bypass_regNext_18_2_data_1;
  reg                 io_in_r_bypass_regNext_18_2_load_store_1;
  reg                 io_in_r_bypass_regNext_18_2_df_is_ws_1;
  reg                 io_in_r_bypass_regNext_18_2_stall_1;
  reg        [15:0]   io_in_r_bypass_regNext_18_3_data_1;
  reg                 io_in_r_bypass_regNext_18_3_load_store_1;
  reg                 io_in_r_bypass_regNext_18_3_df_is_ws_1;
  reg                 io_in_r_bypass_regNext_18_3_stall_1;
  reg        [15:0]   io_in_r_bypass_regNext_19_0_data_1;
  reg                 io_in_r_bypass_regNext_19_0_load_store_1;
  reg                 io_in_r_bypass_regNext_19_0_df_is_ws_1;
  reg                 io_in_r_bypass_regNext_19_0_stall_1;
  reg        [15:0]   io_in_r_bypass_regNext_19_1_data_1;
  reg                 io_in_r_bypass_regNext_19_1_load_store_1;
  reg                 io_in_r_bypass_regNext_19_1_df_is_ws_1;
  reg                 io_in_r_bypass_regNext_19_1_stall_1;
  reg        [15:0]   io_in_r_bypass_regNext_19_2_data_1;
  reg                 io_in_r_bypass_regNext_19_2_load_store_1;
  reg                 io_in_r_bypass_regNext_19_2_df_is_ws_1;
  reg                 io_in_r_bypass_regNext_19_2_stall_1;
  reg        [15:0]   io_in_r_bypass_regNext_19_3_data_1;
  reg                 io_in_r_bypass_regNext_19_3_load_store_1;
  reg                 io_in_r_bypass_regNext_19_3_df_is_ws_1;
  reg                 io_in_r_bypass_regNext_19_3_stall_1;
  reg        [15:0]   io_in_r_bypass_regNext_20_0_data_1;
  reg                 io_in_r_bypass_regNext_20_0_load_store_1;
  reg                 io_in_r_bypass_regNext_20_0_df_is_ws_1;
  reg                 io_in_r_bypass_regNext_20_0_stall_1;
  reg        [15:0]   io_in_r_bypass_regNext_20_1_data_1;
  reg                 io_in_r_bypass_regNext_20_1_load_store_1;
  reg                 io_in_r_bypass_regNext_20_1_df_is_ws_1;
  reg                 io_in_r_bypass_regNext_20_1_stall_1;
  reg        [15:0]   io_in_r_bypass_regNext_20_2_data_1;
  reg                 io_in_r_bypass_regNext_20_2_load_store_1;
  reg                 io_in_r_bypass_regNext_20_2_df_is_ws_1;
  reg                 io_in_r_bypass_regNext_20_2_stall_1;
  reg        [15:0]   io_in_r_bypass_regNext_20_3_data_1;
  reg                 io_in_r_bypass_regNext_20_3_load_store_1;
  reg                 io_in_r_bypass_regNext_20_3_df_is_ws_1;
  reg                 io_in_r_bypass_regNext_20_3_stall_1;
  reg        [15:0]   io_in_r_bypass_regNext_21_0_data_1;
  reg                 io_in_r_bypass_regNext_21_0_load_store_1;
  reg                 io_in_r_bypass_regNext_21_0_df_is_ws_1;
  reg                 io_in_r_bypass_regNext_21_0_stall_1;
  reg        [15:0]   io_in_r_bypass_regNext_21_1_data_1;
  reg                 io_in_r_bypass_regNext_21_1_load_store_1;
  reg                 io_in_r_bypass_regNext_21_1_df_is_ws_1;
  reg                 io_in_r_bypass_regNext_21_1_stall_1;
  reg        [15:0]   io_in_r_bypass_regNext_21_2_data_1;
  reg                 io_in_r_bypass_regNext_21_2_load_store_1;
  reg                 io_in_r_bypass_regNext_21_2_df_is_ws_1;
  reg                 io_in_r_bypass_regNext_21_2_stall_1;
  reg        [15:0]   io_in_r_bypass_regNext_21_3_data_1;
  reg                 io_in_r_bypass_regNext_21_3_load_store_1;
  reg                 io_in_r_bypass_regNext_21_3_df_is_ws_1;
  reg                 io_in_r_bypass_regNext_21_3_stall_1;
  reg        [15:0]   io_in_r_bypass_regNext_22_0_data_1;
  reg                 io_in_r_bypass_regNext_22_0_load_store_1;
  reg                 io_in_r_bypass_regNext_22_0_df_is_ws_1;
  reg                 io_in_r_bypass_regNext_22_0_stall_1;
  reg        [15:0]   io_in_r_bypass_regNext_22_1_data_1;
  reg                 io_in_r_bypass_regNext_22_1_load_store_1;
  reg                 io_in_r_bypass_regNext_22_1_df_is_ws_1;
  reg                 io_in_r_bypass_regNext_22_1_stall_1;
  reg        [15:0]   io_in_r_bypass_regNext_22_2_data_1;
  reg                 io_in_r_bypass_regNext_22_2_load_store_1;
  reg                 io_in_r_bypass_regNext_22_2_df_is_ws_1;
  reg                 io_in_r_bypass_regNext_22_2_stall_1;
  reg        [15:0]   io_in_r_bypass_regNext_22_3_data_1;
  reg                 io_in_r_bypass_regNext_22_3_load_store_1;
  reg                 io_in_r_bypass_regNext_22_3_df_is_ws_1;
  reg                 io_in_r_bypass_regNext_22_3_stall_1;
  reg        [15:0]   io_in_r_bypass_regNext_23_0_data_1;
  reg                 io_in_r_bypass_regNext_23_0_load_store_1;
  reg                 io_in_r_bypass_regNext_23_0_df_is_ws_1;
  reg                 io_in_r_bypass_regNext_23_0_stall_1;
  reg        [15:0]   io_in_r_bypass_regNext_23_1_data_1;
  reg                 io_in_r_bypass_regNext_23_1_load_store_1;
  reg                 io_in_r_bypass_regNext_23_1_df_is_ws_1;
  reg                 io_in_r_bypass_regNext_23_1_stall_1;
  reg        [15:0]   io_in_r_bypass_regNext_23_2_data_1;
  reg                 io_in_r_bypass_regNext_23_2_load_store_1;
  reg                 io_in_r_bypass_regNext_23_2_df_is_ws_1;
  reg                 io_in_r_bypass_regNext_23_2_stall_1;
  reg        [15:0]   io_in_r_bypass_regNext_23_3_data_1;
  reg                 io_in_r_bypass_regNext_23_3_load_store_1;
  reg                 io_in_r_bypass_regNext_23_3_df_is_ws_1;
  reg                 io_in_r_bypass_regNext_23_3_stall_1;
  reg        [15:0]   io_in_r_bypass_regNext_24_0_data_1;
  reg                 io_in_r_bypass_regNext_24_0_load_store_1;
  reg                 io_in_r_bypass_regNext_24_0_df_is_ws_1;
  reg                 io_in_r_bypass_regNext_24_0_stall_1;
  reg        [15:0]   io_in_r_bypass_regNext_24_1_data_1;
  reg                 io_in_r_bypass_regNext_24_1_load_store_1;
  reg                 io_in_r_bypass_regNext_24_1_df_is_ws_1;
  reg                 io_in_r_bypass_regNext_24_1_stall_1;
  reg        [15:0]   io_in_r_bypass_regNext_24_2_data_1;
  reg                 io_in_r_bypass_regNext_24_2_load_store_1;
  reg                 io_in_r_bypass_regNext_24_2_df_is_ws_1;
  reg                 io_in_r_bypass_regNext_24_2_stall_1;
  reg        [15:0]   io_in_r_bypass_regNext_24_3_data_1;
  reg                 io_in_r_bypass_regNext_24_3_load_store_1;
  reg                 io_in_r_bypass_regNext_24_3_df_is_ws_1;
  reg                 io_in_r_bypass_regNext_24_3_stall_1;
  reg        [15:0]   io_in_r_bypass_regNext_25_0_data_1;
  reg                 io_in_r_bypass_regNext_25_0_load_store_1;
  reg                 io_in_r_bypass_regNext_25_0_df_is_ws_1;
  reg                 io_in_r_bypass_regNext_25_0_stall_1;
  reg        [15:0]   io_in_r_bypass_regNext_25_1_data_1;
  reg                 io_in_r_bypass_regNext_25_1_load_store_1;
  reg                 io_in_r_bypass_regNext_25_1_df_is_ws_1;
  reg                 io_in_r_bypass_regNext_25_1_stall_1;
  reg        [15:0]   io_in_r_bypass_regNext_25_2_data_1;
  reg                 io_in_r_bypass_regNext_25_2_load_store_1;
  reg                 io_in_r_bypass_regNext_25_2_df_is_ws_1;
  reg                 io_in_r_bypass_regNext_25_2_stall_1;
  reg        [15:0]   io_in_r_bypass_regNext_25_3_data_1;
  reg                 io_in_r_bypass_regNext_25_3_load_store_1;
  reg                 io_in_r_bypass_regNext_25_3_df_is_ws_1;
  reg                 io_in_r_bypass_regNext_25_3_stall_1;
  reg        [15:0]   io_in_r_bypass_regNext_26_0_data_1;
  reg                 io_in_r_bypass_regNext_26_0_load_store_1;
  reg                 io_in_r_bypass_regNext_26_0_df_is_ws_1;
  reg                 io_in_r_bypass_regNext_26_0_stall_1;
  reg        [15:0]   io_in_r_bypass_regNext_26_1_data_1;
  reg                 io_in_r_bypass_regNext_26_1_load_store_1;
  reg                 io_in_r_bypass_regNext_26_1_df_is_ws_1;
  reg                 io_in_r_bypass_regNext_26_1_stall_1;
  reg        [15:0]   io_in_r_bypass_regNext_26_2_data_1;
  reg                 io_in_r_bypass_regNext_26_2_load_store_1;
  reg                 io_in_r_bypass_regNext_26_2_df_is_ws_1;
  reg                 io_in_r_bypass_regNext_26_2_stall_1;
  reg        [15:0]   io_in_r_bypass_regNext_26_3_data_1;
  reg                 io_in_r_bypass_regNext_26_3_load_store_1;
  reg                 io_in_r_bypass_regNext_26_3_df_is_ws_1;
  reg                 io_in_r_bypass_regNext_26_3_stall_1;
  reg        [15:0]   io_in_r_bypass_regNext_27_0_data_1;
  reg                 io_in_r_bypass_regNext_27_0_load_store_1;
  reg                 io_in_r_bypass_regNext_27_0_df_is_ws_1;
  reg                 io_in_r_bypass_regNext_27_0_stall_1;
  reg        [15:0]   io_in_r_bypass_regNext_27_1_data_1;
  reg                 io_in_r_bypass_regNext_27_1_load_store_1;
  reg                 io_in_r_bypass_regNext_27_1_df_is_ws_1;
  reg                 io_in_r_bypass_regNext_27_1_stall_1;
  reg        [15:0]   io_in_r_bypass_regNext_27_2_data_1;
  reg                 io_in_r_bypass_regNext_27_2_load_store_1;
  reg                 io_in_r_bypass_regNext_27_2_df_is_ws_1;
  reg                 io_in_r_bypass_regNext_27_2_stall_1;
  reg        [15:0]   io_in_r_bypass_regNext_27_3_data_1;
  reg                 io_in_r_bypass_regNext_27_3_load_store_1;
  reg                 io_in_r_bypass_regNext_27_3_df_is_ws_1;
  reg                 io_in_r_bypass_regNext_27_3_stall_1;
  reg        [15:0]   io_in_r_bypass_regNext_28_0_data_1;
  reg                 io_in_r_bypass_regNext_28_0_load_store_1;
  reg                 io_in_r_bypass_regNext_28_0_df_is_ws_1;
  reg                 io_in_r_bypass_regNext_28_0_stall_1;
  reg        [15:0]   io_in_r_bypass_regNext_28_1_data_1;
  reg                 io_in_r_bypass_regNext_28_1_load_store_1;
  reg                 io_in_r_bypass_regNext_28_1_df_is_ws_1;
  reg                 io_in_r_bypass_regNext_28_1_stall_1;
  reg        [15:0]   io_in_r_bypass_regNext_28_2_data_1;
  reg                 io_in_r_bypass_regNext_28_2_load_store_1;
  reg                 io_in_r_bypass_regNext_28_2_df_is_ws_1;
  reg                 io_in_r_bypass_regNext_28_2_stall_1;
  reg        [15:0]   io_in_r_bypass_regNext_28_3_data_1;
  reg                 io_in_r_bypass_regNext_28_3_load_store_1;
  reg                 io_in_r_bypass_regNext_28_3_df_is_ws_1;
  reg                 io_in_r_bypass_regNext_28_3_stall_1;
  reg        [15:0]   io_in_r_bypass_regNext_29_0_data_1;
  reg                 io_in_r_bypass_regNext_29_0_load_store_1;
  reg                 io_in_r_bypass_regNext_29_0_df_is_ws_1;
  reg                 io_in_r_bypass_regNext_29_0_stall_1;
  reg        [15:0]   io_in_r_bypass_regNext_29_1_data_1;
  reg                 io_in_r_bypass_regNext_29_1_load_store_1;
  reg                 io_in_r_bypass_regNext_29_1_df_is_ws_1;
  reg                 io_in_r_bypass_regNext_29_1_stall_1;
  reg        [15:0]   io_in_r_bypass_regNext_29_2_data_1;
  reg                 io_in_r_bypass_regNext_29_2_load_store_1;
  reg                 io_in_r_bypass_regNext_29_2_df_is_ws_1;
  reg                 io_in_r_bypass_regNext_29_2_stall_1;
  reg        [15:0]   io_in_r_bypass_regNext_29_3_data_1;
  reg                 io_in_r_bypass_regNext_29_3_load_store_1;
  reg                 io_in_r_bypass_regNext_29_3_df_is_ws_1;
  reg                 io_in_r_bypass_regNext_29_3_stall_1;
  reg        [15:0]   io_in_r_bypass_regNext_30_0_data_1;
  reg                 io_in_r_bypass_regNext_30_0_load_store_1;
  reg                 io_in_r_bypass_regNext_30_0_df_is_ws_1;
  reg                 io_in_r_bypass_regNext_30_0_stall_1;
  reg        [15:0]   io_in_r_bypass_regNext_30_1_data_1;
  reg                 io_in_r_bypass_regNext_30_1_load_store_1;
  reg                 io_in_r_bypass_regNext_30_1_df_is_ws_1;
  reg                 io_in_r_bypass_regNext_30_1_stall_1;
  reg        [15:0]   io_in_r_bypass_regNext_30_2_data_1;
  reg                 io_in_r_bypass_regNext_30_2_load_store_1;
  reg                 io_in_r_bypass_regNext_30_2_df_is_ws_1;
  reg                 io_in_r_bypass_regNext_30_2_stall_1;
  reg        [15:0]   io_in_r_bypass_regNext_30_3_data_1;
  reg                 io_in_r_bypass_regNext_30_3_load_store_1;
  reg                 io_in_r_bypass_regNext_30_3_df_is_ws_1;
  reg                 io_in_r_bypass_regNext_30_3_stall_1;
  reg        [15:0]   io_in_r_bypass_regNext_31_0_data_1;
  reg                 io_in_r_bypass_regNext_31_0_load_store_1;
  reg                 io_in_r_bypass_regNext_31_0_df_is_ws_1;
  reg                 io_in_r_bypass_regNext_31_0_stall_1;
  reg        [15:0]   io_in_r_bypass_regNext_31_1_data_1;
  reg                 io_in_r_bypass_regNext_31_1_load_store_1;
  reg                 io_in_r_bypass_regNext_31_1_df_is_ws_1;
  reg                 io_in_r_bypass_regNext_31_1_stall_1;
  reg        [15:0]   io_in_r_bypass_regNext_31_2_data_1;
  reg                 io_in_r_bypass_regNext_31_2_load_store_1;
  reg                 io_in_r_bypass_regNext_31_2_df_is_ws_1;
  reg                 io_in_r_bypass_regNext_31_2_stall_1;
  reg        [15:0]   io_in_r_bypass_regNext_31_3_data_1;
  reg                 io_in_r_bypass_regNext_31_3_load_store_1;
  reg                 io_in_r_bypass_regNext_31_3_df_is_ws_1;
  reg                 io_in_r_bypass_regNext_31_3_stall_1;
  reg        [15:0]   io_in_r_bypass_regNext_0_0_data_2;
  reg                 io_in_r_bypass_regNext_0_0_load_store_2;
  reg                 io_in_r_bypass_regNext_0_0_df_is_ws_2;
  reg                 io_in_r_bypass_regNext_0_0_stall_2;
  reg        [15:0]   io_in_r_bypass_regNext_0_1_data_2;
  reg                 io_in_r_bypass_regNext_0_1_load_store_2;
  reg                 io_in_r_bypass_regNext_0_1_df_is_ws_2;
  reg                 io_in_r_bypass_regNext_0_1_stall_2;
  reg        [15:0]   io_in_r_bypass_regNext_0_2_data_2;
  reg                 io_in_r_bypass_regNext_0_2_load_store_2;
  reg                 io_in_r_bypass_regNext_0_2_df_is_ws_2;
  reg                 io_in_r_bypass_regNext_0_2_stall_2;
  reg        [15:0]   io_in_r_bypass_regNext_0_3_data_2;
  reg                 io_in_r_bypass_regNext_0_3_load_store_2;
  reg                 io_in_r_bypass_regNext_0_3_df_is_ws_2;
  reg                 io_in_r_bypass_regNext_0_3_stall_2;
  reg        [15:0]   io_in_r_bypass_regNext_1_0_data_2;
  reg                 io_in_r_bypass_regNext_1_0_load_store_2;
  reg                 io_in_r_bypass_regNext_1_0_df_is_ws_2;
  reg                 io_in_r_bypass_regNext_1_0_stall_2;
  reg        [15:0]   io_in_r_bypass_regNext_1_1_data_2;
  reg                 io_in_r_bypass_regNext_1_1_load_store_2;
  reg                 io_in_r_bypass_regNext_1_1_df_is_ws_2;
  reg                 io_in_r_bypass_regNext_1_1_stall_2;
  reg        [15:0]   io_in_r_bypass_regNext_1_2_data_2;
  reg                 io_in_r_bypass_regNext_1_2_load_store_2;
  reg                 io_in_r_bypass_regNext_1_2_df_is_ws_2;
  reg                 io_in_r_bypass_regNext_1_2_stall_2;
  reg        [15:0]   io_in_r_bypass_regNext_1_3_data_2;
  reg                 io_in_r_bypass_regNext_1_3_load_store_2;
  reg                 io_in_r_bypass_regNext_1_3_df_is_ws_2;
  reg                 io_in_r_bypass_regNext_1_3_stall_2;
  reg        [15:0]   io_in_r_bypass_regNext_2_0_data_2;
  reg                 io_in_r_bypass_regNext_2_0_load_store_2;
  reg                 io_in_r_bypass_regNext_2_0_df_is_ws_2;
  reg                 io_in_r_bypass_regNext_2_0_stall_2;
  reg        [15:0]   io_in_r_bypass_regNext_2_1_data_2;
  reg                 io_in_r_bypass_regNext_2_1_load_store_2;
  reg                 io_in_r_bypass_regNext_2_1_df_is_ws_2;
  reg                 io_in_r_bypass_regNext_2_1_stall_2;
  reg        [15:0]   io_in_r_bypass_regNext_2_2_data_2;
  reg                 io_in_r_bypass_regNext_2_2_load_store_2;
  reg                 io_in_r_bypass_regNext_2_2_df_is_ws_2;
  reg                 io_in_r_bypass_regNext_2_2_stall_2;
  reg        [15:0]   io_in_r_bypass_regNext_2_3_data_2;
  reg                 io_in_r_bypass_regNext_2_3_load_store_2;
  reg                 io_in_r_bypass_regNext_2_3_df_is_ws_2;
  reg                 io_in_r_bypass_regNext_2_3_stall_2;
  reg        [15:0]   io_in_r_bypass_regNext_3_0_data_2;
  reg                 io_in_r_bypass_regNext_3_0_load_store_2;
  reg                 io_in_r_bypass_regNext_3_0_df_is_ws_2;
  reg                 io_in_r_bypass_regNext_3_0_stall_2;
  reg        [15:0]   io_in_r_bypass_regNext_3_1_data_2;
  reg                 io_in_r_bypass_regNext_3_1_load_store_2;
  reg                 io_in_r_bypass_regNext_3_1_df_is_ws_2;
  reg                 io_in_r_bypass_regNext_3_1_stall_2;
  reg        [15:0]   io_in_r_bypass_regNext_3_2_data_2;
  reg                 io_in_r_bypass_regNext_3_2_load_store_2;
  reg                 io_in_r_bypass_regNext_3_2_df_is_ws_2;
  reg                 io_in_r_bypass_regNext_3_2_stall_2;
  reg        [15:0]   io_in_r_bypass_regNext_3_3_data_2;
  reg                 io_in_r_bypass_regNext_3_3_load_store_2;
  reg                 io_in_r_bypass_regNext_3_3_df_is_ws_2;
  reg                 io_in_r_bypass_regNext_3_3_stall_2;
  reg        [15:0]   io_in_r_bypass_regNext_4_0_data_2;
  reg                 io_in_r_bypass_regNext_4_0_load_store_2;
  reg                 io_in_r_bypass_regNext_4_0_df_is_ws_2;
  reg                 io_in_r_bypass_regNext_4_0_stall_2;
  reg        [15:0]   io_in_r_bypass_regNext_4_1_data_2;
  reg                 io_in_r_bypass_regNext_4_1_load_store_2;
  reg                 io_in_r_bypass_regNext_4_1_df_is_ws_2;
  reg                 io_in_r_bypass_regNext_4_1_stall_2;
  reg        [15:0]   io_in_r_bypass_regNext_4_2_data_2;
  reg                 io_in_r_bypass_regNext_4_2_load_store_2;
  reg                 io_in_r_bypass_regNext_4_2_df_is_ws_2;
  reg                 io_in_r_bypass_regNext_4_2_stall_2;
  reg        [15:0]   io_in_r_bypass_regNext_4_3_data_2;
  reg                 io_in_r_bypass_regNext_4_3_load_store_2;
  reg                 io_in_r_bypass_regNext_4_3_df_is_ws_2;
  reg                 io_in_r_bypass_regNext_4_3_stall_2;
  reg        [15:0]   io_in_r_bypass_regNext_5_0_data_2;
  reg                 io_in_r_bypass_regNext_5_0_load_store_2;
  reg                 io_in_r_bypass_regNext_5_0_df_is_ws_2;
  reg                 io_in_r_bypass_regNext_5_0_stall_2;
  reg        [15:0]   io_in_r_bypass_regNext_5_1_data_2;
  reg                 io_in_r_bypass_regNext_5_1_load_store_2;
  reg                 io_in_r_bypass_regNext_5_1_df_is_ws_2;
  reg                 io_in_r_bypass_regNext_5_1_stall_2;
  reg        [15:0]   io_in_r_bypass_regNext_5_2_data_2;
  reg                 io_in_r_bypass_regNext_5_2_load_store_2;
  reg                 io_in_r_bypass_regNext_5_2_df_is_ws_2;
  reg                 io_in_r_bypass_regNext_5_2_stall_2;
  reg        [15:0]   io_in_r_bypass_regNext_5_3_data_2;
  reg                 io_in_r_bypass_regNext_5_3_load_store_2;
  reg                 io_in_r_bypass_regNext_5_3_df_is_ws_2;
  reg                 io_in_r_bypass_regNext_5_3_stall_2;
  reg        [15:0]   io_in_r_bypass_regNext_6_0_data_2;
  reg                 io_in_r_bypass_regNext_6_0_load_store_2;
  reg                 io_in_r_bypass_regNext_6_0_df_is_ws_2;
  reg                 io_in_r_bypass_regNext_6_0_stall_2;
  reg        [15:0]   io_in_r_bypass_regNext_6_1_data_2;
  reg                 io_in_r_bypass_regNext_6_1_load_store_2;
  reg                 io_in_r_bypass_regNext_6_1_df_is_ws_2;
  reg                 io_in_r_bypass_regNext_6_1_stall_2;
  reg        [15:0]   io_in_r_bypass_regNext_6_2_data_2;
  reg                 io_in_r_bypass_regNext_6_2_load_store_2;
  reg                 io_in_r_bypass_regNext_6_2_df_is_ws_2;
  reg                 io_in_r_bypass_regNext_6_2_stall_2;
  reg        [15:0]   io_in_r_bypass_regNext_6_3_data_2;
  reg                 io_in_r_bypass_regNext_6_3_load_store_2;
  reg                 io_in_r_bypass_regNext_6_3_df_is_ws_2;
  reg                 io_in_r_bypass_regNext_6_3_stall_2;
  reg        [15:0]   io_in_r_bypass_regNext_7_0_data_2;
  reg                 io_in_r_bypass_regNext_7_0_load_store_2;
  reg                 io_in_r_bypass_regNext_7_0_df_is_ws_2;
  reg                 io_in_r_bypass_regNext_7_0_stall_2;
  reg        [15:0]   io_in_r_bypass_regNext_7_1_data_2;
  reg                 io_in_r_bypass_regNext_7_1_load_store_2;
  reg                 io_in_r_bypass_regNext_7_1_df_is_ws_2;
  reg                 io_in_r_bypass_regNext_7_1_stall_2;
  reg        [15:0]   io_in_r_bypass_regNext_7_2_data_2;
  reg                 io_in_r_bypass_regNext_7_2_load_store_2;
  reg                 io_in_r_bypass_regNext_7_2_df_is_ws_2;
  reg                 io_in_r_bypass_regNext_7_2_stall_2;
  reg        [15:0]   io_in_r_bypass_regNext_7_3_data_2;
  reg                 io_in_r_bypass_regNext_7_3_load_store_2;
  reg                 io_in_r_bypass_regNext_7_3_df_is_ws_2;
  reg                 io_in_r_bypass_regNext_7_3_stall_2;
  reg        [15:0]   io_in_r_bypass_regNext_8_0_data_2;
  reg                 io_in_r_bypass_regNext_8_0_load_store_2;
  reg                 io_in_r_bypass_regNext_8_0_df_is_ws_2;
  reg                 io_in_r_bypass_regNext_8_0_stall_2;
  reg        [15:0]   io_in_r_bypass_regNext_8_1_data_2;
  reg                 io_in_r_bypass_regNext_8_1_load_store_2;
  reg                 io_in_r_bypass_regNext_8_1_df_is_ws_2;
  reg                 io_in_r_bypass_regNext_8_1_stall_2;
  reg        [15:0]   io_in_r_bypass_regNext_8_2_data_2;
  reg                 io_in_r_bypass_regNext_8_2_load_store_2;
  reg                 io_in_r_bypass_regNext_8_2_df_is_ws_2;
  reg                 io_in_r_bypass_regNext_8_2_stall_2;
  reg        [15:0]   io_in_r_bypass_regNext_8_3_data_2;
  reg                 io_in_r_bypass_regNext_8_3_load_store_2;
  reg                 io_in_r_bypass_regNext_8_3_df_is_ws_2;
  reg                 io_in_r_bypass_regNext_8_3_stall_2;
  reg        [15:0]   io_in_r_bypass_regNext_9_0_data_2;
  reg                 io_in_r_bypass_regNext_9_0_load_store_2;
  reg                 io_in_r_bypass_regNext_9_0_df_is_ws_2;
  reg                 io_in_r_bypass_regNext_9_0_stall_2;
  reg        [15:0]   io_in_r_bypass_regNext_9_1_data_2;
  reg                 io_in_r_bypass_regNext_9_1_load_store_2;
  reg                 io_in_r_bypass_regNext_9_1_df_is_ws_2;
  reg                 io_in_r_bypass_regNext_9_1_stall_2;
  reg        [15:0]   io_in_r_bypass_regNext_9_2_data_2;
  reg                 io_in_r_bypass_regNext_9_2_load_store_2;
  reg                 io_in_r_bypass_regNext_9_2_df_is_ws_2;
  reg                 io_in_r_bypass_regNext_9_2_stall_2;
  reg        [15:0]   io_in_r_bypass_regNext_9_3_data_2;
  reg                 io_in_r_bypass_regNext_9_3_load_store_2;
  reg                 io_in_r_bypass_regNext_9_3_df_is_ws_2;
  reg                 io_in_r_bypass_regNext_9_3_stall_2;
  reg        [15:0]   io_in_r_bypass_regNext_10_0_data_2;
  reg                 io_in_r_bypass_regNext_10_0_load_store_2;
  reg                 io_in_r_bypass_regNext_10_0_df_is_ws_2;
  reg                 io_in_r_bypass_regNext_10_0_stall_2;
  reg        [15:0]   io_in_r_bypass_regNext_10_1_data_2;
  reg                 io_in_r_bypass_regNext_10_1_load_store_2;
  reg                 io_in_r_bypass_regNext_10_1_df_is_ws_2;
  reg                 io_in_r_bypass_regNext_10_1_stall_2;
  reg        [15:0]   io_in_r_bypass_regNext_10_2_data_2;
  reg                 io_in_r_bypass_regNext_10_2_load_store_2;
  reg                 io_in_r_bypass_regNext_10_2_df_is_ws_2;
  reg                 io_in_r_bypass_regNext_10_2_stall_2;
  reg        [15:0]   io_in_r_bypass_regNext_10_3_data_2;
  reg                 io_in_r_bypass_regNext_10_3_load_store_2;
  reg                 io_in_r_bypass_regNext_10_3_df_is_ws_2;
  reg                 io_in_r_bypass_regNext_10_3_stall_2;
  reg        [15:0]   io_in_r_bypass_regNext_11_0_data_2;
  reg                 io_in_r_bypass_regNext_11_0_load_store_2;
  reg                 io_in_r_bypass_regNext_11_0_df_is_ws_2;
  reg                 io_in_r_bypass_regNext_11_0_stall_2;
  reg        [15:0]   io_in_r_bypass_regNext_11_1_data_2;
  reg                 io_in_r_bypass_regNext_11_1_load_store_2;
  reg                 io_in_r_bypass_regNext_11_1_df_is_ws_2;
  reg                 io_in_r_bypass_regNext_11_1_stall_2;
  reg        [15:0]   io_in_r_bypass_regNext_11_2_data_2;
  reg                 io_in_r_bypass_regNext_11_2_load_store_2;
  reg                 io_in_r_bypass_regNext_11_2_df_is_ws_2;
  reg                 io_in_r_bypass_regNext_11_2_stall_2;
  reg        [15:0]   io_in_r_bypass_regNext_11_3_data_2;
  reg                 io_in_r_bypass_regNext_11_3_load_store_2;
  reg                 io_in_r_bypass_regNext_11_3_df_is_ws_2;
  reg                 io_in_r_bypass_regNext_11_3_stall_2;
  reg        [15:0]   io_in_r_bypass_regNext_12_0_data_2;
  reg                 io_in_r_bypass_regNext_12_0_load_store_2;
  reg                 io_in_r_bypass_regNext_12_0_df_is_ws_2;
  reg                 io_in_r_bypass_regNext_12_0_stall_2;
  reg        [15:0]   io_in_r_bypass_regNext_12_1_data_2;
  reg                 io_in_r_bypass_regNext_12_1_load_store_2;
  reg                 io_in_r_bypass_regNext_12_1_df_is_ws_2;
  reg                 io_in_r_bypass_regNext_12_1_stall_2;
  reg        [15:0]   io_in_r_bypass_regNext_12_2_data_2;
  reg                 io_in_r_bypass_regNext_12_2_load_store_2;
  reg                 io_in_r_bypass_regNext_12_2_df_is_ws_2;
  reg                 io_in_r_bypass_regNext_12_2_stall_2;
  reg        [15:0]   io_in_r_bypass_regNext_12_3_data_2;
  reg                 io_in_r_bypass_regNext_12_3_load_store_2;
  reg                 io_in_r_bypass_regNext_12_3_df_is_ws_2;
  reg                 io_in_r_bypass_regNext_12_3_stall_2;
  reg        [15:0]   io_in_r_bypass_regNext_13_0_data_2;
  reg                 io_in_r_bypass_regNext_13_0_load_store_2;
  reg                 io_in_r_bypass_regNext_13_0_df_is_ws_2;
  reg                 io_in_r_bypass_regNext_13_0_stall_2;
  reg        [15:0]   io_in_r_bypass_regNext_13_1_data_2;
  reg                 io_in_r_bypass_regNext_13_1_load_store_2;
  reg                 io_in_r_bypass_regNext_13_1_df_is_ws_2;
  reg                 io_in_r_bypass_regNext_13_1_stall_2;
  reg        [15:0]   io_in_r_bypass_regNext_13_2_data_2;
  reg                 io_in_r_bypass_regNext_13_2_load_store_2;
  reg                 io_in_r_bypass_regNext_13_2_df_is_ws_2;
  reg                 io_in_r_bypass_regNext_13_2_stall_2;
  reg        [15:0]   io_in_r_bypass_regNext_13_3_data_2;
  reg                 io_in_r_bypass_regNext_13_3_load_store_2;
  reg                 io_in_r_bypass_regNext_13_3_df_is_ws_2;
  reg                 io_in_r_bypass_regNext_13_3_stall_2;
  reg        [15:0]   io_in_r_bypass_regNext_14_0_data_2;
  reg                 io_in_r_bypass_regNext_14_0_load_store_2;
  reg                 io_in_r_bypass_regNext_14_0_df_is_ws_2;
  reg                 io_in_r_bypass_regNext_14_0_stall_2;
  reg        [15:0]   io_in_r_bypass_regNext_14_1_data_2;
  reg                 io_in_r_bypass_regNext_14_1_load_store_2;
  reg                 io_in_r_bypass_regNext_14_1_df_is_ws_2;
  reg                 io_in_r_bypass_regNext_14_1_stall_2;
  reg        [15:0]   io_in_r_bypass_regNext_14_2_data_2;
  reg                 io_in_r_bypass_regNext_14_2_load_store_2;
  reg                 io_in_r_bypass_regNext_14_2_df_is_ws_2;
  reg                 io_in_r_bypass_regNext_14_2_stall_2;
  reg        [15:0]   io_in_r_bypass_regNext_14_3_data_2;
  reg                 io_in_r_bypass_regNext_14_3_load_store_2;
  reg                 io_in_r_bypass_regNext_14_3_df_is_ws_2;
  reg                 io_in_r_bypass_regNext_14_3_stall_2;
  reg        [15:0]   io_in_r_bypass_regNext_15_0_data_2;
  reg                 io_in_r_bypass_regNext_15_0_load_store_2;
  reg                 io_in_r_bypass_regNext_15_0_df_is_ws_2;
  reg                 io_in_r_bypass_regNext_15_0_stall_2;
  reg        [15:0]   io_in_r_bypass_regNext_15_1_data_2;
  reg                 io_in_r_bypass_regNext_15_1_load_store_2;
  reg                 io_in_r_bypass_regNext_15_1_df_is_ws_2;
  reg                 io_in_r_bypass_regNext_15_1_stall_2;
  reg        [15:0]   io_in_r_bypass_regNext_15_2_data_2;
  reg                 io_in_r_bypass_regNext_15_2_load_store_2;
  reg                 io_in_r_bypass_regNext_15_2_df_is_ws_2;
  reg                 io_in_r_bypass_regNext_15_2_stall_2;
  reg        [15:0]   io_in_r_bypass_regNext_15_3_data_2;
  reg                 io_in_r_bypass_regNext_15_3_load_store_2;
  reg                 io_in_r_bypass_regNext_15_3_df_is_ws_2;
  reg                 io_in_r_bypass_regNext_15_3_stall_2;
  reg        [15:0]   io_in_r_bypass_regNext_16_0_data_2;
  reg                 io_in_r_bypass_regNext_16_0_load_store_2;
  reg                 io_in_r_bypass_regNext_16_0_df_is_ws_2;
  reg                 io_in_r_bypass_regNext_16_0_stall_2;
  reg        [15:0]   io_in_r_bypass_regNext_16_1_data_2;
  reg                 io_in_r_bypass_regNext_16_1_load_store_2;
  reg                 io_in_r_bypass_regNext_16_1_df_is_ws_2;
  reg                 io_in_r_bypass_regNext_16_1_stall_2;
  reg        [15:0]   io_in_r_bypass_regNext_16_2_data_2;
  reg                 io_in_r_bypass_regNext_16_2_load_store_2;
  reg                 io_in_r_bypass_regNext_16_2_df_is_ws_2;
  reg                 io_in_r_bypass_regNext_16_2_stall_2;
  reg        [15:0]   io_in_r_bypass_regNext_16_3_data_2;
  reg                 io_in_r_bypass_regNext_16_3_load_store_2;
  reg                 io_in_r_bypass_regNext_16_3_df_is_ws_2;
  reg                 io_in_r_bypass_regNext_16_3_stall_2;
  reg        [15:0]   io_in_r_bypass_regNext_17_0_data_2;
  reg                 io_in_r_bypass_regNext_17_0_load_store_2;
  reg                 io_in_r_bypass_regNext_17_0_df_is_ws_2;
  reg                 io_in_r_bypass_regNext_17_0_stall_2;
  reg        [15:0]   io_in_r_bypass_regNext_17_1_data_2;
  reg                 io_in_r_bypass_regNext_17_1_load_store_2;
  reg                 io_in_r_bypass_regNext_17_1_df_is_ws_2;
  reg                 io_in_r_bypass_regNext_17_1_stall_2;
  reg        [15:0]   io_in_r_bypass_regNext_17_2_data_2;
  reg                 io_in_r_bypass_regNext_17_2_load_store_2;
  reg                 io_in_r_bypass_regNext_17_2_df_is_ws_2;
  reg                 io_in_r_bypass_regNext_17_2_stall_2;
  reg        [15:0]   io_in_r_bypass_regNext_17_3_data_2;
  reg                 io_in_r_bypass_regNext_17_3_load_store_2;
  reg                 io_in_r_bypass_regNext_17_3_df_is_ws_2;
  reg                 io_in_r_bypass_regNext_17_3_stall_2;
  reg        [15:0]   io_in_r_bypass_regNext_18_0_data_2;
  reg                 io_in_r_bypass_regNext_18_0_load_store_2;
  reg                 io_in_r_bypass_regNext_18_0_df_is_ws_2;
  reg                 io_in_r_bypass_regNext_18_0_stall_2;
  reg        [15:0]   io_in_r_bypass_regNext_18_1_data_2;
  reg                 io_in_r_bypass_regNext_18_1_load_store_2;
  reg                 io_in_r_bypass_regNext_18_1_df_is_ws_2;
  reg                 io_in_r_bypass_regNext_18_1_stall_2;
  reg        [15:0]   io_in_r_bypass_regNext_18_2_data_2;
  reg                 io_in_r_bypass_regNext_18_2_load_store_2;
  reg                 io_in_r_bypass_regNext_18_2_df_is_ws_2;
  reg                 io_in_r_bypass_regNext_18_2_stall_2;
  reg        [15:0]   io_in_r_bypass_regNext_18_3_data_2;
  reg                 io_in_r_bypass_regNext_18_3_load_store_2;
  reg                 io_in_r_bypass_regNext_18_3_df_is_ws_2;
  reg                 io_in_r_bypass_regNext_18_3_stall_2;
  reg        [15:0]   io_in_r_bypass_regNext_19_0_data_2;
  reg                 io_in_r_bypass_regNext_19_0_load_store_2;
  reg                 io_in_r_bypass_regNext_19_0_df_is_ws_2;
  reg                 io_in_r_bypass_regNext_19_0_stall_2;
  reg        [15:0]   io_in_r_bypass_regNext_19_1_data_2;
  reg                 io_in_r_bypass_regNext_19_1_load_store_2;
  reg                 io_in_r_bypass_regNext_19_1_df_is_ws_2;
  reg                 io_in_r_bypass_regNext_19_1_stall_2;
  reg        [15:0]   io_in_r_bypass_regNext_19_2_data_2;
  reg                 io_in_r_bypass_regNext_19_2_load_store_2;
  reg                 io_in_r_bypass_regNext_19_2_df_is_ws_2;
  reg                 io_in_r_bypass_regNext_19_2_stall_2;
  reg        [15:0]   io_in_r_bypass_regNext_19_3_data_2;
  reg                 io_in_r_bypass_regNext_19_3_load_store_2;
  reg                 io_in_r_bypass_regNext_19_3_df_is_ws_2;
  reg                 io_in_r_bypass_regNext_19_3_stall_2;
  reg        [15:0]   io_in_r_bypass_regNext_20_0_data_2;
  reg                 io_in_r_bypass_regNext_20_0_load_store_2;
  reg                 io_in_r_bypass_regNext_20_0_df_is_ws_2;
  reg                 io_in_r_bypass_regNext_20_0_stall_2;
  reg        [15:0]   io_in_r_bypass_regNext_20_1_data_2;
  reg                 io_in_r_bypass_regNext_20_1_load_store_2;
  reg                 io_in_r_bypass_regNext_20_1_df_is_ws_2;
  reg                 io_in_r_bypass_regNext_20_1_stall_2;
  reg        [15:0]   io_in_r_bypass_regNext_20_2_data_2;
  reg                 io_in_r_bypass_regNext_20_2_load_store_2;
  reg                 io_in_r_bypass_regNext_20_2_df_is_ws_2;
  reg                 io_in_r_bypass_regNext_20_2_stall_2;
  reg        [15:0]   io_in_r_bypass_regNext_20_3_data_2;
  reg                 io_in_r_bypass_regNext_20_3_load_store_2;
  reg                 io_in_r_bypass_regNext_20_3_df_is_ws_2;
  reg                 io_in_r_bypass_regNext_20_3_stall_2;
  reg        [15:0]   io_in_r_bypass_regNext_21_0_data_2;
  reg                 io_in_r_bypass_regNext_21_0_load_store_2;
  reg                 io_in_r_bypass_regNext_21_0_df_is_ws_2;
  reg                 io_in_r_bypass_regNext_21_0_stall_2;
  reg        [15:0]   io_in_r_bypass_regNext_21_1_data_2;
  reg                 io_in_r_bypass_regNext_21_1_load_store_2;
  reg                 io_in_r_bypass_regNext_21_1_df_is_ws_2;
  reg                 io_in_r_bypass_regNext_21_1_stall_2;
  reg        [15:0]   io_in_r_bypass_regNext_21_2_data_2;
  reg                 io_in_r_bypass_regNext_21_2_load_store_2;
  reg                 io_in_r_bypass_regNext_21_2_df_is_ws_2;
  reg                 io_in_r_bypass_regNext_21_2_stall_2;
  reg        [15:0]   io_in_r_bypass_regNext_21_3_data_2;
  reg                 io_in_r_bypass_regNext_21_3_load_store_2;
  reg                 io_in_r_bypass_regNext_21_3_df_is_ws_2;
  reg                 io_in_r_bypass_regNext_21_3_stall_2;
  reg        [15:0]   io_in_r_bypass_regNext_22_0_data_2;
  reg                 io_in_r_bypass_regNext_22_0_load_store_2;
  reg                 io_in_r_bypass_regNext_22_0_df_is_ws_2;
  reg                 io_in_r_bypass_regNext_22_0_stall_2;
  reg        [15:0]   io_in_r_bypass_regNext_22_1_data_2;
  reg                 io_in_r_bypass_regNext_22_1_load_store_2;
  reg                 io_in_r_bypass_regNext_22_1_df_is_ws_2;
  reg                 io_in_r_bypass_regNext_22_1_stall_2;
  reg        [15:0]   io_in_r_bypass_regNext_22_2_data_2;
  reg                 io_in_r_bypass_regNext_22_2_load_store_2;
  reg                 io_in_r_bypass_regNext_22_2_df_is_ws_2;
  reg                 io_in_r_bypass_regNext_22_2_stall_2;
  reg        [15:0]   io_in_r_bypass_regNext_22_3_data_2;
  reg                 io_in_r_bypass_regNext_22_3_load_store_2;
  reg                 io_in_r_bypass_regNext_22_3_df_is_ws_2;
  reg                 io_in_r_bypass_regNext_22_3_stall_2;
  reg        [15:0]   io_in_r_bypass_regNext_23_0_data_2;
  reg                 io_in_r_bypass_regNext_23_0_load_store_2;
  reg                 io_in_r_bypass_regNext_23_0_df_is_ws_2;
  reg                 io_in_r_bypass_regNext_23_0_stall_2;
  reg        [15:0]   io_in_r_bypass_regNext_23_1_data_2;
  reg                 io_in_r_bypass_regNext_23_1_load_store_2;
  reg                 io_in_r_bypass_regNext_23_1_df_is_ws_2;
  reg                 io_in_r_bypass_regNext_23_1_stall_2;
  reg        [15:0]   io_in_r_bypass_regNext_23_2_data_2;
  reg                 io_in_r_bypass_regNext_23_2_load_store_2;
  reg                 io_in_r_bypass_regNext_23_2_df_is_ws_2;
  reg                 io_in_r_bypass_regNext_23_2_stall_2;
  reg        [15:0]   io_in_r_bypass_regNext_23_3_data_2;
  reg                 io_in_r_bypass_regNext_23_3_load_store_2;
  reg                 io_in_r_bypass_regNext_23_3_df_is_ws_2;
  reg                 io_in_r_bypass_regNext_23_3_stall_2;
  reg        [15:0]   io_in_r_bypass_regNext_24_0_data_2;
  reg                 io_in_r_bypass_regNext_24_0_load_store_2;
  reg                 io_in_r_bypass_regNext_24_0_df_is_ws_2;
  reg                 io_in_r_bypass_regNext_24_0_stall_2;
  reg        [15:0]   io_in_r_bypass_regNext_24_1_data_2;
  reg                 io_in_r_bypass_regNext_24_1_load_store_2;
  reg                 io_in_r_bypass_regNext_24_1_df_is_ws_2;
  reg                 io_in_r_bypass_regNext_24_1_stall_2;
  reg        [15:0]   io_in_r_bypass_regNext_24_2_data_2;
  reg                 io_in_r_bypass_regNext_24_2_load_store_2;
  reg                 io_in_r_bypass_regNext_24_2_df_is_ws_2;
  reg                 io_in_r_bypass_regNext_24_2_stall_2;
  reg        [15:0]   io_in_r_bypass_regNext_24_3_data_2;
  reg                 io_in_r_bypass_regNext_24_3_load_store_2;
  reg                 io_in_r_bypass_regNext_24_3_df_is_ws_2;
  reg                 io_in_r_bypass_regNext_24_3_stall_2;
  reg        [15:0]   io_in_r_bypass_regNext_25_0_data_2;
  reg                 io_in_r_bypass_regNext_25_0_load_store_2;
  reg                 io_in_r_bypass_regNext_25_0_df_is_ws_2;
  reg                 io_in_r_bypass_regNext_25_0_stall_2;
  reg        [15:0]   io_in_r_bypass_regNext_25_1_data_2;
  reg                 io_in_r_bypass_regNext_25_1_load_store_2;
  reg                 io_in_r_bypass_regNext_25_1_df_is_ws_2;
  reg                 io_in_r_bypass_regNext_25_1_stall_2;
  reg        [15:0]   io_in_r_bypass_regNext_25_2_data_2;
  reg                 io_in_r_bypass_regNext_25_2_load_store_2;
  reg                 io_in_r_bypass_regNext_25_2_df_is_ws_2;
  reg                 io_in_r_bypass_regNext_25_2_stall_2;
  reg        [15:0]   io_in_r_bypass_regNext_25_3_data_2;
  reg                 io_in_r_bypass_regNext_25_3_load_store_2;
  reg                 io_in_r_bypass_regNext_25_3_df_is_ws_2;
  reg                 io_in_r_bypass_regNext_25_3_stall_2;
  reg        [15:0]   io_in_r_bypass_regNext_26_0_data_2;
  reg                 io_in_r_bypass_regNext_26_0_load_store_2;
  reg                 io_in_r_bypass_regNext_26_0_df_is_ws_2;
  reg                 io_in_r_bypass_regNext_26_0_stall_2;
  reg        [15:0]   io_in_r_bypass_regNext_26_1_data_2;
  reg                 io_in_r_bypass_regNext_26_1_load_store_2;
  reg                 io_in_r_bypass_regNext_26_1_df_is_ws_2;
  reg                 io_in_r_bypass_regNext_26_1_stall_2;
  reg        [15:0]   io_in_r_bypass_regNext_26_2_data_2;
  reg                 io_in_r_bypass_regNext_26_2_load_store_2;
  reg                 io_in_r_bypass_regNext_26_2_df_is_ws_2;
  reg                 io_in_r_bypass_regNext_26_2_stall_2;
  reg        [15:0]   io_in_r_bypass_regNext_26_3_data_2;
  reg                 io_in_r_bypass_regNext_26_3_load_store_2;
  reg                 io_in_r_bypass_regNext_26_3_df_is_ws_2;
  reg                 io_in_r_bypass_regNext_26_3_stall_2;
  reg        [15:0]   io_in_r_bypass_regNext_27_0_data_2;
  reg                 io_in_r_bypass_regNext_27_0_load_store_2;
  reg                 io_in_r_bypass_regNext_27_0_df_is_ws_2;
  reg                 io_in_r_bypass_regNext_27_0_stall_2;
  reg        [15:0]   io_in_r_bypass_regNext_27_1_data_2;
  reg                 io_in_r_bypass_regNext_27_1_load_store_2;
  reg                 io_in_r_bypass_regNext_27_1_df_is_ws_2;
  reg                 io_in_r_bypass_regNext_27_1_stall_2;
  reg        [15:0]   io_in_r_bypass_regNext_27_2_data_2;
  reg                 io_in_r_bypass_regNext_27_2_load_store_2;
  reg                 io_in_r_bypass_regNext_27_2_df_is_ws_2;
  reg                 io_in_r_bypass_regNext_27_2_stall_2;
  reg        [15:0]   io_in_r_bypass_regNext_27_3_data_2;
  reg                 io_in_r_bypass_regNext_27_3_load_store_2;
  reg                 io_in_r_bypass_regNext_27_3_df_is_ws_2;
  reg                 io_in_r_bypass_regNext_27_3_stall_2;
  reg        [15:0]   io_in_r_bypass_regNext_28_0_data_2;
  reg                 io_in_r_bypass_regNext_28_0_load_store_2;
  reg                 io_in_r_bypass_regNext_28_0_df_is_ws_2;
  reg                 io_in_r_bypass_regNext_28_0_stall_2;
  reg        [15:0]   io_in_r_bypass_regNext_28_1_data_2;
  reg                 io_in_r_bypass_regNext_28_1_load_store_2;
  reg                 io_in_r_bypass_regNext_28_1_df_is_ws_2;
  reg                 io_in_r_bypass_regNext_28_1_stall_2;
  reg        [15:0]   io_in_r_bypass_regNext_28_2_data_2;
  reg                 io_in_r_bypass_regNext_28_2_load_store_2;
  reg                 io_in_r_bypass_regNext_28_2_df_is_ws_2;
  reg                 io_in_r_bypass_regNext_28_2_stall_2;
  reg        [15:0]   io_in_r_bypass_regNext_28_3_data_2;
  reg                 io_in_r_bypass_regNext_28_3_load_store_2;
  reg                 io_in_r_bypass_regNext_28_3_df_is_ws_2;
  reg                 io_in_r_bypass_regNext_28_3_stall_2;
  reg        [15:0]   io_in_r_bypass_regNext_29_0_data_2;
  reg                 io_in_r_bypass_regNext_29_0_load_store_2;
  reg                 io_in_r_bypass_regNext_29_0_df_is_ws_2;
  reg                 io_in_r_bypass_regNext_29_0_stall_2;
  reg        [15:0]   io_in_r_bypass_regNext_29_1_data_2;
  reg                 io_in_r_bypass_regNext_29_1_load_store_2;
  reg                 io_in_r_bypass_regNext_29_1_df_is_ws_2;
  reg                 io_in_r_bypass_regNext_29_1_stall_2;
  reg        [15:0]   io_in_r_bypass_regNext_29_2_data_2;
  reg                 io_in_r_bypass_regNext_29_2_load_store_2;
  reg                 io_in_r_bypass_regNext_29_2_df_is_ws_2;
  reg                 io_in_r_bypass_regNext_29_2_stall_2;
  reg        [15:0]   io_in_r_bypass_regNext_29_3_data_2;
  reg                 io_in_r_bypass_regNext_29_3_load_store_2;
  reg                 io_in_r_bypass_regNext_29_3_df_is_ws_2;
  reg                 io_in_r_bypass_regNext_29_3_stall_2;
  reg        [15:0]   io_in_r_bypass_regNext_30_0_data_2;
  reg                 io_in_r_bypass_regNext_30_0_load_store_2;
  reg                 io_in_r_bypass_regNext_30_0_df_is_ws_2;
  reg                 io_in_r_bypass_regNext_30_0_stall_2;
  reg        [15:0]   io_in_r_bypass_regNext_30_1_data_2;
  reg                 io_in_r_bypass_regNext_30_1_load_store_2;
  reg                 io_in_r_bypass_regNext_30_1_df_is_ws_2;
  reg                 io_in_r_bypass_regNext_30_1_stall_2;
  reg        [15:0]   io_in_r_bypass_regNext_30_2_data_2;
  reg                 io_in_r_bypass_regNext_30_2_load_store_2;
  reg                 io_in_r_bypass_regNext_30_2_df_is_ws_2;
  reg                 io_in_r_bypass_regNext_30_2_stall_2;
  reg        [15:0]   io_in_r_bypass_regNext_30_3_data_2;
  reg                 io_in_r_bypass_regNext_30_3_load_store_2;
  reg                 io_in_r_bypass_regNext_30_3_df_is_ws_2;
  reg                 io_in_r_bypass_regNext_30_3_stall_2;
  reg        [15:0]   io_in_r_bypass_regNext_31_0_data_2;
  reg                 io_in_r_bypass_regNext_31_0_load_store_2;
  reg                 io_in_r_bypass_regNext_31_0_df_is_ws_2;
  reg                 io_in_r_bypass_regNext_31_0_stall_2;
  reg        [15:0]   io_in_r_bypass_regNext_31_1_data_2;
  reg                 io_in_r_bypass_regNext_31_1_load_store_2;
  reg                 io_in_r_bypass_regNext_31_1_df_is_ws_2;
  reg                 io_in_r_bypass_regNext_31_1_stall_2;
  reg        [15:0]   io_in_r_bypass_regNext_31_2_data_2;
  reg                 io_in_r_bypass_regNext_31_2_load_store_2;
  reg                 io_in_r_bypass_regNext_31_2_df_is_ws_2;
  reg                 io_in_r_bypass_regNext_31_2_stall_2;
  reg        [15:0]   io_in_r_bypass_regNext_31_3_data_2;
  reg                 io_in_r_bypass_regNext_31_3_load_store_2;
  reg                 io_in_r_bypass_regNext_31_3_df_is_ws_2;
  reg                 io_in_r_bypass_regNext_31_3_stall_2;
  reg        [15:0]   io_in_r_bypass_regNext_0_0_data_3;
  reg                 io_in_r_bypass_regNext_0_0_load_store_3;
  reg                 io_in_r_bypass_regNext_0_0_df_is_ws_3;
  reg                 io_in_r_bypass_regNext_0_0_stall_3;
  reg        [15:0]   io_in_r_bypass_regNext_0_1_data_3;
  reg                 io_in_r_bypass_regNext_0_1_load_store_3;
  reg                 io_in_r_bypass_regNext_0_1_df_is_ws_3;
  reg                 io_in_r_bypass_regNext_0_1_stall_3;
  reg        [15:0]   io_in_r_bypass_regNext_0_2_data_3;
  reg                 io_in_r_bypass_regNext_0_2_load_store_3;
  reg                 io_in_r_bypass_regNext_0_2_df_is_ws_3;
  reg                 io_in_r_bypass_regNext_0_2_stall_3;
  reg        [15:0]   io_in_r_bypass_regNext_0_3_data_3;
  reg                 io_in_r_bypass_regNext_0_3_load_store_3;
  reg                 io_in_r_bypass_regNext_0_3_df_is_ws_3;
  reg                 io_in_r_bypass_regNext_0_3_stall_3;
  reg        [15:0]   io_in_r_bypass_regNext_1_0_data_3;
  reg                 io_in_r_bypass_regNext_1_0_load_store_3;
  reg                 io_in_r_bypass_regNext_1_0_df_is_ws_3;
  reg                 io_in_r_bypass_regNext_1_0_stall_3;
  reg        [15:0]   io_in_r_bypass_regNext_1_1_data_3;
  reg                 io_in_r_bypass_regNext_1_1_load_store_3;
  reg                 io_in_r_bypass_regNext_1_1_df_is_ws_3;
  reg                 io_in_r_bypass_regNext_1_1_stall_3;
  reg        [15:0]   io_in_r_bypass_regNext_1_2_data_3;
  reg                 io_in_r_bypass_regNext_1_2_load_store_3;
  reg                 io_in_r_bypass_regNext_1_2_df_is_ws_3;
  reg                 io_in_r_bypass_regNext_1_2_stall_3;
  reg        [15:0]   io_in_r_bypass_regNext_1_3_data_3;
  reg                 io_in_r_bypass_regNext_1_3_load_store_3;
  reg                 io_in_r_bypass_regNext_1_3_df_is_ws_3;
  reg                 io_in_r_bypass_regNext_1_3_stall_3;
  reg        [15:0]   io_in_r_bypass_regNext_2_0_data_3;
  reg                 io_in_r_bypass_regNext_2_0_load_store_3;
  reg                 io_in_r_bypass_regNext_2_0_df_is_ws_3;
  reg                 io_in_r_bypass_regNext_2_0_stall_3;
  reg        [15:0]   io_in_r_bypass_regNext_2_1_data_3;
  reg                 io_in_r_bypass_regNext_2_1_load_store_3;
  reg                 io_in_r_bypass_regNext_2_1_df_is_ws_3;
  reg                 io_in_r_bypass_regNext_2_1_stall_3;
  reg        [15:0]   io_in_r_bypass_regNext_2_2_data_3;
  reg                 io_in_r_bypass_regNext_2_2_load_store_3;
  reg                 io_in_r_bypass_regNext_2_2_df_is_ws_3;
  reg                 io_in_r_bypass_regNext_2_2_stall_3;
  reg        [15:0]   io_in_r_bypass_regNext_2_3_data_3;
  reg                 io_in_r_bypass_regNext_2_3_load_store_3;
  reg                 io_in_r_bypass_regNext_2_3_df_is_ws_3;
  reg                 io_in_r_bypass_regNext_2_3_stall_3;
  reg        [15:0]   io_in_r_bypass_regNext_3_0_data_3;
  reg                 io_in_r_bypass_regNext_3_0_load_store_3;
  reg                 io_in_r_bypass_regNext_3_0_df_is_ws_3;
  reg                 io_in_r_bypass_regNext_3_0_stall_3;
  reg        [15:0]   io_in_r_bypass_regNext_3_1_data_3;
  reg                 io_in_r_bypass_regNext_3_1_load_store_3;
  reg                 io_in_r_bypass_regNext_3_1_df_is_ws_3;
  reg                 io_in_r_bypass_regNext_3_1_stall_3;
  reg        [15:0]   io_in_r_bypass_regNext_3_2_data_3;
  reg                 io_in_r_bypass_regNext_3_2_load_store_3;
  reg                 io_in_r_bypass_regNext_3_2_df_is_ws_3;
  reg                 io_in_r_bypass_regNext_3_2_stall_3;
  reg        [15:0]   io_in_r_bypass_regNext_3_3_data_3;
  reg                 io_in_r_bypass_regNext_3_3_load_store_3;
  reg                 io_in_r_bypass_regNext_3_3_df_is_ws_3;
  reg                 io_in_r_bypass_regNext_3_3_stall_3;
  reg        [15:0]   io_in_r_bypass_regNext_4_0_data_3;
  reg                 io_in_r_bypass_regNext_4_0_load_store_3;
  reg                 io_in_r_bypass_regNext_4_0_df_is_ws_3;
  reg                 io_in_r_bypass_regNext_4_0_stall_3;
  reg        [15:0]   io_in_r_bypass_regNext_4_1_data_3;
  reg                 io_in_r_bypass_regNext_4_1_load_store_3;
  reg                 io_in_r_bypass_regNext_4_1_df_is_ws_3;
  reg                 io_in_r_bypass_regNext_4_1_stall_3;
  reg        [15:0]   io_in_r_bypass_regNext_4_2_data_3;
  reg                 io_in_r_bypass_regNext_4_2_load_store_3;
  reg                 io_in_r_bypass_regNext_4_2_df_is_ws_3;
  reg                 io_in_r_bypass_regNext_4_2_stall_3;
  reg        [15:0]   io_in_r_bypass_regNext_4_3_data_3;
  reg                 io_in_r_bypass_regNext_4_3_load_store_3;
  reg                 io_in_r_bypass_regNext_4_3_df_is_ws_3;
  reg                 io_in_r_bypass_regNext_4_3_stall_3;
  reg        [15:0]   io_in_r_bypass_regNext_5_0_data_3;
  reg                 io_in_r_bypass_regNext_5_0_load_store_3;
  reg                 io_in_r_bypass_regNext_5_0_df_is_ws_3;
  reg                 io_in_r_bypass_regNext_5_0_stall_3;
  reg        [15:0]   io_in_r_bypass_regNext_5_1_data_3;
  reg                 io_in_r_bypass_regNext_5_1_load_store_3;
  reg                 io_in_r_bypass_regNext_5_1_df_is_ws_3;
  reg                 io_in_r_bypass_regNext_5_1_stall_3;
  reg        [15:0]   io_in_r_bypass_regNext_5_2_data_3;
  reg                 io_in_r_bypass_regNext_5_2_load_store_3;
  reg                 io_in_r_bypass_regNext_5_2_df_is_ws_3;
  reg                 io_in_r_bypass_regNext_5_2_stall_3;
  reg        [15:0]   io_in_r_bypass_regNext_5_3_data_3;
  reg                 io_in_r_bypass_regNext_5_3_load_store_3;
  reg                 io_in_r_bypass_regNext_5_3_df_is_ws_3;
  reg                 io_in_r_bypass_regNext_5_3_stall_3;
  reg        [15:0]   io_in_r_bypass_regNext_6_0_data_3;
  reg                 io_in_r_bypass_regNext_6_0_load_store_3;
  reg                 io_in_r_bypass_regNext_6_0_df_is_ws_3;
  reg                 io_in_r_bypass_regNext_6_0_stall_3;
  reg        [15:0]   io_in_r_bypass_regNext_6_1_data_3;
  reg                 io_in_r_bypass_regNext_6_1_load_store_3;
  reg                 io_in_r_bypass_regNext_6_1_df_is_ws_3;
  reg                 io_in_r_bypass_regNext_6_1_stall_3;
  reg        [15:0]   io_in_r_bypass_regNext_6_2_data_3;
  reg                 io_in_r_bypass_regNext_6_2_load_store_3;
  reg                 io_in_r_bypass_regNext_6_2_df_is_ws_3;
  reg                 io_in_r_bypass_regNext_6_2_stall_3;
  reg        [15:0]   io_in_r_bypass_regNext_6_3_data_3;
  reg                 io_in_r_bypass_regNext_6_3_load_store_3;
  reg                 io_in_r_bypass_regNext_6_3_df_is_ws_3;
  reg                 io_in_r_bypass_regNext_6_3_stall_3;
  reg        [15:0]   io_in_r_bypass_regNext_7_0_data_3;
  reg                 io_in_r_bypass_regNext_7_0_load_store_3;
  reg                 io_in_r_bypass_regNext_7_0_df_is_ws_3;
  reg                 io_in_r_bypass_regNext_7_0_stall_3;
  reg        [15:0]   io_in_r_bypass_regNext_7_1_data_3;
  reg                 io_in_r_bypass_regNext_7_1_load_store_3;
  reg                 io_in_r_bypass_regNext_7_1_df_is_ws_3;
  reg                 io_in_r_bypass_regNext_7_1_stall_3;
  reg        [15:0]   io_in_r_bypass_regNext_7_2_data_3;
  reg                 io_in_r_bypass_regNext_7_2_load_store_3;
  reg                 io_in_r_bypass_regNext_7_2_df_is_ws_3;
  reg                 io_in_r_bypass_regNext_7_2_stall_3;
  reg        [15:0]   io_in_r_bypass_regNext_7_3_data_3;
  reg                 io_in_r_bypass_regNext_7_3_load_store_3;
  reg                 io_in_r_bypass_regNext_7_3_df_is_ws_3;
  reg                 io_in_r_bypass_regNext_7_3_stall_3;
  reg        [15:0]   io_in_r_bypass_regNext_8_0_data_3;
  reg                 io_in_r_bypass_regNext_8_0_load_store_3;
  reg                 io_in_r_bypass_regNext_8_0_df_is_ws_3;
  reg                 io_in_r_bypass_regNext_8_0_stall_3;
  reg        [15:0]   io_in_r_bypass_regNext_8_1_data_3;
  reg                 io_in_r_bypass_regNext_8_1_load_store_3;
  reg                 io_in_r_bypass_regNext_8_1_df_is_ws_3;
  reg                 io_in_r_bypass_regNext_8_1_stall_3;
  reg        [15:0]   io_in_r_bypass_regNext_8_2_data_3;
  reg                 io_in_r_bypass_regNext_8_2_load_store_3;
  reg                 io_in_r_bypass_regNext_8_2_df_is_ws_3;
  reg                 io_in_r_bypass_regNext_8_2_stall_3;
  reg        [15:0]   io_in_r_bypass_regNext_8_3_data_3;
  reg                 io_in_r_bypass_regNext_8_3_load_store_3;
  reg                 io_in_r_bypass_regNext_8_3_df_is_ws_3;
  reg                 io_in_r_bypass_regNext_8_3_stall_3;
  reg        [15:0]   io_in_r_bypass_regNext_9_0_data_3;
  reg                 io_in_r_bypass_regNext_9_0_load_store_3;
  reg                 io_in_r_bypass_regNext_9_0_df_is_ws_3;
  reg                 io_in_r_bypass_regNext_9_0_stall_3;
  reg        [15:0]   io_in_r_bypass_regNext_9_1_data_3;
  reg                 io_in_r_bypass_regNext_9_1_load_store_3;
  reg                 io_in_r_bypass_regNext_9_1_df_is_ws_3;
  reg                 io_in_r_bypass_regNext_9_1_stall_3;
  reg        [15:0]   io_in_r_bypass_regNext_9_2_data_3;
  reg                 io_in_r_bypass_regNext_9_2_load_store_3;
  reg                 io_in_r_bypass_regNext_9_2_df_is_ws_3;
  reg                 io_in_r_bypass_regNext_9_2_stall_3;
  reg        [15:0]   io_in_r_bypass_regNext_9_3_data_3;
  reg                 io_in_r_bypass_regNext_9_3_load_store_3;
  reg                 io_in_r_bypass_regNext_9_3_df_is_ws_3;
  reg                 io_in_r_bypass_regNext_9_3_stall_3;
  reg        [15:0]   io_in_r_bypass_regNext_10_0_data_3;
  reg                 io_in_r_bypass_regNext_10_0_load_store_3;
  reg                 io_in_r_bypass_regNext_10_0_df_is_ws_3;
  reg                 io_in_r_bypass_regNext_10_0_stall_3;
  reg        [15:0]   io_in_r_bypass_regNext_10_1_data_3;
  reg                 io_in_r_bypass_regNext_10_1_load_store_3;
  reg                 io_in_r_bypass_regNext_10_1_df_is_ws_3;
  reg                 io_in_r_bypass_regNext_10_1_stall_3;
  reg        [15:0]   io_in_r_bypass_regNext_10_2_data_3;
  reg                 io_in_r_bypass_regNext_10_2_load_store_3;
  reg                 io_in_r_bypass_regNext_10_2_df_is_ws_3;
  reg                 io_in_r_bypass_regNext_10_2_stall_3;
  reg        [15:0]   io_in_r_bypass_regNext_10_3_data_3;
  reg                 io_in_r_bypass_regNext_10_3_load_store_3;
  reg                 io_in_r_bypass_regNext_10_3_df_is_ws_3;
  reg                 io_in_r_bypass_regNext_10_3_stall_3;
  reg        [15:0]   io_in_r_bypass_regNext_11_0_data_3;
  reg                 io_in_r_bypass_regNext_11_0_load_store_3;
  reg                 io_in_r_bypass_regNext_11_0_df_is_ws_3;
  reg                 io_in_r_bypass_regNext_11_0_stall_3;
  reg        [15:0]   io_in_r_bypass_regNext_11_1_data_3;
  reg                 io_in_r_bypass_regNext_11_1_load_store_3;
  reg                 io_in_r_bypass_regNext_11_1_df_is_ws_3;
  reg                 io_in_r_bypass_regNext_11_1_stall_3;
  reg        [15:0]   io_in_r_bypass_regNext_11_2_data_3;
  reg                 io_in_r_bypass_regNext_11_2_load_store_3;
  reg                 io_in_r_bypass_regNext_11_2_df_is_ws_3;
  reg                 io_in_r_bypass_regNext_11_2_stall_3;
  reg        [15:0]   io_in_r_bypass_regNext_11_3_data_3;
  reg                 io_in_r_bypass_regNext_11_3_load_store_3;
  reg                 io_in_r_bypass_regNext_11_3_df_is_ws_3;
  reg                 io_in_r_bypass_regNext_11_3_stall_3;
  reg        [15:0]   io_in_r_bypass_regNext_12_0_data_3;
  reg                 io_in_r_bypass_regNext_12_0_load_store_3;
  reg                 io_in_r_bypass_regNext_12_0_df_is_ws_3;
  reg                 io_in_r_bypass_regNext_12_0_stall_3;
  reg        [15:0]   io_in_r_bypass_regNext_12_1_data_3;
  reg                 io_in_r_bypass_regNext_12_1_load_store_3;
  reg                 io_in_r_bypass_regNext_12_1_df_is_ws_3;
  reg                 io_in_r_bypass_regNext_12_1_stall_3;
  reg        [15:0]   io_in_r_bypass_regNext_12_2_data_3;
  reg                 io_in_r_bypass_regNext_12_2_load_store_3;
  reg                 io_in_r_bypass_regNext_12_2_df_is_ws_3;
  reg                 io_in_r_bypass_regNext_12_2_stall_3;
  reg        [15:0]   io_in_r_bypass_regNext_12_3_data_3;
  reg                 io_in_r_bypass_regNext_12_3_load_store_3;
  reg                 io_in_r_bypass_regNext_12_3_df_is_ws_3;
  reg                 io_in_r_bypass_regNext_12_3_stall_3;
  reg        [15:0]   io_in_r_bypass_regNext_13_0_data_3;
  reg                 io_in_r_bypass_regNext_13_0_load_store_3;
  reg                 io_in_r_bypass_regNext_13_0_df_is_ws_3;
  reg                 io_in_r_bypass_regNext_13_0_stall_3;
  reg        [15:0]   io_in_r_bypass_regNext_13_1_data_3;
  reg                 io_in_r_bypass_regNext_13_1_load_store_3;
  reg                 io_in_r_bypass_regNext_13_1_df_is_ws_3;
  reg                 io_in_r_bypass_regNext_13_1_stall_3;
  reg        [15:0]   io_in_r_bypass_regNext_13_2_data_3;
  reg                 io_in_r_bypass_regNext_13_2_load_store_3;
  reg                 io_in_r_bypass_regNext_13_2_df_is_ws_3;
  reg                 io_in_r_bypass_regNext_13_2_stall_3;
  reg        [15:0]   io_in_r_bypass_regNext_13_3_data_3;
  reg                 io_in_r_bypass_regNext_13_3_load_store_3;
  reg                 io_in_r_bypass_regNext_13_3_df_is_ws_3;
  reg                 io_in_r_bypass_regNext_13_3_stall_3;
  reg        [15:0]   io_in_r_bypass_regNext_14_0_data_3;
  reg                 io_in_r_bypass_regNext_14_0_load_store_3;
  reg                 io_in_r_bypass_regNext_14_0_df_is_ws_3;
  reg                 io_in_r_bypass_regNext_14_0_stall_3;
  reg        [15:0]   io_in_r_bypass_regNext_14_1_data_3;
  reg                 io_in_r_bypass_regNext_14_1_load_store_3;
  reg                 io_in_r_bypass_regNext_14_1_df_is_ws_3;
  reg                 io_in_r_bypass_regNext_14_1_stall_3;
  reg        [15:0]   io_in_r_bypass_regNext_14_2_data_3;
  reg                 io_in_r_bypass_regNext_14_2_load_store_3;
  reg                 io_in_r_bypass_regNext_14_2_df_is_ws_3;
  reg                 io_in_r_bypass_regNext_14_2_stall_3;
  reg        [15:0]   io_in_r_bypass_regNext_14_3_data_3;
  reg                 io_in_r_bypass_regNext_14_3_load_store_3;
  reg                 io_in_r_bypass_regNext_14_3_df_is_ws_3;
  reg                 io_in_r_bypass_regNext_14_3_stall_3;
  reg        [15:0]   io_in_r_bypass_regNext_15_0_data_3;
  reg                 io_in_r_bypass_regNext_15_0_load_store_3;
  reg                 io_in_r_bypass_regNext_15_0_df_is_ws_3;
  reg                 io_in_r_bypass_regNext_15_0_stall_3;
  reg        [15:0]   io_in_r_bypass_regNext_15_1_data_3;
  reg                 io_in_r_bypass_regNext_15_1_load_store_3;
  reg                 io_in_r_bypass_regNext_15_1_df_is_ws_3;
  reg                 io_in_r_bypass_regNext_15_1_stall_3;
  reg        [15:0]   io_in_r_bypass_regNext_15_2_data_3;
  reg                 io_in_r_bypass_regNext_15_2_load_store_3;
  reg                 io_in_r_bypass_regNext_15_2_df_is_ws_3;
  reg                 io_in_r_bypass_regNext_15_2_stall_3;
  reg        [15:0]   io_in_r_bypass_regNext_15_3_data_3;
  reg                 io_in_r_bypass_regNext_15_3_load_store_3;
  reg                 io_in_r_bypass_regNext_15_3_df_is_ws_3;
  reg                 io_in_r_bypass_regNext_15_3_stall_3;
  reg        [15:0]   io_in_r_bypass_regNext_16_0_data_3;
  reg                 io_in_r_bypass_regNext_16_0_load_store_3;
  reg                 io_in_r_bypass_regNext_16_0_df_is_ws_3;
  reg                 io_in_r_bypass_regNext_16_0_stall_3;
  reg        [15:0]   io_in_r_bypass_regNext_16_1_data_3;
  reg                 io_in_r_bypass_regNext_16_1_load_store_3;
  reg                 io_in_r_bypass_regNext_16_1_df_is_ws_3;
  reg                 io_in_r_bypass_regNext_16_1_stall_3;
  reg        [15:0]   io_in_r_bypass_regNext_16_2_data_3;
  reg                 io_in_r_bypass_regNext_16_2_load_store_3;
  reg                 io_in_r_bypass_regNext_16_2_df_is_ws_3;
  reg                 io_in_r_bypass_regNext_16_2_stall_3;
  reg        [15:0]   io_in_r_bypass_regNext_16_3_data_3;
  reg                 io_in_r_bypass_regNext_16_3_load_store_3;
  reg                 io_in_r_bypass_regNext_16_3_df_is_ws_3;
  reg                 io_in_r_bypass_regNext_16_3_stall_3;
  reg        [15:0]   io_in_r_bypass_regNext_17_0_data_3;
  reg                 io_in_r_bypass_regNext_17_0_load_store_3;
  reg                 io_in_r_bypass_regNext_17_0_df_is_ws_3;
  reg                 io_in_r_bypass_regNext_17_0_stall_3;
  reg        [15:0]   io_in_r_bypass_regNext_17_1_data_3;
  reg                 io_in_r_bypass_regNext_17_1_load_store_3;
  reg                 io_in_r_bypass_regNext_17_1_df_is_ws_3;
  reg                 io_in_r_bypass_regNext_17_1_stall_3;
  reg        [15:0]   io_in_r_bypass_regNext_17_2_data_3;
  reg                 io_in_r_bypass_regNext_17_2_load_store_3;
  reg                 io_in_r_bypass_regNext_17_2_df_is_ws_3;
  reg                 io_in_r_bypass_regNext_17_2_stall_3;
  reg        [15:0]   io_in_r_bypass_regNext_17_3_data_3;
  reg                 io_in_r_bypass_regNext_17_3_load_store_3;
  reg                 io_in_r_bypass_regNext_17_3_df_is_ws_3;
  reg                 io_in_r_bypass_regNext_17_3_stall_3;
  reg        [15:0]   io_in_r_bypass_regNext_18_0_data_3;
  reg                 io_in_r_bypass_regNext_18_0_load_store_3;
  reg                 io_in_r_bypass_regNext_18_0_df_is_ws_3;
  reg                 io_in_r_bypass_regNext_18_0_stall_3;
  reg        [15:0]   io_in_r_bypass_regNext_18_1_data_3;
  reg                 io_in_r_bypass_regNext_18_1_load_store_3;
  reg                 io_in_r_bypass_regNext_18_1_df_is_ws_3;
  reg                 io_in_r_bypass_regNext_18_1_stall_3;
  reg        [15:0]   io_in_r_bypass_regNext_18_2_data_3;
  reg                 io_in_r_bypass_regNext_18_2_load_store_3;
  reg                 io_in_r_bypass_regNext_18_2_df_is_ws_3;
  reg                 io_in_r_bypass_regNext_18_2_stall_3;
  reg        [15:0]   io_in_r_bypass_regNext_18_3_data_3;
  reg                 io_in_r_bypass_regNext_18_3_load_store_3;
  reg                 io_in_r_bypass_regNext_18_3_df_is_ws_3;
  reg                 io_in_r_bypass_regNext_18_3_stall_3;
  reg        [15:0]   io_in_r_bypass_regNext_19_0_data_3;
  reg                 io_in_r_bypass_regNext_19_0_load_store_3;
  reg                 io_in_r_bypass_regNext_19_0_df_is_ws_3;
  reg                 io_in_r_bypass_regNext_19_0_stall_3;
  reg        [15:0]   io_in_r_bypass_regNext_19_1_data_3;
  reg                 io_in_r_bypass_regNext_19_1_load_store_3;
  reg                 io_in_r_bypass_regNext_19_1_df_is_ws_3;
  reg                 io_in_r_bypass_regNext_19_1_stall_3;
  reg        [15:0]   io_in_r_bypass_regNext_19_2_data_3;
  reg                 io_in_r_bypass_regNext_19_2_load_store_3;
  reg                 io_in_r_bypass_regNext_19_2_df_is_ws_3;
  reg                 io_in_r_bypass_regNext_19_2_stall_3;
  reg        [15:0]   io_in_r_bypass_regNext_19_3_data_3;
  reg                 io_in_r_bypass_regNext_19_3_load_store_3;
  reg                 io_in_r_bypass_regNext_19_3_df_is_ws_3;
  reg                 io_in_r_bypass_regNext_19_3_stall_3;
  reg        [15:0]   io_in_r_bypass_regNext_20_0_data_3;
  reg                 io_in_r_bypass_regNext_20_0_load_store_3;
  reg                 io_in_r_bypass_regNext_20_0_df_is_ws_3;
  reg                 io_in_r_bypass_regNext_20_0_stall_3;
  reg        [15:0]   io_in_r_bypass_regNext_20_1_data_3;
  reg                 io_in_r_bypass_regNext_20_1_load_store_3;
  reg                 io_in_r_bypass_regNext_20_1_df_is_ws_3;
  reg                 io_in_r_bypass_regNext_20_1_stall_3;
  reg        [15:0]   io_in_r_bypass_regNext_20_2_data_3;
  reg                 io_in_r_bypass_regNext_20_2_load_store_3;
  reg                 io_in_r_bypass_regNext_20_2_df_is_ws_3;
  reg                 io_in_r_bypass_regNext_20_2_stall_3;
  reg        [15:0]   io_in_r_bypass_regNext_20_3_data_3;
  reg                 io_in_r_bypass_regNext_20_3_load_store_3;
  reg                 io_in_r_bypass_regNext_20_3_df_is_ws_3;
  reg                 io_in_r_bypass_regNext_20_3_stall_3;
  reg        [15:0]   io_in_r_bypass_regNext_21_0_data_3;
  reg                 io_in_r_bypass_regNext_21_0_load_store_3;
  reg                 io_in_r_bypass_regNext_21_0_df_is_ws_3;
  reg                 io_in_r_bypass_regNext_21_0_stall_3;
  reg        [15:0]   io_in_r_bypass_regNext_21_1_data_3;
  reg                 io_in_r_bypass_regNext_21_1_load_store_3;
  reg                 io_in_r_bypass_regNext_21_1_df_is_ws_3;
  reg                 io_in_r_bypass_regNext_21_1_stall_3;
  reg        [15:0]   io_in_r_bypass_regNext_21_2_data_3;
  reg                 io_in_r_bypass_regNext_21_2_load_store_3;
  reg                 io_in_r_bypass_regNext_21_2_df_is_ws_3;
  reg                 io_in_r_bypass_regNext_21_2_stall_3;
  reg        [15:0]   io_in_r_bypass_regNext_21_3_data_3;
  reg                 io_in_r_bypass_regNext_21_3_load_store_3;
  reg                 io_in_r_bypass_regNext_21_3_df_is_ws_3;
  reg                 io_in_r_bypass_regNext_21_3_stall_3;
  reg        [15:0]   io_in_r_bypass_regNext_22_0_data_3;
  reg                 io_in_r_bypass_regNext_22_0_load_store_3;
  reg                 io_in_r_bypass_regNext_22_0_df_is_ws_3;
  reg                 io_in_r_bypass_regNext_22_0_stall_3;
  reg        [15:0]   io_in_r_bypass_regNext_22_1_data_3;
  reg                 io_in_r_bypass_regNext_22_1_load_store_3;
  reg                 io_in_r_bypass_regNext_22_1_df_is_ws_3;
  reg                 io_in_r_bypass_regNext_22_1_stall_3;
  reg        [15:0]   io_in_r_bypass_regNext_22_2_data_3;
  reg                 io_in_r_bypass_regNext_22_2_load_store_3;
  reg                 io_in_r_bypass_regNext_22_2_df_is_ws_3;
  reg                 io_in_r_bypass_regNext_22_2_stall_3;
  reg        [15:0]   io_in_r_bypass_regNext_22_3_data_3;
  reg                 io_in_r_bypass_regNext_22_3_load_store_3;
  reg                 io_in_r_bypass_regNext_22_3_df_is_ws_3;
  reg                 io_in_r_bypass_regNext_22_3_stall_3;
  reg        [15:0]   io_in_r_bypass_regNext_23_0_data_3;
  reg                 io_in_r_bypass_regNext_23_0_load_store_3;
  reg                 io_in_r_bypass_regNext_23_0_df_is_ws_3;
  reg                 io_in_r_bypass_regNext_23_0_stall_3;
  reg        [15:0]   io_in_r_bypass_regNext_23_1_data_3;
  reg                 io_in_r_bypass_regNext_23_1_load_store_3;
  reg                 io_in_r_bypass_regNext_23_1_df_is_ws_3;
  reg                 io_in_r_bypass_regNext_23_1_stall_3;
  reg        [15:0]   io_in_r_bypass_regNext_23_2_data_3;
  reg                 io_in_r_bypass_regNext_23_2_load_store_3;
  reg                 io_in_r_bypass_regNext_23_2_df_is_ws_3;
  reg                 io_in_r_bypass_regNext_23_2_stall_3;
  reg        [15:0]   io_in_r_bypass_regNext_23_3_data_3;
  reg                 io_in_r_bypass_regNext_23_3_load_store_3;
  reg                 io_in_r_bypass_regNext_23_3_df_is_ws_3;
  reg                 io_in_r_bypass_regNext_23_3_stall_3;
  reg        [15:0]   io_in_r_bypass_regNext_24_0_data_3;
  reg                 io_in_r_bypass_regNext_24_0_load_store_3;
  reg                 io_in_r_bypass_regNext_24_0_df_is_ws_3;
  reg                 io_in_r_bypass_regNext_24_0_stall_3;
  reg        [15:0]   io_in_r_bypass_regNext_24_1_data_3;
  reg                 io_in_r_bypass_regNext_24_1_load_store_3;
  reg                 io_in_r_bypass_regNext_24_1_df_is_ws_3;
  reg                 io_in_r_bypass_regNext_24_1_stall_3;
  reg        [15:0]   io_in_r_bypass_regNext_24_2_data_3;
  reg                 io_in_r_bypass_regNext_24_2_load_store_3;
  reg                 io_in_r_bypass_regNext_24_2_df_is_ws_3;
  reg                 io_in_r_bypass_regNext_24_2_stall_3;
  reg        [15:0]   io_in_r_bypass_regNext_24_3_data_3;
  reg                 io_in_r_bypass_regNext_24_3_load_store_3;
  reg                 io_in_r_bypass_regNext_24_3_df_is_ws_3;
  reg                 io_in_r_bypass_regNext_24_3_stall_3;
  reg        [15:0]   io_in_r_bypass_regNext_25_0_data_3;
  reg                 io_in_r_bypass_regNext_25_0_load_store_3;
  reg                 io_in_r_bypass_regNext_25_0_df_is_ws_3;
  reg                 io_in_r_bypass_regNext_25_0_stall_3;
  reg        [15:0]   io_in_r_bypass_regNext_25_1_data_3;
  reg                 io_in_r_bypass_regNext_25_1_load_store_3;
  reg                 io_in_r_bypass_regNext_25_1_df_is_ws_3;
  reg                 io_in_r_bypass_regNext_25_1_stall_3;
  reg        [15:0]   io_in_r_bypass_regNext_25_2_data_3;
  reg                 io_in_r_bypass_regNext_25_2_load_store_3;
  reg                 io_in_r_bypass_regNext_25_2_df_is_ws_3;
  reg                 io_in_r_bypass_regNext_25_2_stall_3;
  reg        [15:0]   io_in_r_bypass_regNext_25_3_data_3;
  reg                 io_in_r_bypass_regNext_25_3_load_store_3;
  reg                 io_in_r_bypass_regNext_25_3_df_is_ws_3;
  reg                 io_in_r_bypass_regNext_25_3_stall_3;
  reg        [15:0]   io_in_r_bypass_regNext_26_0_data_3;
  reg                 io_in_r_bypass_regNext_26_0_load_store_3;
  reg                 io_in_r_bypass_regNext_26_0_df_is_ws_3;
  reg                 io_in_r_bypass_regNext_26_0_stall_3;
  reg        [15:0]   io_in_r_bypass_regNext_26_1_data_3;
  reg                 io_in_r_bypass_regNext_26_1_load_store_3;
  reg                 io_in_r_bypass_regNext_26_1_df_is_ws_3;
  reg                 io_in_r_bypass_regNext_26_1_stall_3;
  reg        [15:0]   io_in_r_bypass_regNext_26_2_data_3;
  reg                 io_in_r_bypass_regNext_26_2_load_store_3;
  reg                 io_in_r_bypass_regNext_26_2_df_is_ws_3;
  reg                 io_in_r_bypass_regNext_26_2_stall_3;
  reg        [15:0]   io_in_r_bypass_regNext_26_3_data_3;
  reg                 io_in_r_bypass_regNext_26_3_load_store_3;
  reg                 io_in_r_bypass_regNext_26_3_df_is_ws_3;
  reg                 io_in_r_bypass_regNext_26_3_stall_3;
  reg        [15:0]   io_in_r_bypass_regNext_27_0_data_3;
  reg                 io_in_r_bypass_regNext_27_0_load_store_3;
  reg                 io_in_r_bypass_regNext_27_0_df_is_ws_3;
  reg                 io_in_r_bypass_regNext_27_0_stall_3;
  reg        [15:0]   io_in_r_bypass_regNext_27_1_data_3;
  reg                 io_in_r_bypass_regNext_27_1_load_store_3;
  reg                 io_in_r_bypass_regNext_27_1_df_is_ws_3;
  reg                 io_in_r_bypass_regNext_27_1_stall_3;
  reg        [15:0]   io_in_r_bypass_regNext_27_2_data_3;
  reg                 io_in_r_bypass_regNext_27_2_load_store_3;
  reg                 io_in_r_bypass_regNext_27_2_df_is_ws_3;
  reg                 io_in_r_bypass_regNext_27_2_stall_3;
  reg        [15:0]   io_in_r_bypass_regNext_27_3_data_3;
  reg                 io_in_r_bypass_regNext_27_3_load_store_3;
  reg                 io_in_r_bypass_regNext_27_3_df_is_ws_3;
  reg                 io_in_r_bypass_regNext_27_3_stall_3;
  reg        [15:0]   io_in_r_bypass_regNext_28_0_data_3;
  reg                 io_in_r_bypass_regNext_28_0_load_store_3;
  reg                 io_in_r_bypass_regNext_28_0_df_is_ws_3;
  reg                 io_in_r_bypass_regNext_28_0_stall_3;
  reg        [15:0]   io_in_r_bypass_regNext_28_1_data_3;
  reg                 io_in_r_bypass_regNext_28_1_load_store_3;
  reg                 io_in_r_bypass_regNext_28_1_df_is_ws_3;
  reg                 io_in_r_bypass_regNext_28_1_stall_3;
  reg        [15:0]   io_in_r_bypass_regNext_28_2_data_3;
  reg                 io_in_r_bypass_regNext_28_2_load_store_3;
  reg                 io_in_r_bypass_regNext_28_2_df_is_ws_3;
  reg                 io_in_r_bypass_regNext_28_2_stall_3;
  reg        [15:0]   io_in_r_bypass_regNext_28_3_data_3;
  reg                 io_in_r_bypass_regNext_28_3_load_store_3;
  reg                 io_in_r_bypass_regNext_28_3_df_is_ws_3;
  reg                 io_in_r_bypass_regNext_28_3_stall_3;
  reg        [15:0]   io_in_r_bypass_regNext_29_0_data_3;
  reg                 io_in_r_bypass_regNext_29_0_load_store_3;
  reg                 io_in_r_bypass_regNext_29_0_df_is_ws_3;
  reg                 io_in_r_bypass_regNext_29_0_stall_3;
  reg        [15:0]   io_in_r_bypass_regNext_29_1_data_3;
  reg                 io_in_r_bypass_regNext_29_1_load_store_3;
  reg                 io_in_r_bypass_regNext_29_1_df_is_ws_3;
  reg                 io_in_r_bypass_regNext_29_1_stall_3;
  reg        [15:0]   io_in_r_bypass_regNext_29_2_data_3;
  reg                 io_in_r_bypass_regNext_29_2_load_store_3;
  reg                 io_in_r_bypass_regNext_29_2_df_is_ws_3;
  reg                 io_in_r_bypass_regNext_29_2_stall_3;
  reg        [15:0]   io_in_r_bypass_regNext_29_3_data_3;
  reg                 io_in_r_bypass_regNext_29_3_load_store_3;
  reg                 io_in_r_bypass_regNext_29_3_df_is_ws_3;
  reg                 io_in_r_bypass_regNext_29_3_stall_3;
  reg        [15:0]   io_in_r_bypass_regNext_30_0_data_3;
  reg                 io_in_r_bypass_regNext_30_0_load_store_3;
  reg                 io_in_r_bypass_regNext_30_0_df_is_ws_3;
  reg                 io_in_r_bypass_regNext_30_0_stall_3;
  reg        [15:0]   io_in_r_bypass_regNext_30_1_data_3;
  reg                 io_in_r_bypass_regNext_30_1_load_store_3;
  reg                 io_in_r_bypass_regNext_30_1_df_is_ws_3;
  reg                 io_in_r_bypass_regNext_30_1_stall_3;
  reg        [15:0]   io_in_r_bypass_regNext_30_2_data_3;
  reg                 io_in_r_bypass_regNext_30_2_load_store_3;
  reg                 io_in_r_bypass_regNext_30_2_df_is_ws_3;
  reg                 io_in_r_bypass_regNext_30_2_stall_3;
  reg        [15:0]   io_in_r_bypass_regNext_30_3_data_3;
  reg                 io_in_r_bypass_regNext_30_3_load_store_3;
  reg                 io_in_r_bypass_regNext_30_3_df_is_ws_3;
  reg                 io_in_r_bypass_regNext_30_3_stall_3;
  reg        [15:0]   io_in_r_bypass_regNext_31_0_data_3;
  reg                 io_in_r_bypass_regNext_31_0_load_store_3;
  reg                 io_in_r_bypass_regNext_31_0_df_is_ws_3;
  reg                 io_in_r_bypass_regNext_31_0_stall_3;
  reg        [15:0]   io_in_r_bypass_regNext_31_1_data_3;
  reg                 io_in_r_bypass_regNext_31_1_load_store_3;
  reg                 io_in_r_bypass_regNext_31_1_df_is_ws_3;
  reg                 io_in_r_bypass_regNext_31_1_stall_3;
  reg        [15:0]   io_in_r_bypass_regNext_31_2_data_3;
  reg                 io_in_r_bypass_regNext_31_2_load_store_3;
  reg                 io_in_r_bypass_regNext_31_2_df_is_ws_3;
  reg                 io_in_r_bypass_regNext_31_2_stall_3;
  reg        [15:0]   io_in_r_bypass_regNext_31_3_data_3;
  reg                 io_in_r_bypass_regNext_31_3_load_store_3;
  reg                 io_in_r_bypass_regNext_31_3_df_is_ws_3;
  reg                 io_in_r_bypass_regNext_31_3_stall_3;
  reg        [15:0]   io_in_r_bypass_regNext_0_0_data_4;
  reg                 io_in_r_bypass_regNext_0_0_load_store_4;
  reg                 io_in_r_bypass_regNext_0_0_df_is_ws_4;
  reg                 io_in_r_bypass_regNext_0_0_stall_4;
  reg        [15:0]   io_in_r_bypass_regNext_0_1_data_4;
  reg                 io_in_r_bypass_regNext_0_1_load_store_4;
  reg                 io_in_r_bypass_regNext_0_1_df_is_ws_4;
  reg                 io_in_r_bypass_regNext_0_1_stall_4;
  reg        [15:0]   io_in_r_bypass_regNext_0_2_data_4;
  reg                 io_in_r_bypass_regNext_0_2_load_store_4;
  reg                 io_in_r_bypass_regNext_0_2_df_is_ws_4;
  reg                 io_in_r_bypass_regNext_0_2_stall_4;
  reg        [15:0]   io_in_r_bypass_regNext_0_3_data_4;
  reg                 io_in_r_bypass_regNext_0_3_load_store_4;
  reg                 io_in_r_bypass_regNext_0_3_df_is_ws_4;
  reg                 io_in_r_bypass_regNext_0_3_stall_4;
  reg        [15:0]   io_in_r_bypass_regNext_1_0_data_4;
  reg                 io_in_r_bypass_regNext_1_0_load_store_4;
  reg                 io_in_r_bypass_regNext_1_0_df_is_ws_4;
  reg                 io_in_r_bypass_regNext_1_0_stall_4;
  reg        [15:0]   io_in_r_bypass_regNext_1_1_data_4;
  reg                 io_in_r_bypass_regNext_1_1_load_store_4;
  reg                 io_in_r_bypass_regNext_1_1_df_is_ws_4;
  reg                 io_in_r_bypass_regNext_1_1_stall_4;
  reg        [15:0]   io_in_r_bypass_regNext_1_2_data_4;
  reg                 io_in_r_bypass_regNext_1_2_load_store_4;
  reg                 io_in_r_bypass_regNext_1_2_df_is_ws_4;
  reg                 io_in_r_bypass_regNext_1_2_stall_4;
  reg        [15:0]   io_in_r_bypass_regNext_1_3_data_4;
  reg                 io_in_r_bypass_regNext_1_3_load_store_4;
  reg                 io_in_r_bypass_regNext_1_3_df_is_ws_4;
  reg                 io_in_r_bypass_regNext_1_3_stall_4;
  reg        [15:0]   io_in_r_bypass_regNext_2_0_data_4;
  reg                 io_in_r_bypass_regNext_2_0_load_store_4;
  reg                 io_in_r_bypass_regNext_2_0_df_is_ws_4;
  reg                 io_in_r_bypass_regNext_2_0_stall_4;
  reg        [15:0]   io_in_r_bypass_regNext_2_1_data_4;
  reg                 io_in_r_bypass_regNext_2_1_load_store_4;
  reg                 io_in_r_bypass_regNext_2_1_df_is_ws_4;
  reg                 io_in_r_bypass_regNext_2_1_stall_4;
  reg        [15:0]   io_in_r_bypass_regNext_2_2_data_4;
  reg                 io_in_r_bypass_regNext_2_2_load_store_4;
  reg                 io_in_r_bypass_regNext_2_2_df_is_ws_4;
  reg                 io_in_r_bypass_regNext_2_2_stall_4;
  reg        [15:0]   io_in_r_bypass_regNext_2_3_data_4;
  reg                 io_in_r_bypass_regNext_2_3_load_store_4;
  reg                 io_in_r_bypass_regNext_2_3_df_is_ws_4;
  reg                 io_in_r_bypass_regNext_2_3_stall_4;
  reg        [15:0]   io_in_r_bypass_regNext_3_0_data_4;
  reg                 io_in_r_bypass_regNext_3_0_load_store_4;
  reg                 io_in_r_bypass_regNext_3_0_df_is_ws_4;
  reg                 io_in_r_bypass_regNext_3_0_stall_4;
  reg        [15:0]   io_in_r_bypass_regNext_3_1_data_4;
  reg                 io_in_r_bypass_regNext_3_1_load_store_4;
  reg                 io_in_r_bypass_regNext_3_1_df_is_ws_4;
  reg                 io_in_r_bypass_regNext_3_1_stall_4;
  reg        [15:0]   io_in_r_bypass_regNext_3_2_data_4;
  reg                 io_in_r_bypass_regNext_3_2_load_store_4;
  reg                 io_in_r_bypass_regNext_3_2_df_is_ws_4;
  reg                 io_in_r_bypass_regNext_3_2_stall_4;
  reg        [15:0]   io_in_r_bypass_regNext_3_3_data_4;
  reg                 io_in_r_bypass_regNext_3_3_load_store_4;
  reg                 io_in_r_bypass_regNext_3_3_df_is_ws_4;
  reg                 io_in_r_bypass_regNext_3_3_stall_4;
  reg        [15:0]   io_in_r_bypass_regNext_4_0_data_4;
  reg                 io_in_r_bypass_regNext_4_0_load_store_4;
  reg                 io_in_r_bypass_regNext_4_0_df_is_ws_4;
  reg                 io_in_r_bypass_regNext_4_0_stall_4;
  reg        [15:0]   io_in_r_bypass_regNext_4_1_data_4;
  reg                 io_in_r_bypass_regNext_4_1_load_store_4;
  reg                 io_in_r_bypass_regNext_4_1_df_is_ws_4;
  reg                 io_in_r_bypass_regNext_4_1_stall_4;
  reg        [15:0]   io_in_r_bypass_regNext_4_2_data_4;
  reg                 io_in_r_bypass_regNext_4_2_load_store_4;
  reg                 io_in_r_bypass_regNext_4_2_df_is_ws_4;
  reg                 io_in_r_bypass_regNext_4_2_stall_4;
  reg        [15:0]   io_in_r_bypass_regNext_4_3_data_4;
  reg                 io_in_r_bypass_regNext_4_3_load_store_4;
  reg                 io_in_r_bypass_regNext_4_3_df_is_ws_4;
  reg                 io_in_r_bypass_regNext_4_3_stall_4;
  reg        [15:0]   io_in_r_bypass_regNext_5_0_data_4;
  reg                 io_in_r_bypass_regNext_5_0_load_store_4;
  reg                 io_in_r_bypass_regNext_5_0_df_is_ws_4;
  reg                 io_in_r_bypass_regNext_5_0_stall_4;
  reg        [15:0]   io_in_r_bypass_regNext_5_1_data_4;
  reg                 io_in_r_bypass_regNext_5_1_load_store_4;
  reg                 io_in_r_bypass_regNext_5_1_df_is_ws_4;
  reg                 io_in_r_bypass_regNext_5_1_stall_4;
  reg        [15:0]   io_in_r_bypass_regNext_5_2_data_4;
  reg                 io_in_r_bypass_regNext_5_2_load_store_4;
  reg                 io_in_r_bypass_regNext_5_2_df_is_ws_4;
  reg                 io_in_r_bypass_regNext_5_2_stall_4;
  reg        [15:0]   io_in_r_bypass_regNext_5_3_data_4;
  reg                 io_in_r_bypass_regNext_5_3_load_store_4;
  reg                 io_in_r_bypass_regNext_5_3_df_is_ws_4;
  reg                 io_in_r_bypass_regNext_5_3_stall_4;
  reg        [15:0]   io_in_r_bypass_regNext_6_0_data_4;
  reg                 io_in_r_bypass_regNext_6_0_load_store_4;
  reg                 io_in_r_bypass_regNext_6_0_df_is_ws_4;
  reg                 io_in_r_bypass_regNext_6_0_stall_4;
  reg        [15:0]   io_in_r_bypass_regNext_6_1_data_4;
  reg                 io_in_r_bypass_regNext_6_1_load_store_4;
  reg                 io_in_r_bypass_regNext_6_1_df_is_ws_4;
  reg                 io_in_r_bypass_regNext_6_1_stall_4;
  reg        [15:0]   io_in_r_bypass_regNext_6_2_data_4;
  reg                 io_in_r_bypass_regNext_6_2_load_store_4;
  reg                 io_in_r_bypass_regNext_6_2_df_is_ws_4;
  reg                 io_in_r_bypass_regNext_6_2_stall_4;
  reg        [15:0]   io_in_r_bypass_regNext_6_3_data_4;
  reg                 io_in_r_bypass_regNext_6_3_load_store_4;
  reg                 io_in_r_bypass_regNext_6_3_df_is_ws_4;
  reg                 io_in_r_bypass_regNext_6_3_stall_4;
  reg        [15:0]   io_in_r_bypass_regNext_7_0_data_4;
  reg                 io_in_r_bypass_regNext_7_0_load_store_4;
  reg                 io_in_r_bypass_regNext_7_0_df_is_ws_4;
  reg                 io_in_r_bypass_regNext_7_0_stall_4;
  reg        [15:0]   io_in_r_bypass_regNext_7_1_data_4;
  reg                 io_in_r_bypass_regNext_7_1_load_store_4;
  reg                 io_in_r_bypass_regNext_7_1_df_is_ws_4;
  reg                 io_in_r_bypass_regNext_7_1_stall_4;
  reg        [15:0]   io_in_r_bypass_regNext_7_2_data_4;
  reg                 io_in_r_bypass_regNext_7_2_load_store_4;
  reg                 io_in_r_bypass_regNext_7_2_df_is_ws_4;
  reg                 io_in_r_bypass_regNext_7_2_stall_4;
  reg        [15:0]   io_in_r_bypass_regNext_7_3_data_4;
  reg                 io_in_r_bypass_regNext_7_3_load_store_4;
  reg                 io_in_r_bypass_regNext_7_3_df_is_ws_4;
  reg                 io_in_r_bypass_regNext_7_3_stall_4;
  reg        [15:0]   io_in_r_bypass_regNext_8_0_data_4;
  reg                 io_in_r_bypass_regNext_8_0_load_store_4;
  reg                 io_in_r_bypass_regNext_8_0_df_is_ws_4;
  reg                 io_in_r_bypass_regNext_8_0_stall_4;
  reg        [15:0]   io_in_r_bypass_regNext_8_1_data_4;
  reg                 io_in_r_bypass_regNext_8_1_load_store_4;
  reg                 io_in_r_bypass_regNext_8_1_df_is_ws_4;
  reg                 io_in_r_bypass_regNext_8_1_stall_4;
  reg        [15:0]   io_in_r_bypass_regNext_8_2_data_4;
  reg                 io_in_r_bypass_regNext_8_2_load_store_4;
  reg                 io_in_r_bypass_regNext_8_2_df_is_ws_4;
  reg                 io_in_r_bypass_regNext_8_2_stall_4;
  reg        [15:0]   io_in_r_bypass_regNext_8_3_data_4;
  reg                 io_in_r_bypass_regNext_8_3_load_store_4;
  reg                 io_in_r_bypass_regNext_8_3_df_is_ws_4;
  reg                 io_in_r_bypass_regNext_8_3_stall_4;
  reg        [15:0]   io_in_r_bypass_regNext_9_0_data_4;
  reg                 io_in_r_bypass_regNext_9_0_load_store_4;
  reg                 io_in_r_bypass_regNext_9_0_df_is_ws_4;
  reg                 io_in_r_bypass_regNext_9_0_stall_4;
  reg        [15:0]   io_in_r_bypass_regNext_9_1_data_4;
  reg                 io_in_r_bypass_regNext_9_1_load_store_4;
  reg                 io_in_r_bypass_regNext_9_1_df_is_ws_4;
  reg                 io_in_r_bypass_regNext_9_1_stall_4;
  reg        [15:0]   io_in_r_bypass_regNext_9_2_data_4;
  reg                 io_in_r_bypass_regNext_9_2_load_store_4;
  reg                 io_in_r_bypass_regNext_9_2_df_is_ws_4;
  reg                 io_in_r_bypass_regNext_9_2_stall_4;
  reg        [15:0]   io_in_r_bypass_regNext_9_3_data_4;
  reg                 io_in_r_bypass_regNext_9_3_load_store_4;
  reg                 io_in_r_bypass_regNext_9_3_df_is_ws_4;
  reg                 io_in_r_bypass_regNext_9_3_stall_4;
  reg        [15:0]   io_in_r_bypass_regNext_10_0_data_4;
  reg                 io_in_r_bypass_regNext_10_0_load_store_4;
  reg                 io_in_r_bypass_regNext_10_0_df_is_ws_4;
  reg                 io_in_r_bypass_regNext_10_0_stall_4;
  reg        [15:0]   io_in_r_bypass_regNext_10_1_data_4;
  reg                 io_in_r_bypass_regNext_10_1_load_store_4;
  reg                 io_in_r_bypass_regNext_10_1_df_is_ws_4;
  reg                 io_in_r_bypass_regNext_10_1_stall_4;
  reg        [15:0]   io_in_r_bypass_regNext_10_2_data_4;
  reg                 io_in_r_bypass_regNext_10_2_load_store_4;
  reg                 io_in_r_bypass_regNext_10_2_df_is_ws_4;
  reg                 io_in_r_bypass_regNext_10_2_stall_4;
  reg        [15:0]   io_in_r_bypass_regNext_10_3_data_4;
  reg                 io_in_r_bypass_regNext_10_3_load_store_4;
  reg                 io_in_r_bypass_regNext_10_3_df_is_ws_4;
  reg                 io_in_r_bypass_regNext_10_3_stall_4;
  reg        [15:0]   io_in_r_bypass_regNext_11_0_data_4;
  reg                 io_in_r_bypass_regNext_11_0_load_store_4;
  reg                 io_in_r_bypass_regNext_11_0_df_is_ws_4;
  reg                 io_in_r_bypass_regNext_11_0_stall_4;
  reg        [15:0]   io_in_r_bypass_regNext_11_1_data_4;
  reg                 io_in_r_bypass_regNext_11_1_load_store_4;
  reg                 io_in_r_bypass_regNext_11_1_df_is_ws_4;
  reg                 io_in_r_bypass_regNext_11_1_stall_4;
  reg        [15:0]   io_in_r_bypass_regNext_11_2_data_4;
  reg                 io_in_r_bypass_regNext_11_2_load_store_4;
  reg                 io_in_r_bypass_regNext_11_2_df_is_ws_4;
  reg                 io_in_r_bypass_regNext_11_2_stall_4;
  reg        [15:0]   io_in_r_bypass_regNext_11_3_data_4;
  reg                 io_in_r_bypass_regNext_11_3_load_store_4;
  reg                 io_in_r_bypass_regNext_11_3_df_is_ws_4;
  reg                 io_in_r_bypass_regNext_11_3_stall_4;
  reg        [15:0]   io_in_r_bypass_regNext_12_0_data_4;
  reg                 io_in_r_bypass_regNext_12_0_load_store_4;
  reg                 io_in_r_bypass_regNext_12_0_df_is_ws_4;
  reg                 io_in_r_bypass_regNext_12_0_stall_4;
  reg        [15:0]   io_in_r_bypass_regNext_12_1_data_4;
  reg                 io_in_r_bypass_regNext_12_1_load_store_4;
  reg                 io_in_r_bypass_regNext_12_1_df_is_ws_4;
  reg                 io_in_r_bypass_regNext_12_1_stall_4;
  reg        [15:0]   io_in_r_bypass_regNext_12_2_data_4;
  reg                 io_in_r_bypass_regNext_12_2_load_store_4;
  reg                 io_in_r_bypass_regNext_12_2_df_is_ws_4;
  reg                 io_in_r_bypass_regNext_12_2_stall_4;
  reg        [15:0]   io_in_r_bypass_regNext_12_3_data_4;
  reg                 io_in_r_bypass_regNext_12_3_load_store_4;
  reg                 io_in_r_bypass_regNext_12_3_df_is_ws_4;
  reg                 io_in_r_bypass_regNext_12_3_stall_4;
  reg        [15:0]   io_in_r_bypass_regNext_13_0_data_4;
  reg                 io_in_r_bypass_regNext_13_0_load_store_4;
  reg                 io_in_r_bypass_regNext_13_0_df_is_ws_4;
  reg                 io_in_r_bypass_regNext_13_0_stall_4;
  reg        [15:0]   io_in_r_bypass_regNext_13_1_data_4;
  reg                 io_in_r_bypass_regNext_13_1_load_store_4;
  reg                 io_in_r_bypass_regNext_13_1_df_is_ws_4;
  reg                 io_in_r_bypass_regNext_13_1_stall_4;
  reg        [15:0]   io_in_r_bypass_regNext_13_2_data_4;
  reg                 io_in_r_bypass_regNext_13_2_load_store_4;
  reg                 io_in_r_bypass_regNext_13_2_df_is_ws_4;
  reg                 io_in_r_bypass_regNext_13_2_stall_4;
  reg        [15:0]   io_in_r_bypass_regNext_13_3_data_4;
  reg                 io_in_r_bypass_regNext_13_3_load_store_4;
  reg                 io_in_r_bypass_regNext_13_3_df_is_ws_4;
  reg                 io_in_r_bypass_regNext_13_3_stall_4;
  reg        [15:0]   io_in_r_bypass_regNext_14_0_data_4;
  reg                 io_in_r_bypass_regNext_14_0_load_store_4;
  reg                 io_in_r_bypass_regNext_14_0_df_is_ws_4;
  reg                 io_in_r_bypass_regNext_14_0_stall_4;
  reg        [15:0]   io_in_r_bypass_regNext_14_1_data_4;
  reg                 io_in_r_bypass_regNext_14_1_load_store_4;
  reg                 io_in_r_bypass_regNext_14_1_df_is_ws_4;
  reg                 io_in_r_bypass_regNext_14_1_stall_4;
  reg        [15:0]   io_in_r_bypass_regNext_14_2_data_4;
  reg                 io_in_r_bypass_regNext_14_2_load_store_4;
  reg                 io_in_r_bypass_regNext_14_2_df_is_ws_4;
  reg                 io_in_r_bypass_regNext_14_2_stall_4;
  reg        [15:0]   io_in_r_bypass_regNext_14_3_data_4;
  reg                 io_in_r_bypass_regNext_14_3_load_store_4;
  reg                 io_in_r_bypass_regNext_14_3_df_is_ws_4;
  reg                 io_in_r_bypass_regNext_14_3_stall_4;
  reg        [15:0]   io_in_r_bypass_regNext_15_0_data_4;
  reg                 io_in_r_bypass_regNext_15_0_load_store_4;
  reg                 io_in_r_bypass_regNext_15_0_df_is_ws_4;
  reg                 io_in_r_bypass_regNext_15_0_stall_4;
  reg        [15:0]   io_in_r_bypass_regNext_15_1_data_4;
  reg                 io_in_r_bypass_regNext_15_1_load_store_4;
  reg                 io_in_r_bypass_regNext_15_1_df_is_ws_4;
  reg                 io_in_r_bypass_regNext_15_1_stall_4;
  reg        [15:0]   io_in_r_bypass_regNext_15_2_data_4;
  reg                 io_in_r_bypass_regNext_15_2_load_store_4;
  reg                 io_in_r_bypass_regNext_15_2_df_is_ws_4;
  reg                 io_in_r_bypass_regNext_15_2_stall_4;
  reg        [15:0]   io_in_r_bypass_regNext_15_3_data_4;
  reg                 io_in_r_bypass_regNext_15_3_load_store_4;
  reg                 io_in_r_bypass_regNext_15_3_df_is_ws_4;
  reg                 io_in_r_bypass_regNext_15_3_stall_4;
  reg        [15:0]   io_in_r_bypass_regNext_16_0_data_4;
  reg                 io_in_r_bypass_regNext_16_0_load_store_4;
  reg                 io_in_r_bypass_regNext_16_0_df_is_ws_4;
  reg                 io_in_r_bypass_regNext_16_0_stall_4;
  reg        [15:0]   io_in_r_bypass_regNext_16_1_data_4;
  reg                 io_in_r_bypass_regNext_16_1_load_store_4;
  reg                 io_in_r_bypass_regNext_16_1_df_is_ws_4;
  reg                 io_in_r_bypass_regNext_16_1_stall_4;
  reg        [15:0]   io_in_r_bypass_regNext_16_2_data_4;
  reg                 io_in_r_bypass_regNext_16_2_load_store_4;
  reg                 io_in_r_bypass_regNext_16_2_df_is_ws_4;
  reg                 io_in_r_bypass_regNext_16_2_stall_4;
  reg        [15:0]   io_in_r_bypass_regNext_16_3_data_4;
  reg                 io_in_r_bypass_regNext_16_3_load_store_4;
  reg                 io_in_r_bypass_regNext_16_3_df_is_ws_4;
  reg                 io_in_r_bypass_regNext_16_3_stall_4;
  reg        [15:0]   io_in_r_bypass_regNext_17_0_data_4;
  reg                 io_in_r_bypass_regNext_17_0_load_store_4;
  reg                 io_in_r_bypass_regNext_17_0_df_is_ws_4;
  reg                 io_in_r_bypass_regNext_17_0_stall_4;
  reg        [15:0]   io_in_r_bypass_regNext_17_1_data_4;
  reg                 io_in_r_bypass_regNext_17_1_load_store_4;
  reg                 io_in_r_bypass_regNext_17_1_df_is_ws_4;
  reg                 io_in_r_bypass_regNext_17_1_stall_4;
  reg        [15:0]   io_in_r_bypass_regNext_17_2_data_4;
  reg                 io_in_r_bypass_regNext_17_2_load_store_4;
  reg                 io_in_r_bypass_regNext_17_2_df_is_ws_4;
  reg                 io_in_r_bypass_regNext_17_2_stall_4;
  reg        [15:0]   io_in_r_bypass_regNext_17_3_data_4;
  reg                 io_in_r_bypass_regNext_17_3_load_store_4;
  reg                 io_in_r_bypass_regNext_17_3_df_is_ws_4;
  reg                 io_in_r_bypass_regNext_17_3_stall_4;
  reg        [15:0]   io_in_r_bypass_regNext_18_0_data_4;
  reg                 io_in_r_bypass_regNext_18_0_load_store_4;
  reg                 io_in_r_bypass_regNext_18_0_df_is_ws_4;
  reg                 io_in_r_bypass_regNext_18_0_stall_4;
  reg        [15:0]   io_in_r_bypass_regNext_18_1_data_4;
  reg                 io_in_r_bypass_regNext_18_1_load_store_4;
  reg                 io_in_r_bypass_regNext_18_1_df_is_ws_4;
  reg                 io_in_r_bypass_regNext_18_1_stall_4;
  reg        [15:0]   io_in_r_bypass_regNext_18_2_data_4;
  reg                 io_in_r_bypass_regNext_18_2_load_store_4;
  reg                 io_in_r_bypass_regNext_18_2_df_is_ws_4;
  reg                 io_in_r_bypass_regNext_18_2_stall_4;
  reg        [15:0]   io_in_r_bypass_regNext_18_3_data_4;
  reg                 io_in_r_bypass_regNext_18_3_load_store_4;
  reg                 io_in_r_bypass_regNext_18_3_df_is_ws_4;
  reg                 io_in_r_bypass_regNext_18_3_stall_4;
  reg        [15:0]   io_in_r_bypass_regNext_19_0_data_4;
  reg                 io_in_r_bypass_regNext_19_0_load_store_4;
  reg                 io_in_r_bypass_regNext_19_0_df_is_ws_4;
  reg                 io_in_r_bypass_regNext_19_0_stall_4;
  reg        [15:0]   io_in_r_bypass_regNext_19_1_data_4;
  reg                 io_in_r_bypass_regNext_19_1_load_store_4;
  reg                 io_in_r_bypass_regNext_19_1_df_is_ws_4;
  reg                 io_in_r_bypass_regNext_19_1_stall_4;
  reg        [15:0]   io_in_r_bypass_regNext_19_2_data_4;
  reg                 io_in_r_bypass_regNext_19_2_load_store_4;
  reg                 io_in_r_bypass_regNext_19_2_df_is_ws_4;
  reg                 io_in_r_bypass_regNext_19_2_stall_4;
  reg        [15:0]   io_in_r_bypass_regNext_19_3_data_4;
  reg                 io_in_r_bypass_regNext_19_3_load_store_4;
  reg                 io_in_r_bypass_regNext_19_3_df_is_ws_4;
  reg                 io_in_r_bypass_regNext_19_3_stall_4;
  reg        [15:0]   io_in_r_bypass_regNext_20_0_data_4;
  reg                 io_in_r_bypass_regNext_20_0_load_store_4;
  reg                 io_in_r_bypass_regNext_20_0_df_is_ws_4;
  reg                 io_in_r_bypass_regNext_20_0_stall_4;
  reg        [15:0]   io_in_r_bypass_regNext_20_1_data_4;
  reg                 io_in_r_bypass_regNext_20_1_load_store_4;
  reg                 io_in_r_bypass_regNext_20_1_df_is_ws_4;
  reg                 io_in_r_bypass_regNext_20_1_stall_4;
  reg        [15:0]   io_in_r_bypass_regNext_20_2_data_4;
  reg                 io_in_r_bypass_regNext_20_2_load_store_4;
  reg                 io_in_r_bypass_regNext_20_2_df_is_ws_4;
  reg                 io_in_r_bypass_regNext_20_2_stall_4;
  reg        [15:0]   io_in_r_bypass_regNext_20_3_data_4;
  reg                 io_in_r_bypass_regNext_20_3_load_store_4;
  reg                 io_in_r_bypass_regNext_20_3_df_is_ws_4;
  reg                 io_in_r_bypass_regNext_20_3_stall_4;
  reg        [15:0]   io_in_r_bypass_regNext_21_0_data_4;
  reg                 io_in_r_bypass_regNext_21_0_load_store_4;
  reg                 io_in_r_bypass_regNext_21_0_df_is_ws_4;
  reg                 io_in_r_bypass_regNext_21_0_stall_4;
  reg        [15:0]   io_in_r_bypass_regNext_21_1_data_4;
  reg                 io_in_r_bypass_regNext_21_1_load_store_4;
  reg                 io_in_r_bypass_regNext_21_1_df_is_ws_4;
  reg                 io_in_r_bypass_regNext_21_1_stall_4;
  reg        [15:0]   io_in_r_bypass_regNext_21_2_data_4;
  reg                 io_in_r_bypass_regNext_21_2_load_store_4;
  reg                 io_in_r_bypass_regNext_21_2_df_is_ws_4;
  reg                 io_in_r_bypass_regNext_21_2_stall_4;
  reg        [15:0]   io_in_r_bypass_regNext_21_3_data_4;
  reg                 io_in_r_bypass_regNext_21_3_load_store_4;
  reg                 io_in_r_bypass_regNext_21_3_df_is_ws_4;
  reg                 io_in_r_bypass_regNext_21_3_stall_4;
  reg        [15:0]   io_in_r_bypass_regNext_22_0_data_4;
  reg                 io_in_r_bypass_regNext_22_0_load_store_4;
  reg                 io_in_r_bypass_regNext_22_0_df_is_ws_4;
  reg                 io_in_r_bypass_regNext_22_0_stall_4;
  reg        [15:0]   io_in_r_bypass_regNext_22_1_data_4;
  reg                 io_in_r_bypass_regNext_22_1_load_store_4;
  reg                 io_in_r_bypass_regNext_22_1_df_is_ws_4;
  reg                 io_in_r_bypass_regNext_22_1_stall_4;
  reg        [15:0]   io_in_r_bypass_regNext_22_2_data_4;
  reg                 io_in_r_bypass_regNext_22_2_load_store_4;
  reg                 io_in_r_bypass_regNext_22_2_df_is_ws_4;
  reg                 io_in_r_bypass_regNext_22_2_stall_4;
  reg        [15:0]   io_in_r_bypass_regNext_22_3_data_4;
  reg                 io_in_r_bypass_regNext_22_3_load_store_4;
  reg                 io_in_r_bypass_regNext_22_3_df_is_ws_4;
  reg                 io_in_r_bypass_regNext_22_3_stall_4;
  reg        [15:0]   io_in_r_bypass_regNext_23_0_data_4;
  reg                 io_in_r_bypass_regNext_23_0_load_store_4;
  reg                 io_in_r_bypass_regNext_23_0_df_is_ws_4;
  reg                 io_in_r_bypass_regNext_23_0_stall_4;
  reg        [15:0]   io_in_r_bypass_regNext_23_1_data_4;
  reg                 io_in_r_bypass_regNext_23_1_load_store_4;
  reg                 io_in_r_bypass_regNext_23_1_df_is_ws_4;
  reg                 io_in_r_bypass_regNext_23_1_stall_4;
  reg        [15:0]   io_in_r_bypass_regNext_23_2_data_4;
  reg                 io_in_r_bypass_regNext_23_2_load_store_4;
  reg                 io_in_r_bypass_regNext_23_2_df_is_ws_4;
  reg                 io_in_r_bypass_regNext_23_2_stall_4;
  reg        [15:0]   io_in_r_bypass_regNext_23_3_data_4;
  reg                 io_in_r_bypass_regNext_23_3_load_store_4;
  reg                 io_in_r_bypass_regNext_23_3_df_is_ws_4;
  reg                 io_in_r_bypass_regNext_23_3_stall_4;
  reg        [15:0]   io_in_r_bypass_regNext_24_0_data_4;
  reg                 io_in_r_bypass_regNext_24_0_load_store_4;
  reg                 io_in_r_bypass_regNext_24_0_df_is_ws_4;
  reg                 io_in_r_bypass_regNext_24_0_stall_4;
  reg        [15:0]   io_in_r_bypass_regNext_24_1_data_4;
  reg                 io_in_r_bypass_regNext_24_1_load_store_4;
  reg                 io_in_r_bypass_regNext_24_1_df_is_ws_4;
  reg                 io_in_r_bypass_regNext_24_1_stall_4;
  reg        [15:0]   io_in_r_bypass_regNext_24_2_data_4;
  reg                 io_in_r_bypass_regNext_24_2_load_store_4;
  reg                 io_in_r_bypass_regNext_24_2_df_is_ws_4;
  reg                 io_in_r_bypass_regNext_24_2_stall_4;
  reg        [15:0]   io_in_r_bypass_regNext_24_3_data_4;
  reg                 io_in_r_bypass_regNext_24_3_load_store_4;
  reg                 io_in_r_bypass_regNext_24_3_df_is_ws_4;
  reg                 io_in_r_bypass_regNext_24_3_stall_4;
  reg        [15:0]   io_in_r_bypass_regNext_25_0_data_4;
  reg                 io_in_r_bypass_regNext_25_0_load_store_4;
  reg                 io_in_r_bypass_regNext_25_0_df_is_ws_4;
  reg                 io_in_r_bypass_regNext_25_0_stall_4;
  reg        [15:0]   io_in_r_bypass_regNext_25_1_data_4;
  reg                 io_in_r_bypass_regNext_25_1_load_store_4;
  reg                 io_in_r_bypass_regNext_25_1_df_is_ws_4;
  reg                 io_in_r_bypass_regNext_25_1_stall_4;
  reg        [15:0]   io_in_r_bypass_regNext_25_2_data_4;
  reg                 io_in_r_bypass_regNext_25_2_load_store_4;
  reg                 io_in_r_bypass_regNext_25_2_df_is_ws_4;
  reg                 io_in_r_bypass_regNext_25_2_stall_4;
  reg        [15:0]   io_in_r_bypass_regNext_25_3_data_4;
  reg                 io_in_r_bypass_regNext_25_3_load_store_4;
  reg                 io_in_r_bypass_regNext_25_3_df_is_ws_4;
  reg                 io_in_r_bypass_regNext_25_3_stall_4;
  reg        [15:0]   io_in_r_bypass_regNext_26_0_data_4;
  reg                 io_in_r_bypass_regNext_26_0_load_store_4;
  reg                 io_in_r_bypass_regNext_26_0_df_is_ws_4;
  reg                 io_in_r_bypass_regNext_26_0_stall_4;
  reg        [15:0]   io_in_r_bypass_regNext_26_1_data_4;
  reg                 io_in_r_bypass_regNext_26_1_load_store_4;
  reg                 io_in_r_bypass_regNext_26_1_df_is_ws_4;
  reg                 io_in_r_bypass_regNext_26_1_stall_4;
  reg        [15:0]   io_in_r_bypass_regNext_26_2_data_4;
  reg                 io_in_r_bypass_regNext_26_2_load_store_4;
  reg                 io_in_r_bypass_regNext_26_2_df_is_ws_4;
  reg                 io_in_r_bypass_regNext_26_2_stall_4;
  reg        [15:0]   io_in_r_bypass_regNext_26_3_data_4;
  reg                 io_in_r_bypass_regNext_26_3_load_store_4;
  reg                 io_in_r_bypass_regNext_26_3_df_is_ws_4;
  reg                 io_in_r_bypass_regNext_26_3_stall_4;
  reg        [15:0]   io_in_r_bypass_regNext_27_0_data_4;
  reg                 io_in_r_bypass_regNext_27_0_load_store_4;
  reg                 io_in_r_bypass_regNext_27_0_df_is_ws_4;
  reg                 io_in_r_bypass_regNext_27_0_stall_4;
  reg        [15:0]   io_in_r_bypass_regNext_27_1_data_4;
  reg                 io_in_r_bypass_regNext_27_1_load_store_4;
  reg                 io_in_r_bypass_regNext_27_1_df_is_ws_4;
  reg                 io_in_r_bypass_regNext_27_1_stall_4;
  reg        [15:0]   io_in_r_bypass_regNext_27_2_data_4;
  reg                 io_in_r_bypass_regNext_27_2_load_store_4;
  reg                 io_in_r_bypass_regNext_27_2_df_is_ws_4;
  reg                 io_in_r_bypass_regNext_27_2_stall_4;
  reg        [15:0]   io_in_r_bypass_regNext_27_3_data_4;
  reg                 io_in_r_bypass_regNext_27_3_load_store_4;
  reg                 io_in_r_bypass_regNext_27_3_df_is_ws_4;
  reg                 io_in_r_bypass_regNext_27_3_stall_4;
  reg        [15:0]   io_in_r_bypass_regNext_28_0_data_4;
  reg                 io_in_r_bypass_regNext_28_0_load_store_4;
  reg                 io_in_r_bypass_regNext_28_0_df_is_ws_4;
  reg                 io_in_r_bypass_regNext_28_0_stall_4;
  reg        [15:0]   io_in_r_bypass_regNext_28_1_data_4;
  reg                 io_in_r_bypass_regNext_28_1_load_store_4;
  reg                 io_in_r_bypass_regNext_28_1_df_is_ws_4;
  reg                 io_in_r_bypass_regNext_28_1_stall_4;
  reg        [15:0]   io_in_r_bypass_regNext_28_2_data_4;
  reg                 io_in_r_bypass_regNext_28_2_load_store_4;
  reg                 io_in_r_bypass_regNext_28_2_df_is_ws_4;
  reg                 io_in_r_bypass_regNext_28_2_stall_4;
  reg        [15:0]   io_in_r_bypass_regNext_28_3_data_4;
  reg                 io_in_r_bypass_regNext_28_3_load_store_4;
  reg                 io_in_r_bypass_regNext_28_3_df_is_ws_4;
  reg                 io_in_r_bypass_regNext_28_3_stall_4;
  reg        [15:0]   io_in_r_bypass_regNext_29_0_data_4;
  reg                 io_in_r_bypass_regNext_29_0_load_store_4;
  reg                 io_in_r_bypass_regNext_29_0_df_is_ws_4;
  reg                 io_in_r_bypass_regNext_29_0_stall_4;
  reg        [15:0]   io_in_r_bypass_regNext_29_1_data_4;
  reg                 io_in_r_bypass_regNext_29_1_load_store_4;
  reg                 io_in_r_bypass_regNext_29_1_df_is_ws_4;
  reg                 io_in_r_bypass_regNext_29_1_stall_4;
  reg        [15:0]   io_in_r_bypass_regNext_29_2_data_4;
  reg                 io_in_r_bypass_regNext_29_2_load_store_4;
  reg                 io_in_r_bypass_regNext_29_2_df_is_ws_4;
  reg                 io_in_r_bypass_regNext_29_2_stall_4;
  reg        [15:0]   io_in_r_bypass_regNext_29_3_data_4;
  reg                 io_in_r_bypass_regNext_29_3_load_store_4;
  reg                 io_in_r_bypass_regNext_29_3_df_is_ws_4;
  reg                 io_in_r_bypass_regNext_29_3_stall_4;
  reg        [15:0]   io_in_r_bypass_regNext_30_0_data_4;
  reg                 io_in_r_bypass_regNext_30_0_load_store_4;
  reg                 io_in_r_bypass_regNext_30_0_df_is_ws_4;
  reg                 io_in_r_bypass_regNext_30_0_stall_4;
  reg        [15:0]   io_in_r_bypass_regNext_30_1_data_4;
  reg                 io_in_r_bypass_regNext_30_1_load_store_4;
  reg                 io_in_r_bypass_regNext_30_1_df_is_ws_4;
  reg                 io_in_r_bypass_regNext_30_1_stall_4;
  reg        [15:0]   io_in_r_bypass_regNext_30_2_data_4;
  reg                 io_in_r_bypass_regNext_30_2_load_store_4;
  reg                 io_in_r_bypass_regNext_30_2_df_is_ws_4;
  reg                 io_in_r_bypass_regNext_30_2_stall_4;
  reg        [15:0]   io_in_r_bypass_regNext_30_3_data_4;
  reg                 io_in_r_bypass_regNext_30_3_load_store_4;
  reg                 io_in_r_bypass_regNext_30_3_df_is_ws_4;
  reg                 io_in_r_bypass_regNext_30_3_stall_4;
  reg        [15:0]   io_in_r_bypass_regNext_31_0_data_4;
  reg                 io_in_r_bypass_regNext_31_0_load_store_4;
  reg                 io_in_r_bypass_regNext_31_0_df_is_ws_4;
  reg                 io_in_r_bypass_regNext_31_0_stall_4;
  reg        [15:0]   io_in_r_bypass_regNext_31_1_data_4;
  reg                 io_in_r_bypass_regNext_31_1_load_store_4;
  reg                 io_in_r_bypass_regNext_31_1_df_is_ws_4;
  reg                 io_in_r_bypass_regNext_31_1_stall_4;
  reg        [15:0]   io_in_r_bypass_regNext_31_2_data_4;
  reg                 io_in_r_bypass_regNext_31_2_load_store_4;
  reg                 io_in_r_bypass_regNext_31_2_df_is_ws_4;
  reg                 io_in_r_bypass_regNext_31_2_stall_4;
  reg        [15:0]   io_in_r_bypass_regNext_31_3_data_4;
  reg                 io_in_r_bypass_regNext_31_3_load_store_4;
  reg                 io_in_r_bypass_regNext_31_3_df_is_ws_4;
  reg                 io_in_r_bypass_regNext_31_3_stall_4;
  reg        [15:0]   io_in_r_bypass_regNext_0_0_data_5;
  reg                 io_in_r_bypass_regNext_0_0_load_store_5;
  reg                 io_in_r_bypass_regNext_0_0_df_is_ws_5;
  reg                 io_in_r_bypass_regNext_0_0_stall_5;
  reg        [15:0]   io_in_r_bypass_regNext_0_1_data_5;
  reg                 io_in_r_bypass_regNext_0_1_load_store_5;
  reg                 io_in_r_bypass_regNext_0_1_df_is_ws_5;
  reg                 io_in_r_bypass_regNext_0_1_stall_5;
  reg        [15:0]   io_in_r_bypass_regNext_0_2_data_5;
  reg                 io_in_r_bypass_regNext_0_2_load_store_5;
  reg                 io_in_r_bypass_regNext_0_2_df_is_ws_5;
  reg                 io_in_r_bypass_regNext_0_2_stall_5;
  reg        [15:0]   io_in_r_bypass_regNext_0_3_data_5;
  reg                 io_in_r_bypass_regNext_0_3_load_store_5;
  reg                 io_in_r_bypass_regNext_0_3_df_is_ws_5;
  reg                 io_in_r_bypass_regNext_0_3_stall_5;
  reg        [15:0]   io_in_r_bypass_regNext_1_0_data_5;
  reg                 io_in_r_bypass_regNext_1_0_load_store_5;
  reg                 io_in_r_bypass_regNext_1_0_df_is_ws_5;
  reg                 io_in_r_bypass_regNext_1_0_stall_5;
  reg        [15:0]   io_in_r_bypass_regNext_1_1_data_5;
  reg                 io_in_r_bypass_regNext_1_1_load_store_5;
  reg                 io_in_r_bypass_regNext_1_1_df_is_ws_5;
  reg                 io_in_r_bypass_regNext_1_1_stall_5;
  reg        [15:0]   io_in_r_bypass_regNext_1_2_data_5;
  reg                 io_in_r_bypass_regNext_1_2_load_store_5;
  reg                 io_in_r_bypass_regNext_1_2_df_is_ws_5;
  reg                 io_in_r_bypass_regNext_1_2_stall_5;
  reg        [15:0]   io_in_r_bypass_regNext_1_3_data_5;
  reg                 io_in_r_bypass_regNext_1_3_load_store_5;
  reg                 io_in_r_bypass_regNext_1_3_df_is_ws_5;
  reg                 io_in_r_bypass_regNext_1_3_stall_5;
  reg        [15:0]   io_in_r_bypass_regNext_2_0_data_5;
  reg                 io_in_r_bypass_regNext_2_0_load_store_5;
  reg                 io_in_r_bypass_regNext_2_0_df_is_ws_5;
  reg                 io_in_r_bypass_regNext_2_0_stall_5;
  reg        [15:0]   io_in_r_bypass_regNext_2_1_data_5;
  reg                 io_in_r_bypass_regNext_2_1_load_store_5;
  reg                 io_in_r_bypass_regNext_2_1_df_is_ws_5;
  reg                 io_in_r_bypass_regNext_2_1_stall_5;
  reg        [15:0]   io_in_r_bypass_regNext_2_2_data_5;
  reg                 io_in_r_bypass_regNext_2_2_load_store_5;
  reg                 io_in_r_bypass_regNext_2_2_df_is_ws_5;
  reg                 io_in_r_bypass_regNext_2_2_stall_5;
  reg        [15:0]   io_in_r_bypass_regNext_2_3_data_5;
  reg                 io_in_r_bypass_regNext_2_3_load_store_5;
  reg                 io_in_r_bypass_regNext_2_3_df_is_ws_5;
  reg                 io_in_r_bypass_regNext_2_3_stall_5;
  reg        [15:0]   io_in_r_bypass_regNext_3_0_data_5;
  reg                 io_in_r_bypass_regNext_3_0_load_store_5;
  reg                 io_in_r_bypass_regNext_3_0_df_is_ws_5;
  reg                 io_in_r_bypass_regNext_3_0_stall_5;
  reg        [15:0]   io_in_r_bypass_regNext_3_1_data_5;
  reg                 io_in_r_bypass_regNext_3_1_load_store_5;
  reg                 io_in_r_bypass_regNext_3_1_df_is_ws_5;
  reg                 io_in_r_bypass_regNext_3_1_stall_5;
  reg        [15:0]   io_in_r_bypass_regNext_3_2_data_5;
  reg                 io_in_r_bypass_regNext_3_2_load_store_5;
  reg                 io_in_r_bypass_regNext_3_2_df_is_ws_5;
  reg                 io_in_r_bypass_regNext_3_2_stall_5;
  reg        [15:0]   io_in_r_bypass_regNext_3_3_data_5;
  reg                 io_in_r_bypass_regNext_3_3_load_store_5;
  reg                 io_in_r_bypass_regNext_3_3_df_is_ws_5;
  reg                 io_in_r_bypass_regNext_3_3_stall_5;
  reg        [15:0]   io_in_r_bypass_regNext_4_0_data_5;
  reg                 io_in_r_bypass_regNext_4_0_load_store_5;
  reg                 io_in_r_bypass_regNext_4_0_df_is_ws_5;
  reg                 io_in_r_bypass_regNext_4_0_stall_5;
  reg        [15:0]   io_in_r_bypass_regNext_4_1_data_5;
  reg                 io_in_r_bypass_regNext_4_1_load_store_5;
  reg                 io_in_r_bypass_regNext_4_1_df_is_ws_5;
  reg                 io_in_r_bypass_regNext_4_1_stall_5;
  reg        [15:0]   io_in_r_bypass_regNext_4_2_data_5;
  reg                 io_in_r_bypass_regNext_4_2_load_store_5;
  reg                 io_in_r_bypass_regNext_4_2_df_is_ws_5;
  reg                 io_in_r_bypass_regNext_4_2_stall_5;
  reg        [15:0]   io_in_r_bypass_regNext_4_3_data_5;
  reg                 io_in_r_bypass_regNext_4_3_load_store_5;
  reg                 io_in_r_bypass_regNext_4_3_df_is_ws_5;
  reg                 io_in_r_bypass_regNext_4_3_stall_5;
  reg        [15:0]   io_in_r_bypass_regNext_5_0_data_5;
  reg                 io_in_r_bypass_regNext_5_0_load_store_5;
  reg                 io_in_r_bypass_regNext_5_0_df_is_ws_5;
  reg                 io_in_r_bypass_regNext_5_0_stall_5;
  reg        [15:0]   io_in_r_bypass_regNext_5_1_data_5;
  reg                 io_in_r_bypass_regNext_5_1_load_store_5;
  reg                 io_in_r_bypass_regNext_5_1_df_is_ws_5;
  reg                 io_in_r_bypass_regNext_5_1_stall_5;
  reg        [15:0]   io_in_r_bypass_regNext_5_2_data_5;
  reg                 io_in_r_bypass_regNext_5_2_load_store_5;
  reg                 io_in_r_bypass_regNext_5_2_df_is_ws_5;
  reg                 io_in_r_bypass_regNext_5_2_stall_5;
  reg        [15:0]   io_in_r_bypass_regNext_5_3_data_5;
  reg                 io_in_r_bypass_regNext_5_3_load_store_5;
  reg                 io_in_r_bypass_regNext_5_3_df_is_ws_5;
  reg                 io_in_r_bypass_regNext_5_3_stall_5;
  reg        [15:0]   io_in_r_bypass_regNext_6_0_data_5;
  reg                 io_in_r_bypass_regNext_6_0_load_store_5;
  reg                 io_in_r_bypass_regNext_6_0_df_is_ws_5;
  reg                 io_in_r_bypass_regNext_6_0_stall_5;
  reg        [15:0]   io_in_r_bypass_regNext_6_1_data_5;
  reg                 io_in_r_bypass_regNext_6_1_load_store_5;
  reg                 io_in_r_bypass_regNext_6_1_df_is_ws_5;
  reg                 io_in_r_bypass_regNext_6_1_stall_5;
  reg        [15:0]   io_in_r_bypass_regNext_6_2_data_5;
  reg                 io_in_r_bypass_regNext_6_2_load_store_5;
  reg                 io_in_r_bypass_regNext_6_2_df_is_ws_5;
  reg                 io_in_r_bypass_regNext_6_2_stall_5;
  reg        [15:0]   io_in_r_bypass_regNext_6_3_data_5;
  reg                 io_in_r_bypass_regNext_6_3_load_store_5;
  reg                 io_in_r_bypass_regNext_6_3_df_is_ws_5;
  reg                 io_in_r_bypass_regNext_6_3_stall_5;
  reg        [15:0]   io_in_r_bypass_regNext_7_0_data_5;
  reg                 io_in_r_bypass_regNext_7_0_load_store_5;
  reg                 io_in_r_bypass_regNext_7_0_df_is_ws_5;
  reg                 io_in_r_bypass_regNext_7_0_stall_5;
  reg        [15:0]   io_in_r_bypass_regNext_7_1_data_5;
  reg                 io_in_r_bypass_regNext_7_1_load_store_5;
  reg                 io_in_r_bypass_regNext_7_1_df_is_ws_5;
  reg                 io_in_r_bypass_regNext_7_1_stall_5;
  reg        [15:0]   io_in_r_bypass_regNext_7_2_data_5;
  reg                 io_in_r_bypass_regNext_7_2_load_store_5;
  reg                 io_in_r_bypass_regNext_7_2_df_is_ws_5;
  reg                 io_in_r_bypass_regNext_7_2_stall_5;
  reg        [15:0]   io_in_r_bypass_regNext_7_3_data_5;
  reg                 io_in_r_bypass_regNext_7_3_load_store_5;
  reg                 io_in_r_bypass_regNext_7_3_df_is_ws_5;
  reg                 io_in_r_bypass_regNext_7_3_stall_5;
  reg        [15:0]   io_in_r_bypass_regNext_8_0_data_5;
  reg                 io_in_r_bypass_regNext_8_0_load_store_5;
  reg                 io_in_r_bypass_regNext_8_0_df_is_ws_5;
  reg                 io_in_r_bypass_regNext_8_0_stall_5;
  reg        [15:0]   io_in_r_bypass_regNext_8_1_data_5;
  reg                 io_in_r_bypass_regNext_8_1_load_store_5;
  reg                 io_in_r_bypass_regNext_8_1_df_is_ws_5;
  reg                 io_in_r_bypass_regNext_8_1_stall_5;
  reg        [15:0]   io_in_r_bypass_regNext_8_2_data_5;
  reg                 io_in_r_bypass_regNext_8_2_load_store_5;
  reg                 io_in_r_bypass_regNext_8_2_df_is_ws_5;
  reg                 io_in_r_bypass_regNext_8_2_stall_5;
  reg        [15:0]   io_in_r_bypass_regNext_8_3_data_5;
  reg                 io_in_r_bypass_regNext_8_3_load_store_5;
  reg                 io_in_r_bypass_regNext_8_3_df_is_ws_5;
  reg                 io_in_r_bypass_regNext_8_3_stall_5;
  reg        [15:0]   io_in_r_bypass_regNext_9_0_data_5;
  reg                 io_in_r_bypass_regNext_9_0_load_store_5;
  reg                 io_in_r_bypass_regNext_9_0_df_is_ws_5;
  reg                 io_in_r_bypass_regNext_9_0_stall_5;
  reg        [15:0]   io_in_r_bypass_regNext_9_1_data_5;
  reg                 io_in_r_bypass_regNext_9_1_load_store_5;
  reg                 io_in_r_bypass_regNext_9_1_df_is_ws_5;
  reg                 io_in_r_bypass_regNext_9_1_stall_5;
  reg        [15:0]   io_in_r_bypass_regNext_9_2_data_5;
  reg                 io_in_r_bypass_regNext_9_2_load_store_5;
  reg                 io_in_r_bypass_regNext_9_2_df_is_ws_5;
  reg                 io_in_r_bypass_regNext_9_2_stall_5;
  reg        [15:0]   io_in_r_bypass_regNext_9_3_data_5;
  reg                 io_in_r_bypass_regNext_9_3_load_store_5;
  reg                 io_in_r_bypass_regNext_9_3_df_is_ws_5;
  reg                 io_in_r_bypass_regNext_9_3_stall_5;
  reg        [15:0]   io_in_r_bypass_regNext_10_0_data_5;
  reg                 io_in_r_bypass_regNext_10_0_load_store_5;
  reg                 io_in_r_bypass_regNext_10_0_df_is_ws_5;
  reg                 io_in_r_bypass_regNext_10_0_stall_5;
  reg        [15:0]   io_in_r_bypass_regNext_10_1_data_5;
  reg                 io_in_r_bypass_regNext_10_1_load_store_5;
  reg                 io_in_r_bypass_regNext_10_1_df_is_ws_5;
  reg                 io_in_r_bypass_regNext_10_1_stall_5;
  reg        [15:0]   io_in_r_bypass_regNext_10_2_data_5;
  reg                 io_in_r_bypass_regNext_10_2_load_store_5;
  reg                 io_in_r_bypass_regNext_10_2_df_is_ws_5;
  reg                 io_in_r_bypass_regNext_10_2_stall_5;
  reg        [15:0]   io_in_r_bypass_regNext_10_3_data_5;
  reg                 io_in_r_bypass_regNext_10_3_load_store_5;
  reg                 io_in_r_bypass_regNext_10_3_df_is_ws_5;
  reg                 io_in_r_bypass_regNext_10_3_stall_5;
  reg        [15:0]   io_in_r_bypass_regNext_11_0_data_5;
  reg                 io_in_r_bypass_regNext_11_0_load_store_5;
  reg                 io_in_r_bypass_regNext_11_0_df_is_ws_5;
  reg                 io_in_r_bypass_regNext_11_0_stall_5;
  reg        [15:0]   io_in_r_bypass_regNext_11_1_data_5;
  reg                 io_in_r_bypass_regNext_11_1_load_store_5;
  reg                 io_in_r_bypass_regNext_11_1_df_is_ws_5;
  reg                 io_in_r_bypass_regNext_11_1_stall_5;
  reg        [15:0]   io_in_r_bypass_regNext_11_2_data_5;
  reg                 io_in_r_bypass_regNext_11_2_load_store_5;
  reg                 io_in_r_bypass_regNext_11_2_df_is_ws_5;
  reg                 io_in_r_bypass_regNext_11_2_stall_5;
  reg        [15:0]   io_in_r_bypass_regNext_11_3_data_5;
  reg                 io_in_r_bypass_regNext_11_3_load_store_5;
  reg                 io_in_r_bypass_regNext_11_3_df_is_ws_5;
  reg                 io_in_r_bypass_regNext_11_3_stall_5;
  reg        [15:0]   io_in_r_bypass_regNext_12_0_data_5;
  reg                 io_in_r_bypass_regNext_12_0_load_store_5;
  reg                 io_in_r_bypass_regNext_12_0_df_is_ws_5;
  reg                 io_in_r_bypass_regNext_12_0_stall_5;
  reg        [15:0]   io_in_r_bypass_regNext_12_1_data_5;
  reg                 io_in_r_bypass_regNext_12_1_load_store_5;
  reg                 io_in_r_bypass_regNext_12_1_df_is_ws_5;
  reg                 io_in_r_bypass_regNext_12_1_stall_5;
  reg        [15:0]   io_in_r_bypass_regNext_12_2_data_5;
  reg                 io_in_r_bypass_regNext_12_2_load_store_5;
  reg                 io_in_r_bypass_regNext_12_2_df_is_ws_5;
  reg                 io_in_r_bypass_regNext_12_2_stall_5;
  reg        [15:0]   io_in_r_bypass_regNext_12_3_data_5;
  reg                 io_in_r_bypass_regNext_12_3_load_store_5;
  reg                 io_in_r_bypass_regNext_12_3_df_is_ws_5;
  reg                 io_in_r_bypass_regNext_12_3_stall_5;
  reg        [15:0]   io_in_r_bypass_regNext_13_0_data_5;
  reg                 io_in_r_bypass_regNext_13_0_load_store_5;
  reg                 io_in_r_bypass_regNext_13_0_df_is_ws_5;
  reg                 io_in_r_bypass_regNext_13_0_stall_5;
  reg        [15:0]   io_in_r_bypass_regNext_13_1_data_5;
  reg                 io_in_r_bypass_regNext_13_1_load_store_5;
  reg                 io_in_r_bypass_regNext_13_1_df_is_ws_5;
  reg                 io_in_r_bypass_regNext_13_1_stall_5;
  reg        [15:0]   io_in_r_bypass_regNext_13_2_data_5;
  reg                 io_in_r_bypass_regNext_13_2_load_store_5;
  reg                 io_in_r_bypass_regNext_13_2_df_is_ws_5;
  reg                 io_in_r_bypass_regNext_13_2_stall_5;
  reg        [15:0]   io_in_r_bypass_regNext_13_3_data_5;
  reg                 io_in_r_bypass_regNext_13_3_load_store_5;
  reg                 io_in_r_bypass_regNext_13_3_df_is_ws_5;
  reg                 io_in_r_bypass_regNext_13_3_stall_5;
  reg        [15:0]   io_in_r_bypass_regNext_14_0_data_5;
  reg                 io_in_r_bypass_regNext_14_0_load_store_5;
  reg                 io_in_r_bypass_regNext_14_0_df_is_ws_5;
  reg                 io_in_r_bypass_regNext_14_0_stall_5;
  reg        [15:0]   io_in_r_bypass_regNext_14_1_data_5;
  reg                 io_in_r_bypass_regNext_14_1_load_store_5;
  reg                 io_in_r_bypass_regNext_14_1_df_is_ws_5;
  reg                 io_in_r_bypass_regNext_14_1_stall_5;
  reg        [15:0]   io_in_r_bypass_regNext_14_2_data_5;
  reg                 io_in_r_bypass_regNext_14_2_load_store_5;
  reg                 io_in_r_bypass_regNext_14_2_df_is_ws_5;
  reg                 io_in_r_bypass_regNext_14_2_stall_5;
  reg        [15:0]   io_in_r_bypass_regNext_14_3_data_5;
  reg                 io_in_r_bypass_regNext_14_3_load_store_5;
  reg                 io_in_r_bypass_regNext_14_3_df_is_ws_5;
  reg                 io_in_r_bypass_regNext_14_3_stall_5;
  reg        [15:0]   io_in_r_bypass_regNext_15_0_data_5;
  reg                 io_in_r_bypass_regNext_15_0_load_store_5;
  reg                 io_in_r_bypass_regNext_15_0_df_is_ws_5;
  reg                 io_in_r_bypass_regNext_15_0_stall_5;
  reg        [15:0]   io_in_r_bypass_regNext_15_1_data_5;
  reg                 io_in_r_bypass_regNext_15_1_load_store_5;
  reg                 io_in_r_bypass_regNext_15_1_df_is_ws_5;
  reg                 io_in_r_bypass_regNext_15_1_stall_5;
  reg        [15:0]   io_in_r_bypass_regNext_15_2_data_5;
  reg                 io_in_r_bypass_regNext_15_2_load_store_5;
  reg                 io_in_r_bypass_regNext_15_2_df_is_ws_5;
  reg                 io_in_r_bypass_regNext_15_2_stall_5;
  reg        [15:0]   io_in_r_bypass_regNext_15_3_data_5;
  reg                 io_in_r_bypass_regNext_15_3_load_store_5;
  reg                 io_in_r_bypass_regNext_15_3_df_is_ws_5;
  reg                 io_in_r_bypass_regNext_15_3_stall_5;
  reg        [15:0]   io_in_r_bypass_regNext_16_0_data_5;
  reg                 io_in_r_bypass_regNext_16_0_load_store_5;
  reg                 io_in_r_bypass_regNext_16_0_df_is_ws_5;
  reg                 io_in_r_bypass_regNext_16_0_stall_5;
  reg        [15:0]   io_in_r_bypass_regNext_16_1_data_5;
  reg                 io_in_r_bypass_regNext_16_1_load_store_5;
  reg                 io_in_r_bypass_regNext_16_1_df_is_ws_5;
  reg                 io_in_r_bypass_regNext_16_1_stall_5;
  reg        [15:0]   io_in_r_bypass_regNext_16_2_data_5;
  reg                 io_in_r_bypass_regNext_16_2_load_store_5;
  reg                 io_in_r_bypass_regNext_16_2_df_is_ws_5;
  reg                 io_in_r_bypass_regNext_16_2_stall_5;
  reg        [15:0]   io_in_r_bypass_regNext_16_3_data_5;
  reg                 io_in_r_bypass_regNext_16_3_load_store_5;
  reg                 io_in_r_bypass_regNext_16_3_df_is_ws_5;
  reg                 io_in_r_bypass_regNext_16_3_stall_5;
  reg        [15:0]   io_in_r_bypass_regNext_17_0_data_5;
  reg                 io_in_r_bypass_regNext_17_0_load_store_5;
  reg                 io_in_r_bypass_regNext_17_0_df_is_ws_5;
  reg                 io_in_r_bypass_regNext_17_0_stall_5;
  reg        [15:0]   io_in_r_bypass_regNext_17_1_data_5;
  reg                 io_in_r_bypass_regNext_17_1_load_store_5;
  reg                 io_in_r_bypass_regNext_17_1_df_is_ws_5;
  reg                 io_in_r_bypass_regNext_17_1_stall_5;
  reg        [15:0]   io_in_r_bypass_regNext_17_2_data_5;
  reg                 io_in_r_bypass_regNext_17_2_load_store_5;
  reg                 io_in_r_bypass_regNext_17_2_df_is_ws_5;
  reg                 io_in_r_bypass_regNext_17_2_stall_5;
  reg        [15:0]   io_in_r_bypass_regNext_17_3_data_5;
  reg                 io_in_r_bypass_regNext_17_3_load_store_5;
  reg                 io_in_r_bypass_regNext_17_3_df_is_ws_5;
  reg                 io_in_r_bypass_regNext_17_3_stall_5;
  reg        [15:0]   io_in_r_bypass_regNext_18_0_data_5;
  reg                 io_in_r_bypass_regNext_18_0_load_store_5;
  reg                 io_in_r_bypass_regNext_18_0_df_is_ws_5;
  reg                 io_in_r_bypass_regNext_18_0_stall_5;
  reg        [15:0]   io_in_r_bypass_regNext_18_1_data_5;
  reg                 io_in_r_bypass_regNext_18_1_load_store_5;
  reg                 io_in_r_bypass_regNext_18_1_df_is_ws_5;
  reg                 io_in_r_bypass_regNext_18_1_stall_5;
  reg        [15:0]   io_in_r_bypass_regNext_18_2_data_5;
  reg                 io_in_r_bypass_regNext_18_2_load_store_5;
  reg                 io_in_r_bypass_regNext_18_2_df_is_ws_5;
  reg                 io_in_r_bypass_regNext_18_2_stall_5;
  reg        [15:0]   io_in_r_bypass_regNext_18_3_data_5;
  reg                 io_in_r_bypass_regNext_18_3_load_store_5;
  reg                 io_in_r_bypass_regNext_18_3_df_is_ws_5;
  reg                 io_in_r_bypass_regNext_18_3_stall_5;
  reg        [15:0]   io_in_r_bypass_regNext_19_0_data_5;
  reg                 io_in_r_bypass_regNext_19_0_load_store_5;
  reg                 io_in_r_bypass_regNext_19_0_df_is_ws_5;
  reg                 io_in_r_bypass_regNext_19_0_stall_5;
  reg        [15:0]   io_in_r_bypass_regNext_19_1_data_5;
  reg                 io_in_r_bypass_regNext_19_1_load_store_5;
  reg                 io_in_r_bypass_regNext_19_1_df_is_ws_5;
  reg                 io_in_r_bypass_regNext_19_1_stall_5;
  reg        [15:0]   io_in_r_bypass_regNext_19_2_data_5;
  reg                 io_in_r_bypass_regNext_19_2_load_store_5;
  reg                 io_in_r_bypass_regNext_19_2_df_is_ws_5;
  reg                 io_in_r_bypass_regNext_19_2_stall_5;
  reg        [15:0]   io_in_r_bypass_regNext_19_3_data_5;
  reg                 io_in_r_bypass_regNext_19_3_load_store_5;
  reg                 io_in_r_bypass_regNext_19_3_df_is_ws_5;
  reg                 io_in_r_bypass_regNext_19_3_stall_5;
  reg        [15:0]   io_in_r_bypass_regNext_20_0_data_5;
  reg                 io_in_r_bypass_regNext_20_0_load_store_5;
  reg                 io_in_r_bypass_regNext_20_0_df_is_ws_5;
  reg                 io_in_r_bypass_regNext_20_0_stall_5;
  reg        [15:0]   io_in_r_bypass_regNext_20_1_data_5;
  reg                 io_in_r_bypass_regNext_20_1_load_store_5;
  reg                 io_in_r_bypass_regNext_20_1_df_is_ws_5;
  reg                 io_in_r_bypass_regNext_20_1_stall_5;
  reg        [15:0]   io_in_r_bypass_regNext_20_2_data_5;
  reg                 io_in_r_bypass_regNext_20_2_load_store_5;
  reg                 io_in_r_bypass_regNext_20_2_df_is_ws_5;
  reg                 io_in_r_bypass_regNext_20_2_stall_5;
  reg        [15:0]   io_in_r_bypass_regNext_20_3_data_5;
  reg                 io_in_r_bypass_regNext_20_3_load_store_5;
  reg                 io_in_r_bypass_regNext_20_3_df_is_ws_5;
  reg                 io_in_r_bypass_regNext_20_3_stall_5;
  reg        [15:0]   io_in_r_bypass_regNext_21_0_data_5;
  reg                 io_in_r_bypass_regNext_21_0_load_store_5;
  reg                 io_in_r_bypass_regNext_21_0_df_is_ws_5;
  reg                 io_in_r_bypass_regNext_21_0_stall_5;
  reg        [15:0]   io_in_r_bypass_regNext_21_1_data_5;
  reg                 io_in_r_bypass_regNext_21_1_load_store_5;
  reg                 io_in_r_bypass_regNext_21_1_df_is_ws_5;
  reg                 io_in_r_bypass_regNext_21_1_stall_5;
  reg        [15:0]   io_in_r_bypass_regNext_21_2_data_5;
  reg                 io_in_r_bypass_regNext_21_2_load_store_5;
  reg                 io_in_r_bypass_regNext_21_2_df_is_ws_5;
  reg                 io_in_r_bypass_regNext_21_2_stall_5;
  reg        [15:0]   io_in_r_bypass_regNext_21_3_data_5;
  reg                 io_in_r_bypass_regNext_21_3_load_store_5;
  reg                 io_in_r_bypass_regNext_21_3_df_is_ws_5;
  reg                 io_in_r_bypass_regNext_21_3_stall_5;
  reg        [15:0]   io_in_r_bypass_regNext_22_0_data_5;
  reg                 io_in_r_bypass_regNext_22_0_load_store_5;
  reg                 io_in_r_bypass_regNext_22_0_df_is_ws_5;
  reg                 io_in_r_bypass_regNext_22_0_stall_5;
  reg        [15:0]   io_in_r_bypass_regNext_22_1_data_5;
  reg                 io_in_r_bypass_regNext_22_1_load_store_5;
  reg                 io_in_r_bypass_regNext_22_1_df_is_ws_5;
  reg                 io_in_r_bypass_regNext_22_1_stall_5;
  reg        [15:0]   io_in_r_bypass_regNext_22_2_data_5;
  reg                 io_in_r_bypass_regNext_22_2_load_store_5;
  reg                 io_in_r_bypass_regNext_22_2_df_is_ws_5;
  reg                 io_in_r_bypass_regNext_22_2_stall_5;
  reg        [15:0]   io_in_r_bypass_regNext_22_3_data_5;
  reg                 io_in_r_bypass_regNext_22_3_load_store_5;
  reg                 io_in_r_bypass_regNext_22_3_df_is_ws_5;
  reg                 io_in_r_bypass_regNext_22_3_stall_5;
  reg        [15:0]   io_in_r_bypass_regNext_23_0_data_5;
  reg                 io_in_r_bypass_regNext_23_0_load_store_5;
  reg                 io_in_r_bypass_regNext_23_0_df_is_ws_5;
  reg                 io_in_r_bypass_regNext_23_0_stall_5;
  reg        [15:0]   io_in_r_bypass_regNext_23_1_data_5;
  reg                 io_in_r_bypass_regNext_23_1_load_store_5;
  reg                 io_in_r_bypass_regNext_23_1_df_is_ws_5;
  reg                 io_in_r_bypass_regNext_23_1_stall_5;
  reg        [15:0]   io_in_r_bypass_regNext_23_2_data_5;
  reg                 io_in_r_bypass_regNext_23_2_load_store_5;
  reg                 io_in_r_bypass_regNext_23_2_df_is_ws_5;
  reg                 io_in_r_bypass_regNext_23_2_stall_5;
  reg        [15:0]   io_in_r_bypass_regNext_23_3_data_5;
  reg                 io_in_r_bypass_regNext_23_3_load_store_5;
  reg                 io_in_r_bypass_regNext_23_3_df_is_ws_5;
  reg                 io_in_r_bypass_regNext_23_3_stall_5;
  reg        [15:0]   io_in_r_bypass_regNext_24_0_data_5;
  reg                 io_in_r_bypass_regNext_24_0_load_store_5;
  reg                 io_in_r_bypass_regNext_24_0_df_is_ws_5;
  reg                 io_in_r_bypass_regNext_24_0_stall_5;
  reg        [15:0]   io_in_r_bypass_regNext_24_1_data_5;
  reg                 io_in_r_bypass_regNext_24_1_load_store_5;
  reg                 io_in_r_bypass_regNext_24_1_df_is_ws_5;
  reg                 io_in_r_bypass_regNext_24_1_stall_5;
  reg        [15:0]   io_in_r_bypass_regNext_24_2_data_5;
  reg                 io_in_r_bypass_regNext_24_2_load_store_5;
  reg                 io_in_r_bypass_regNext_24_2_df_is_ws_5;
  reg                 io_in_r_bypass_regNext_24_2_stall_5;
  reg        [15:0]   io_in_r_bypass_regNext_24_3_data_5;
  reg                 io_in_r_bypass_regNext_24_3_load_store_5;
  reg                 io_in_r_bypass_regNext_24_3_df_is_ws_5;
  reg                 io_in_r_bypass_regNext_24_3_stall_5;
  reg        [15:0]   io_in_r_bypass_regNext_25_0_data_5;
  reg                 io_in_r_bypass_regNext_25_0_load_store_5;
  reg                 io_in_r_bypass_regNext_25_0_df_is_ws_5;
  reg                 io_in_r_bypass_regNext_25_0_stall_5;
  reg        [15:0]   io_in_r_bypass_regNext_25_1_data_5;
  reg                 io_in_r_bypass_regNext_25_1_load_store_5;
  reg                 io_in_r_bypass_regNext_25_1_df_is_ws_5;
  reg                 io_in_r_bypass_regNext_25_1_stall_5;
  reg        [15:0]   io_in_r_bypass_regNext_25_2_data_5;
  reg                 io_in_r_bypass_regNext_25_2_load_store_5;
  reg                 io_in_r_bypass_regNext_25_2_df_is_ws_5;
  reg                 io_in_r_bypass_regNext_25_2_stall_5;
  reg        [15:0]   io_in_r_bypass_regNext_25_3_data_5;
  reg                 io_in_r_bypass_regNext_25_3_load_store_5;
  reg                 io_in_r_bypass_regNext_25_3_df_is_ws_5;
  reg                 io_in_r_bypass_regNext_25_3_stall_5;
  reg        [15:0]   io_in_r_bypass_regNext_26_0_data_5;
  reg                 io_in_r_bypass_regNext_26_0_load_store_5;
  reg                 io_in_r_bypass_regNext_26_0_df_is_ws_5;
  reg                 io_in_r_bypass_regNext_26_0_stall_5;
  reg        [15:0]   io_in_r_bypass_regNext_26_1_data_5;
  reg                 io_in_r_bypass_regNext_26_1_load_store_5;
  reg                 io_in_r_bypass_regNext_26_1_df_is_ws_5;
  reg                 io_in_r_bypass_regNext_26_1_stall_5;
  reg        [15:0]   io_in_r_bypass_regNext_26_2_data_5;
  reg                 io_in_r_bypass_regNext_26_2_load_store_5;
  reg                 io_in_r_bypass_regNext_26_2_df_is_ws_5;
  reg                 io_in_r_bypass_regNext_26_2_stall_5;
  reg        [15:0]   io_in_r_bypass_regNext_26_3_data_5;
  reg                 io_in_r_bypass_regNext_26_3_load_store_5;
  reg                 io_in_r_bypass_regNext_26_3_df_is_ws_5;
  reg                 io_in_r_bypass_regNext_26_3_stall_5;
  reg        [15:0]   io_in_r_bypass_regNext_27_0_data_5;
  reg                 io_in_r_bypass_regNext_27_0_load_store_5;
  reg                 io_in_r_bypass_regNext_27_0_df_is_ws_5;
  reg                 io_in_r_bypass_regNext_27_0_stall_5;
  reg        [15:0]   io_in_r_bypass_regNext_27_1_data_5;
  reg                 io_in_r_bypass_regNext_27_1_load_store_5;
  reg                 io_in_r_bypass_regNext_27_1_df_is_ws_5;
  reg                 io_in_r_bypass_regNext_27_1_stall_5;
  reg        [15:0]   io_in_r_bypass_regNext_27_2_data_5;
  reg                 io_in_r_bypass_regNext_27_2_load_store_5;
  reg                 io_in_r_bypass_regNext_27_2_df_is_ws_5;
  reg                 io_in_r_bypass_regNext_27_2_stall_5;
  reg        [15:0]   io_in_r_bypass_regNext_27_3_data_5;
  reg                 io_in_r_bypass_regNext_27_3_load_store_5;
  reg                 io_in_r_bypass_regNext_27_3_df_is_ws_5;
  reg                 io_in_r_bypass_regNext_27_3_stall_5;
  reg        [15:0]   io_in_r_bypass_regNext_28_0_data_5;
  reg                 io_in_r_bypass_regNext_28_0_load_store_5;
  reg                 io_in_r_bypass_regNext_28_0_df_is_ws_5;
  reg                 io_in_r_bypass_regNext_28_0_stall_5;
  reg        [15:0]   io_in_r_bypass_regNext_28_1_data_5;
  reg                 io_in_r_bypass_regNext_28_1_load_store_5;
  reg                 io_in_r_bypass_regNext_28_1_df_is_ws_5;
  reg                 io_in_r_bypass_regNext_28_1_stall_5;
  reg        [15:0]   io_in_r_bypass_regNext_28_2_data_5;
  reg                 io_in_r_bypass_regNext_28_2_load_store_5;
  reg                 io_in_r_bypass_regNext_28_2_df_is_ws_5;
  reg                 io_in_r_bypass_regNext_28_2_stall_5;
  reg        [15:0]   io_in_r_bypass_regNext_28_3_data_5;
  reg                 io_in_r_bypass_regNext_28_3_load_store_5;
  reg                 io_in_r_bypass_regNext_28_3_df_is_ws_5;
  reg                 io_in_r_bypass_regNext_28_3_stall_5;
  reg        [15:0]   io_in_r_bypass_regNext_29_0_data_5;
  reg                 io_in_r_bypass_regNext_29_0_load_store_5;
  reg                 io_in_r_bypass_regNext_29_0_df_is_ws_5;
  reg                 io_in_r_bypass_regNext_29_0_stall_5;
  reg        [15:0]   io_in_r_bypass_regNext_29_1_data_5;
  reg                 io_in_r_bypass_regNext_29_1_load_store_5;
  reg                 io_in_r_bypass_regNext_29_1_df_is_ws_5;
  reg                 io_in_r_bypass_regNext_29_1_stall_5;
  reg        [15:0]   io_in_r_bypass_regNext_29_2_data_5;
  reg                 io_in_r_bypass_regNext_29_2_load_store_5;
  reg                 io_in_r_bypass_regNext_29_2_df_is_ws_5;
  reg                 io_in_r_bypass_regNext_29_2_stall_5;
  reg        [15:0]   io_in_r_bypass_regNext_29_3_data_5;
  reg                 io_in_r_bypass_regNext_29_3_load_store_5;
  reg                 io_in_r_bypass_regNext_29_3_df_is_ws_5;
  reg                 io_in_r_bypass_regNext_29_3_stall_5;
  reg        [15:0]   io_in_r_bypass_regNext_30_0_data_5;
  reg                 io_in_r_bypass_regNext_30_0_load_store_5;
  reg                 io_in_r_bypass_regNext_30_0_df_is_ws_5;
  reg                 io_in_r_bypass_regNext_30_0_stall_5;
  reg        [15:0]   io_in_r_bypass_regNext_30_1_data_5;
  reg                 io_in_r_bypass_regNext_30_1_load_store_5;
  reg                 io_in_r_bypass_regNext_30_1_df_is_ws_5;
  reg                 io_in_r_bypass_regNext_30_1_stall_5;
  reg        [15:0]   io_in_r_bypass_regNext_30_2_data_5;
  reg                 io_in_r_bypass_regNext_30_2_load_store_5;
  reg                 io_in_r_bypass_regNext_30_2_df_is_ws_5;
  reg                 io_in_r_bypass_regNext_30_2_stall_5;
  reg        [15:0]   io_in_r_bypass_regNext_30_3_data_5;
  reg                 io_in_r_bypass_regNext_30_3_load_store_5;
  reg                 io_in_r_bypass_regNext_30_3_df_is_ws_5;
  reg                 io_in_r_bypass_regNext_30_3_stall_5;
  reg        [15:0]   io_in_r_bypass_regNext_31_0_data_5;
  reg                 io_in_r_bypass_regNext_31_0_load_store_5;
  reg                 io_in_r_bypass_regNext_31_0_df_is_ws_5;
  reg                 io_in_r_bypass_regNext_31_0_stall_5;
  reg        [15:0]   io_in_r_bypass_regNext_31_1_data_5;
  reg                 io_in_r_bypass_regNext_31_1_load_store_5;
  reg                 io_in_r_bypass_regNext_31_1_df_is_ws_5;
  reg                 io_in_r_bypass_regNext_31_1_stall_5;
  reg        [15:0]   io_in_r_bypass_regNext_31_2_data_5;
  reg                 io_in_r_bypass_regNext_31_2_load_store_5;
  reg                 io_in_r_bypass_regNext_31_2_df_is_ws_5;
  reg                 io_in_r_bypass_regNext_31_2_stall_5;
  reg        [15:0]   io_in_r_bypass_regNext_31_3_data_5;
  reg                 io_in_r_bypass_regNext_31_3_load_store_5;
  reg                 io_in_r_bypass_regNext_31_3_df_is_ws_5;
  reg                 io_in_r_bypass_regNext_31_3_stall_5;
  reg        [15:0]   io_in_r_bypass_regNext_0_0_data_6;
  reg                 io_in_r_bypass_regNext_0_0_load_store_6;
  reg                 io_in_r_bypass_regNext_0_0_df_is_ws_6;
  reg                 io_in_r_bypass_regNext_0_0_stall_6;
  reg        [15:0]   io_in_r_bypass_regNext_0_1_data_6;
  reg                 io_in_r_bypass_regNext_0_1_load_store_6;
  reg                 io_in_r_bypass_regNext_0_1_df_is_ws_6;
  reg                 io_in_r_bypass_regNext_0_1_stall_6;
  reg        [15:0]   io_in_r_bypass_regNext_0_2_data_6;
  reg                 io_in_r_bypass_regNext_0_2_load_store_6;
  reg                 io_in_r_bypass_regNext_0_2_df_is_ws_6;
  reg                 io_in_r_bypass_regNext_0_2_stall_6;
  reg        [15:0]   io_in_r_bypass_regNext_0_3_data_6;
  reg                 io_in_r_bypass_regNext_0_3_load_store_6;
  reg                 io_in_r_bypass_regNext_0_3_df_is_ws_6;
  reg                 io_in_r_bypass_regNext_0_3_stall_6;
  reg        [15:0]   io_in_r_bypass_regNext_1_0_data_6;
  reg                 io_in_r_bypass_regNext_1_0_load_store_6;
  reg                 io_in_r_bypass_regNext_1_0_df_is_ws_6;
  reg                 io_in_r_bypass_regNext_1_0_stall_6;
  reg        [15:0]   io_in_r_bypass_regNext_1_1_data_6;
  reg                 io_in_r_bypass_regNext_1_1_load_store_6;
  reg                 io_in_r_bypass_regNext_1_1_df_is_ws_6;
  reg                 io_in_r_bypass_regNext_1_1_stall_6;
  reg        [15:0]   io_in_r_bypass_regNext_1_2_data_6;
  reg                 io_in_r_bypass_regNext_1_2_load_store_6;
  reg                 io_in_r_bypass_regNext_1_2_df_is_ws_6;
  reg                 io_in_r_bypass_regNext_1_2_stall_6;
  reg        [15:0]   io_in_r_bypass_regNext_1_3_data_6;
  reg                 io_in_r_bypass_regNext_1_3_load_store_6;
  reg                 io_in_r_bypass_regNext_1_3_df_is_ws_6;
  reg                 io_in_r_bypass_regNext_1_3_stall_6;
  reg        [15:0]   io_in_r_bypass_regNext_2_0_data_6;
  reg                 io_in_r_bypass_regNext_2_0_load_store_6;
  reg                 io_in_r_bypass_regNext_2_0_df_is_ws_6;
  reg                 io_in_r_bypass_regNext_2_0_stall_6;
  reg        [15:0]   io_in_r_bypass_regNext_2_1_data_6;
  reg                 io_in_r_bypass_regNext_2_1_load_store_6;
  reg                 io_in_r_bypass_regNext_2_1_df_is_ws_6;
  reg                 io_in_r_bypass_regNext_2_1_stall_6;
  reg        [15:0]   io_in_r_bypass_regNext_2_2_data_6;
  reg                 io_in_r_bypass_regNext_2_2_load_store_6;
  reg                 io_in_r_bypass_regNext_2_2_df_is_ws_6;
  reg                 io_in_r_bypass_regNext_2_2_stall_6;
  reg        [15:0]   io_in_r_bypass_regNext_2_3_data_6;
  reg                 io_in_r_bypass_regNext_2_3_load_store_6;
  reg                 io_in_r_bypass_regNext_2_3_df_is_ws_6;
  reg                 io_in_r_bypass_regNext_2_3_stall_6;
  reg        [15:0]   io_in_r_bypass_regNext_3_0_data_6;
  reg                 io_in_r_bypass_regNext_3_0_load_store_6;
  reg                 io_in_r_bypass_regNext_3_0_df_is_ws_6;
  reg                 io_in_r_bypass_regNext_3_0_stall_6;
  reg        [15:0]   io_in_r_bypass_regNext_3_1_data_6;
  reg                 io_in_r_bypass_regNext_3_1_load_store_6;
  reg                 io_in_r_bypass_regNext_3_1_df_is_ws_6;
  reg                 io_in_r_bypass_regNext_3_1_stall_6;
  reg        [15:0]   io_in_r_bypass_regNext_3_2_data_6;
  reg                 io_in_r_bypass_regNext_3_2_load_store_6;
  reg                 io_in_r_bypass_regNext_3_2_df_is_ws_6;
  reg                 io_in_r_bypass_regNext_3_2_stall_6;
  reg        [15:0]   io_in_r_bypass_regNext_3_3_data_6;
  reg                 io_in_r_bypass_regNext_3_3_load_store_6;
  reg                 io_in_r_bypass_regNext_3_3_df_is_ws_6;
  reg                 io_in_r_bypass_regNext_3_3_stall_6;
  reg        [15:0]   io_in_r_bypass_regNext_4_0_data_6;
  reg                 io_in_r_bypass_regNext_4_0_load_store_6;
  reg                 io_in_r_bypass_regNext_4_0_df_is_ws_6;
  reg                 io_in_r_bypass_regNext_4_0_stall_6;
  reg        [15:0]   io_in_r_bypass_regNext_4_1_data_6;
  reg                 io_in_r_bypass_regNext_4_1_load_store_6;
  reg                 io_in_r_bypass_regNext_4_1_df_is_ws_6;
  reg                 io_in_r_bypass_regNext_4_1_stall_6;
  reg        [15:0]   io_in_r_bypass_regNext_4_2_data_6;
  reg                 io_in_r_bypass_regNext_4_2_load_store_6;
  reg                 io_in_r_bypass_regNext_4_2_df_is_ws_6;
  reg                 io_in_r_bypass_regNext_4_2_stall_6;
  reg        [15:0]   io_in_r_bypass_regNext_4_3_data_6;
  reg                 io_in_r_bypass_regNext_4_3_load_store_6;
  reg                 io_in_r_bypass_regNext_4_3_df_is_ws_6;
  reg                 io_in_r_bypass_regNext_4_3_stall_6;
  reg        [15:0]   io_in_r_bypass_regNext_5_0_data_6;
  reg                 io_in_r_bypass_regNext_5_0_load_store_6;
  reg                 io_in_r_bypass_regNext_5_0_df_is_ws_6;
  reg                 io_in_r_bypass_regNext_5_0_stall_6;
  reg        [15:0]   io_in_r_bypass_regNext_5_1_data_6;
  reg                 io_in_r_bypass_regNext_5_1_load_store_6;
  reg                 io_in_r_bypass_regNext_5_1_df_is_ws_6;
  reg                 io_in_r_bypass_regNext_5_1_stall_6;
  reg        [15:0]   io_in_r_bypass_regNext_5_2_data_6;
  reg                 io_in_r_bypass_regNext_5_2_load_store_6;
  reg                 io_in_r_bypass_regNext_5_2_df_is_ws_6;
  reg                 io_in_r_bypass_regNext_5_2_stall_6;
  reg        [15:0]   io_in_r_bypass_regNext_5_3_data_6;
  reg                 io_in_r_bypass_regNext_5_3_load_store_6;
  reg                 io_in_r_bypass_regNext_5_3_df_is_ws_6;
  reg                 io_in_r_bypass_regNext_5_3_stall_6;
  reg        [15:0]   io_in_r_bypass_regNext_6_0_data_6;
  reg                 io_in_r_bypass_regNext_6_0_load_store_6;
  reg                 io_in_r_bypass_regNext_6_0_df_is_ws_6;
  reg                 io_in_r_bypass_regNext_6_0_stall_6;
  reg        [15:0]   io_in_r_bypass_regNext_6_1_data_6;
  reg                 io_in_r_bypass_regNext_6_1_load_store_6;
  reg                 io_in_r_bypass_regNext_6_1_df_is_ws_6;
  reg                 io_in_r_bypass_regNext_6_1_stall_6;
  reg        [15:0]   io_in_r_bypass_regNext_6_2_data_6;
  reg                 io_in_r_bypass_regNext_6_2_load_store_6;
  reg                 io_in_r_bypass_regNext_6_2_df_is_ws_6;
  reg                 io_in_r_bypass_regNext_6_2_stall_6;
  reg        [15:0]   io_in_r_bypass_regNext_6_3_data_6;
  reg                 io_in_r_bypass_regNext_6_3_load_store_6;
  reg                 io_in_r_bypass_regNext_6_3_df_is_ws_6;
  reg                 io_in_r_bypass_regNext_6_3_stall_6;
  reg        [15:0]   io_in_r_bypass_regNext_7_0_data_6;
  reg                 io_in_r_bypass_regNext_7_0_load_store_6;
  reg                 io_in_r_bypass_regNext_7_0_df_is_ws_6;
  reg                 io_in_r_bypass_regNext_7_0_stall_6;
  reg        [15:0]   io_in_r_bypass_regNext_7_1_data_6;
  reg                 io_in_r_bypass_regNext_7_1_load_store_6;
  reg                 io_in_r_bypass_regNext_7_1_df_is_ws_6;
  reg                 io_in_r_bypass_regNext_7_1_stall_6;
  reg        [15:0]   io_in_r_bypass_regNext_7_2_data_6;
  reg                 io_in_r_bypass_regNext_7_2_load_store_6;
  reg                 io_in_r_bypass_regNext_7_2_df_is_ws_6;
  reg                 io_in_r_bypass_regNext_7_2_stall_6;
  reg        [15:0]   io_in_r_bypass_regNext_7_3_data_6;
  reg                 io_in_r_bypass_regNext_7_3_load_store_6;
  reg                 io_in_r_bypass_regNext_7_3_df_is_ws_6;
  reg                 io_in_r_bypass_regNext_7_3_stall_6;
  reg        [15:0]   io_in_r_bypass_regNext_8_0_data_6;
  reg                 io_in_r_bypass_regNext_8_0_load_store_6;
  reg                 io_in_r_bypass_regNext_8_0_df_is_ws_6;
  reg                 io_in_r_bypass_regNext_8_0_stall_6;
  reg        [15:0]   io_in_r_bypass_regNext_8_1_data_6;
  reg                 io_in_r_bypass_regNext_8_1_load_store_6;
  reg                 io_in_r_bypass_regNext_8_1_df_is_ws_6;
  reg                 io_in_r_bypass_regNext_8_1_stall_6;
  reg        [15:0]   io_in_r_bypass_regNext_8_2_data_6;
  reg                 io_in_r_bypass_regNext_8_2_load_store_6;
  reg                 io_in_r_bypass_regNext_8_2_df_is_ws_6;
  reg                 io_in_r_bypass_regNext_8_2_stall_6;
  reg        [15:0]   io_in_r_bypass_regNext_8_3_data_6;
  reg                 io_in_r_bypass_regNext_8_3_load_store_6;
  reg                 io_in_r_bypass_regNext_8_3_df_is_ws_6;
  reg                 io_in_r_bypass_regNext_8_3_stall_6;
  reg        [15:0]   io_in_r_bypass_regNext_9_0_data_6;
  reg                 io_in_r_bypass_regNext_9_0_load_store_6;
  reg                 io_in_r_bypass_regNext_9_0_df_is_ws_6;
  reg                 io_in_r_bypass_regNext_9_0_stall_6;
  reg        [15:0]   io_in_r_bypass_regNext_9_1_data_6;
  reg                 io_in_r_bypass_regNext_9_1_load_store_6;
  reg                 io_in_r_bypass_regNext_9_1_df_is_ws_6;
  reg                 io_in_r_bypass_regNext_9_1_stall_6;
  reg        [15:0]   io_in_r_bypass_regNext_9_2_data_6;
  reg                 io_in_r_bypass_regNext_9_2_load_store_6;
  reg                 io_in_r_bypass_regNext_9_2_df_is_ws_6;
  reg                 io_in_r_bypass_regNext_9_2_stall_6;
  reg        [15:0]   io_in_r_bypass_regNext_9_3_data_6;
  reg                 io_in_r_bypass_regNext_9_3_load_store_6;
  reg                 io_in_r_bypass_regNext_9_3_df_is_ws_6;
  reg                 io_in_r_bypass_regNext_9_3_stall_6;
  reg        [15:0]   io_in_r_bypass_regNext_10_0_data_6;
  reg                 io_in_r_bypass_regNext_10_0_load_store_6;
  reg                 io_in_r_bypass_regNext_10_0_df_is_ws_6;
  reg                 io_in_r_bypass_regNext_10_0_stall_6;
  reg        [15:0]   io_in_r_bypass_regNext_10_1_data_6;
  reg                 io_in_r_bypass_regNext_10_1_load_store_6;
  reg                 io_in_r_bypass_regNext_10_1_df_is_ws_6;
  reg                 io_in_r_bypass_regNext_10_1_stall_6;
  reg        [15:0]   io_in_r_bypass_regNext_10_2_data_6;
  reg                 io_in_r_bypass_regNext_10_2_load_store_6;
  reg                 io_in_r_bypass_regNext_10_2_df_is_ws_6;
  reg                 io_in_r_bypass_regNext_10_2_stall_6;
  reg        [15:0]   io_in_r_bypass_regNext_10_3_data_6;
  reg                 io_in_r_bypass_regNext_10_3_load_store_6;
  reg                 io_in_r_bypass_regNext_10_3_df_is_ws_6;
  reg                 io_in_r_bypass_regNext_10_3_stall_6;
  reg        [15:0]   io_in_r_bypass_regNext_11_0_data_6;
  reg                 io_in_r_bypass_regNext_11_0_load_store_6;
  reg                 io_in_r_bypass_regNext_11_0_df_is_ws_6;
  reg                 io_in_r_bypass_regNext_11_0_stall_6;
  reg        [15:0]   io_in_r_bypass_regNext_11_1_data_6;
  reg                 io_in_r_bypass_regNext_11_1_load_store_6;
  reg                 io_in_r_bypass_regNext_11_1_df_is_ws_6;
  reg                 io_in_r_bypass_regNext_11_1_stall_6;
  reg        [15:0]   io_in_r_bypass_regNext_11_2_data_6;
  reg                 io_in_r_bypass_regNext_11_2_load_store_6;
  reg                 io_in_r_bypass_regNext_11_2_df_is_ws_6;
  reg                 io_in_r_bypass_regNext_11_2_stall_6;
  reg        [15:0]   io_in_r_bypass_regNext_11_3_data_6;
  reg                 io_in_r_bypass_regNext_11_3_load_store_6;
  reg                 io_in_r_bypass_regNext_11_3_df_is_ws_6;
  reg                 io_in_r_bypass_regNext_11_3_stall_6;
  reg        [15:0]   io_in_r_bypass_regNext_12_0_data_6;
  reg                 io_in_r_bypass_regNext_12_0_load_store_6;
  reg                 io_in_r_bypass_regNext_12_0_df_is_ws_6;
  reg                 io_in_r_bypass_regNext_12_0_stall_6;
  reg        [15:0]   io_in_r_bypass_regNext_12_1_data_6;
  reg                 io_in_r_bypass_regNext_12_1_load_store_6;
  reg                 io_in_r_bypass_regNext_12_1_df_is_ws_6;
  reg                 io_in_r_bypass_regNext_12_1_stall_6;
  reg        [15:0]   io_in_r_bypass_regNext_12_2_data_6;
  reg                 io_in_r_bypass_regNext_12_2_load_store_6;
  reg                 io_in_r_bypass_regNext_12_2_df_is_ws_6;
  reg                 io_in_r_bypass_regNext_12_2_stall_6;
  reg        [15:0]   io_in_r_bypass_regNext_12_3_data_6;
  reg                 io_in_r_bypass_regNext_12_3_load_store_6;
  reg                 io_in_r_bypass_regNext_12_3_df_is_ws_6;
  reg                 io_in_r_bypass_regNext_12_3_stall_6;
  reg        [15:0]   io_in_r_bypass_regNext_13_0_data_6;
  reg                 io_in_r_bypass_regNext_13_0_load_store_6;
  reg                 io_in_r_bypass_regNext_13_0_df_is_ws_6;
  reg                 io_in_r_bypass_regNext_13_0_stall_6;
  reg        [15:0]   io_in_r_bypass_regNext_13_1_data_6;
  reg                 io_in_r_bypass_regNext_13_1_load_store_6;
  reg                 io_in_r_bypass_regNext_13_1_df_is_ws_6;
  reg                 io_in_r_bypass_regNext_13_1_stall_6;
  reg        [15:0]   io_in_r_bypass_regNext_13_2_data_6;
  reg                 io_in_r_bypass_regNext_13_2_load_store_6;
  reg                 io_in_r_bypass_regNext_13_2_df_is_ws_6;
  reg                 io_in_r_bypass_regNext_13_2_stall_6;
  reg        [15:0]   io_in_r_bypass_regNext_13_3_data_6;
  reg                 io_in_r_bypass_regNext_13_3_load_store_6;
  reg                 io_in_r_bypass_regNext_13_3_df_is_ws_6;
  reg                 io_in_r_bypass_regNext_13_3_stall_6;
  reg        [15:0]   io_in_r_bypass_regNext_14_0_data_6;
  reg                 io_in_r_bypass_regNext_14_0_load_store_6;
  reg                 io_in_r_bypass_regNext_14_0_df_is_ws_6;
  reg                 io_in_r_bypass_regNext_14_0_stall_6;
  reg        [15:0]   io_in_r_bypass_regNext_14_1_data_6;
  reg                 io_in_r_bypass_regNext_14_1_load_store_6;
  reg                 io_in_r_bypass_regNext_14_1_df_is_ws_6;
  reg                 io_in_r_bypass_regNext_14_1_stall_6;
  reg        [15:0]   io_in_r_bypass_regNext_14_2_data_6;
  reg                 io_in_r_bypass_regNext_14_2_load_store_6;
  reg                 io_in_r_bypass_regNext_14_2_df_is_ws_6;
  reg                 io_in_r_bypass_regNext_14_2_stall_6;
  reg        [15:0]   io_in_r_bypass_regNext_14_3_data_6;
  reg                 io_in_r_bypass_regNext_14_3_load_store_6;
  reg                 io_in_r_bypass_regNext_14_3_df_is_ws_6;
  reg                 io_in_r_bypass_regNext_14_3_stall_6;
  reg        [15:0]   io_in_r_bypass_regNext_15_0_data_6;
  reg                 io_in_r_bypass_regNext_15_0_load_store_6;
  reg                 io_in_r_bypass_regNext_15_0_df_is_ws_6;
  reg                 io_in_r_bypass_regNext_15_0_stall_6;
  reg        [15:0]   io_in_r_bypass_regNext_15_1_data_6;
  reg                 io_in_r_bypass_regNext_15_1_load_store_6;
  reg                 io_in_r_bypass_regNext_15_1_df_is_ws_6;
  reg                 io_in_r_bypass_regNext_15_1_stall_6;
  reg        [15:0]   io_in_r_bypass_regNext_15_2_data_6;
  reg                 io_in_r_bypass_regNext_15_2_load_store_6;
  reg                 io_in_r_bypass_regNext_15_2_df_is_ws_6;
  reg                 io_in_r_bypass_regNext_15_2_stall_6;
  reg        [15:0]   io_in_r_bypass_regNext_15_3_data_6;
  reg                 io_in_r_bypass_regNext_15_3_load_store_6;
  reg                 io_in_r_bypass_regNext_15_3_df_is_ws_6;
  reg                 io_in_r_bypass_regNext_15_3_stall_6;
  reg        [15:0]   io_in_r_bypass_regNext_16_0_data_6;
  reg                 io_in_r_bypass_regNext_16_0_load_store_6;
  reg                 io_in_r_bypass_regNext_16_0_df_is_ws_6;
  reg                 io_in_r_bypass_regNext_16_0_stall_6;
  reg        [15:0]   io_in_r_bypass_regNext_16_1_data_6;
  reg                 io_in_r_bypass_regNext_16_1_load_store_6;
  reg                 io_in_r_bypass_regNext_16_1_df_is_ws_6;
  reg                 io_in_r_bypass_regNext_16_1_stall_6;
  reg        [15:0]   io_in_r_bypass_regNext_16_2_data_6;
  reg                 io_in_r_bypass_regNext_16_2_load_store_6;
  reg                 io_in_r_bypass_regNext_16_2_df_is_ws_6;
  reg                 io_in_r_bypass_regNext_16_2_stall_6;
  reg        [15:0]   io_in_r_bypass_regNext_16_3_data_6;
  reg                 io_in_r_bypass_regNext_16_3_load_store_6;
  reg                 io_in_r_bypass_regNext_16_3_df_is_ws_6;
  reg                 io_in_r_bypass_regNext_16_3_stall_6;
  reg        [15:0]   io_in_r_bypass_regNext_17_0_data_6;
  reg                 io_in_r_bypass_regNext_17_0_load_store_6;
  reg                 io_in_r_bypass_regNext_17_0_df_is_ws_6;
  reg                 io_in_r_bypass_regNext_17_0_stall_6;
  reg        [15:0]   io_in_r_bypass_regNext_17_1_data_6;
  reg                 io_in_r_bypass_regNext_17_1_load_store_6;
  reg                 io_in_r_bypass_regNext_17_1_df_is_ws_6;
  reg                 io_in_r_bypass_regNext_17_1_stall_6;
  reg        [15:0]   io_in_r_bypass_regNext_17_2_data_6;
  reg                 io_in_r_bypass_regNext_17_2_load_store_6;
  reg                 io_in_r_bypass_regNext_17_2_df_is_ws_6;
  reg                 io_in_r_bypass_regNext_17_2_stall_6;
  reg        [15:0]   io_in_r_bypass_regNext_17_3_data_6;
  reg                 io_in_r_bypass_regNext_17_3_load_store_6;
  reg                 io_in_r_bypass_regNext_17_3_df_is_ws_6;
  reg                 io_in_r_bypass_regNext_17_3_stall_6;
  reg        [15:0]   io_in_r_bypass_regNext_18_0_data_6;
  reg                 io_in_r_bypass_regNext_18_0_load_store_6;
  reg                 io_in_r_bypass_regNext_18_0_df_is_ws_6;
  reg                 io_in_r_bypass_regNext_18_0_stall_6;
  reg        [15:0]   io_in_r_bypass_regNext_18_1_data_6;
  reg                 io_in_r_bypass_regNext_18_1_load_store_6;
  reg                 io_in_r_bypass_regNext_18_1_df_is_ws_6;
  reg                 io_in_r_bypass_regNext_18_1_stall_6;
  reg        [15:0]   io_in_r_bypass_regNext_18_2_data_6;
  reg                 io_in_r_bypass_regNext_18_2_load_store_6;
  reg                 io_in_r_bypass_regNext_18_2_df_is_ws_6;
  reg                 io_in_r_bypass_regNext_18_2_stall_6;
  reg        [15:0]   io_in_r_bypass_regNext_18_3_data_6;
  reg                 io_in_r_bypass_regNext_18_3_load_store_6;
  reg                 io_in_r_bypass_regNext_18_3_df_is_ws_6;
  reg                 io_in_r_bypass_regNext_18_3_stall_6;
  reg        [15:0]   io_in_r_bypass_regNext_19_0_data_6;
  reg                 io_in_r_bypass_regNext_19_0_load_store_6;
  reg                 io_in_r_bypass_regNext_19_0_df_is_ws_6;
  reg                 io_in_r_bypass_regNext_19_0_stall_6;
  reg        [15:0]   io_in_r_bypass_regNext_19_1_data_6;
  reg                 io_in_r_bypass_regNext_19_1_load_store_6;
  reg                 io_in_r_bypass_regNext_19_1_df_is_ws_6;
  reg                 io_in_r_bypass_regNext_19_1_stall_6;
  reg        [15:0]   io_in_r_bypass_regNext_19_2_data_6;
  reg                 io_in_r_bypass_regNext_19_2_load_store_6;
  reg                 io_in_r_bypass_regNext_19_2_df_is_ws_6;
  reg                 io_in_r_bypass_regNext_19_2_stall_6;
  reg        [15:0]   io_in_r_bypass_regNext_19_3_data_6;
  reg                 io_in_r_bypass_regNext_19_3_load_store_6;
  reg                 io_in_r_bypass_regNext_19_3_df_is_ws_6;
  reg                 io_in_r_bypass_regNext_19_3_stall_6;
  reg        [15:0]   io_in_r_bypass_regNext_20_0_data_6;
  reg                 io_in_r_bypass_regNext_20_0_load_store_6;
  reg                 io_in_r_bypass_regNext_20_0_df_is_ws_6;
  reg                 io_in_r_bypass_regNext_20_0_stall_6;
  reg        [15:0]   io_in_r_bypass_regNext_20_1_data_6;
  reg                 io_in_r_bypass_regNext_20_1_load_store_6;
  reg                 io_in_r_bypass_regNext_20_1_df_is_ws_6;
  reg                 io_in_r_bypass_regNext_20_1_stall_6;
  reg        [15:0]   io_in_r_bypass_regNext_20_2_data_6;
  reg                 io_in_r_bypass_regNext_20_2_load_store_6;
  reg                 io_in_r_bypass_regNext_20_2_df_is_ws_6;
  reg                 io_in_r_bypass_regNext_20_2_stall_6;
  reg        [15:0]   io_in_r_bypass_regNext_20_3_data_6;
  reg                 io_in_r_bypass_regNext_20_3_load_store_6;
  reg                 io_in_r_bypass_regNext_20_3_df_is_ws_6;
  reg                 io_in_r_bypass_regNext_20_3_stall_6;
  reg        [15:0]   io_in_r_bypass_regNext_21_0_data_6;
  reg                 io_in_r_bypass_regNext_21_0_load_store_6;
  reg                 io_in_r_bypass_regNext_21_0_df_is_ws_6;
  reg                 io_in_r_bypass_regNext_21_0_stall_6;
  reg        [15:0]   io_in_r_bypass_regNext_21_1_data_6;
  reg                 io_in_r_bypass_regNext_21_1_load_store_6;
  reg                 io_in_r_bypass_regNext_21_1_df_is_ws_6;
  reg                 io_in_r_bypass_regNext_21_1_stall_6;
  reg        [15:0]   io_in_r_bypass_regNext_21_2_data_6;
  reg                 io_in_r_bypass_regNext_21_2_load_store_6;
  reg                 io_in_r_bypass_regNext_21_2_df_is_ws_6;
  reg                 io_in_r_bypass_regNext_21_2_stall_6;
  reg        [15:0]   io_in_r_bypass_regNext_21_3_data_6;
  reg                 io_in_r_bypass_regNext_21_3_load_store_6;
  reg                 io_in_r_bypass_regNext_21_3_df_is_ws_6;
  reg                 io_in_r_bypass_regNext_21_3_stall_6;
  reg        [15:0]   io_in_r_bypass_regNext_22_0_data_6;
  reg                 io_in_r_bypass_regNext_22_0_load_store_6;
  reg                 io_in_r_bypass_regNext_22_0_df_is_ws_6;
  reg                 io_in_r_bypass_regNext_22_0_stall_6;
  reg        [15:0]   io_in_r_bypass_regNext_22_1_data_6;
  reg                 io_in_r_bypass_regNext_22_1_load_store_6;
  reg                 io_in_r_bypass_regNext_22_1_df_is_ws_6;
  reg                 io_in_r_bypass_regNext_22_1_stall_6;
  reg        [15:0]   io_in_r_bypass_regNext_22_2_data_6;
  reg                 io_in_r_bypass_regNext_22_2_load_store_6;
  reg                 io_in_r_bypass_regNext_22_2_df_is_ws_6;
  reg                 io_in_r_bypass_regNext_22_2_stall_6;
  reg        [15:0]   io_in_r_bypass_regNext_22_3_data_6;
  reg                 io_in_r_bypass_regNext_22_3_load_store_6;
  reg                 io_in_r_bypass_regNext_22_3_df_is_ws_6;
  reg                 io_in_r_bypass_regNext_22_3_stall_6;
  reg        [15:0]   io_in_r_bypass_regNext_23_0_data_6;
  reg                 io_in_r_bypass_regNext_23_0_load_store_6;
  reg                 io_in_r_bypass_regNext_23_0_df_is_ws_6;
  reg                 io_in_r_bypass_regNext_23_0_stall_6;
  reg        [15:0]   io_in_r_bypass_regNext_23_1_data_6;
  reg                 io_in_r_bypass_regNext_23_1_load_store_6;
  reg                 io_in_r_bypass_regNext_23_1_df_is_ws_6;
  reg                 io_in_r_bypass_regNext_23_1_stall_6;
  reg        [15:0]   io_in_r_bypass_regNext_23_2_data_6;
  reg                 io_in_r_bypass_regNext_23_2_load_store_6;
  reg                 io_in_r_bypass_regNext_23_2_df_is_ws_6;
  reg                 io_in_r_bypass_regNext_23_2_stall_6;
  reg        [15:0]   io_in_r_bypass_regNext_23_3_data_6;
  reg                 io_in_r_bypass_regNext_23_3_load_store_6;
  reg                 io_in_r_bypass_regNext_23_3_df_is_ws_6;
  reg                 io_in_r_bypass_regNext_23_3_stall_6;
  reg        [15:0]   io_in_r_bypass_regNext_24_0_data_6;
  reg                 io_in_r_bypass_regNext_24_0_load_store_6;
  reg                 io_in_r_bypass_regNext_24_0_df_is_ws_6;
  reg                 io_in_r_bypass_regNext_24_0_stall_6;
  reg        [15:0]   io_in_r_bypass_regNext_24_1_data_6;
  reg                 io_in_r_bypass_regNext_24_1_load_store_6;
  reg                 io_in_r_bypass_regNext_24_1_df_is_ws_6;
  reg                 io_in_r_bypass_regNext_24_1_stall_6;
  reg        [15:0]   io_in_r_bypass_regNext_24_2_data_6;
  reg                 io_in_r_bypass_regNext_24_2_load_store_6;
  reg                 io_in_r_bypass_regNext_24_2_df_is_ws_6;
  reg                 io_in_r_bypass_regNext_24_2_stall_6;
  reg        [15:0]   io_in_r_bypass_regNext_24_3_data_6;
  reg                 io_in_r_bypass_regNext_24_3_load_store_6;
  reg                 io_in_r_bypass_regNext_24_3_df_is_ws_6;
  reg                 io_in_r_bypass_regNext_24_3_stall_6;
  reg        [15:0]   io_in_r_bypass_regNext_25_0_data_6;
  reg                 io_in_r_bypass_regNext_25_0_load_store_6;
  reg                 io_in_r_bypass_regNext_25_0_df_is_ws_6;
  reg                 io_in_r_bypass_regNext_25_0_stall_6;
  reg        [15:0]   io_in_r_bypass_regNext_25_1_data_6;
  reg                 io_in_r_bypass_regNext_25_1_load_store_6;
  reg                 io_in_r_bypass_regNext_25_1_df_is_ws_6;
  reg                 io_in_r_bypass_regNext_25_1_stall_6;
  reg        [15:0]   io_in_r_bypass_regNext_25_2_data_6;
  reg                 io_in_r_bypass_regNext_25_2_load_store_6;
  reg                 io_in_r_bypass_regNext_25_2_df_is_ws_6;
  reg                 io_in_r_bypass_regNext_25_2_stall_6;
  reg        [15:0]   io_in_r_bypass_regNext_25_3_data_6;
  reg                 io_in_r_bypass_regNext_25_3_load_store_6;
  reg                 io_in_r_bypass_regNext_25_3_df_is_ws_6;
  reg                 io_in_r_bypass_regNext_25_3_stall_6;
  reg        [15:0]   io_in_r_bypass_regNext_26_0_data_6;
  reg                 io_in_r_bypass_regNext_26_0_load_store_6;
  reg                 io_in_r_bypass_regNext_26_0_df_is_ws_6;
  reg                 io_in_r_bypass_regNext_26_0_stall_6;
  reg        [15:0]   io_in_r_bypass_regNext_26_1_data_6;
  reg                 io_in_r_bypass_regNext_26_1_load_store_6;
  reg                 io_in_r_bypass_regNext_26_1_df_is_ws_6;
  reg                 io_in_r_bypass_regNext_26_1_stall_6;
  reg        [15:0]   io_in_r_bypass_regNext_26_2_data_6;
  reg                 io_in_r_bypass_regNext_26_2_load_store_6;
  reg                 io_in_r_bypass_regNext_26_2_df_is_ws_6;
  reg                 io_in_r_bypass_regNext_26_2_stall_6;
  reg        [15:0]   io_in_r_bypass_regNext_26_3_data_6;
  reg                 io_in_r_bypass_regNext_26_3_load_store_6;
  reg                 io_in_r_bypass_regNext_26_3_df_is_ws_6;
  reg                 io_in_r_bypass_regNext_26_3_stall_6;
  reg        [15:0]   io_in_r_bypass_regNext_27_0_data_6;
  reg                 io_in_r_bypass_regNext_27_0_load_store_6;
  reg                 io_in_r_bypass_regNext_27_0_df_is_ws_6;
  reg                 io_in_r_bypass_regNext_27_0_stall_6;
  reg        [15:0]   io_in_r_bypass_regNext_27_1_data_6;
  reg                 io_in_r_bypass_regNext_27_1_load_store_6;
  reg                 io_in_r_bypass_regNext_27_1_df_is_ws_6;
  reg                 io_in_r_bypass_regNext_27_1_stall_6;
  reg        [15:0]   io_in_r_bypass_regNext_27_2_data_6;
  reg                 io_in_r_bypass_regNext_27_2_load_store_6;
  reg                 io_in_r_bypass_regNext_27_2_df_is_ws_6;
  reg                 io_in_r_bypass_regNext_27_2_stall_6;
  reg        [15:0]   io_in_r_bypass_regNext_27_3_data_6;
  reg                 io_in_r_bypass_regNext_27_3_load_store_6;
  reg                 io_in_r_bypass_regNext_27_3_df_is_ws_6;
  reg                 io_in_r_bypass_regNext_27_3_stall_6;
  reg        [15:0]   io_in_r_bypass_regNext_28_0_data_6;
  reg                 io_in_r_bypass_regNext_28_0_load_store_6;
  reg                 io_in_r_bypass_regNext_28_0_df_is_ws_6;
  reg                 io_in_r_bypass_regNext_28_0_stall_6;
  reg        [15:0]   io_in_r_bypass_regNext_28_1_data_6;
  reg                 io_in_r_bypass_regNext_28_1_load_store_6;
  reg                 io_in_r_bypass_regNext_28_1_df_is_ws_6;
  reg                 io_in_r_bypass_regNext_28_1_stall_6;
  reg        [15:0]   io_in_r_bypass_regNext_28_2_data_6;
  reg                 io_in_r_bypass_regNext_28_2_load_store_6;
  reg                 io_in_r_bypass_regNext_28_2_df_is_ws_6;
  reg                 io_in_r_bypass_regNext_28_2_stall_6;
  reg        [15:0]   io_in_r_bypass_regNext_28_3_data_6;
  reg                 io_in_r_bypass_regNext_28_3_load_store_6;
  reg                 io_in_r_bypass_regNext_28_3_df_is_ws_6;
  reg                 io_in_r_bypass_regNext_28_3_stall_6;
  reg        [15:0]   io_in_r_bypass_regNext_29_0_data_6;
  reg                 io_in_r_bypass_regNext_29_0_load_store_6;
  reg                 io_in_r_bypass_regNext_29_0_df_is_ws_6;
  reg                 io_in_r_bypass_regNext_29_0_stall_6;
  reg        [15:0]   io_in_r_bypass_regNext_29_1_data_6;
  reg                 io_in_r_bypass_regNext_29_1_load_store_6;
  reg                 io_in_r_bypass_regNext_29_1_df_is_ws_6;
  reg                 io_in_r_bypass_regNext_29_1_stall_6;
  reg        [15:0]   io_in_r_bypass_regNext_29_2_data_6;
  reg                 io_in_r_bypass_regNext_29_2_load_store_6;
  reg                 io_in_r_bypass_regNext_29_2_df_is_ws_6;
  reg                 io_in_r_bypass_regNext_29_2_stall_6;
  reg        [15:0]   io_in_r_bypass_regNext_29_3_data_6;
  reg                 io_in_r_bypass_regNext_29_3_load_store_6;
  reg                 io_in_r_bypass_regNext_29_3_df_is_ws_6;
  reg                 io_in_r_bypass_regNext_29_3_stall_6;
  reg        [15:0]   io_in_r_bypass_regNext_30_0_data_6;
  reg                 io_in_r_bypass_regNext_30_0_load_store_6;
  reg                 io_in_r_bypass_regNext_30_0_df_is_ws_6;
  reg                 io_in_r_bypass_regNext_30_0_stall_6;
  reg        [15:0]   io_in_r_bypass_regNext_30_1_data_6;
  reg                 io_in_r_bypass_regNext_30_1_load_store_6;
  reg                 io_in_r_bypass_regNext_30_1_df_is_ws_6;
  reg                 io_in_r_bypass_regNext_30_1_stall_6;
  reg        [15:0]   io_in_r_bypass_regNext_30_2_data_6;
  reg                 io_in_r_bypass_regNext_30_2_load_store_6;
  reg                 io_in_r_bypass_regNext_30_2_df_is_ws_6;
  reg                 io_in_r_bypass_regNext_30_2_stall_6;
  reg        [15:0]   io_in_r_bypass_regNext_30_3_data_6;
  reg                 io_in_r_bypass_regNext_30_3_load_store_6;
  reg                 io_in_r_bypass_regNext_30_3_df_is_ws_6;
  reg                 io_in_r_bypass_regNext_30_3_stall_6;
  reg        [15:0]   io_in_r_bypass_regNext_31_0_data_6;
  reg                 io_in_r_bypass_regNext_31_0_load_store_6;
  reg                 io_in_r_bypass_regNext_31_0_df_is_ws_6;
  reg                 io_in_r_bypass_regNext_31_0_stall_6;
  reg        [15:0]   io_in_r_bypass_regNext_31_1_data_6;
  reg                 io_in_r_bypass_regNext_31_1_load_store_6;
  reg                 io_in_r_bypass_regNext_31_1_df_is_ws_6;
  reg                 io_in_r_bypass_regNext_31_1_stall_6;
  reg        [15:0]   io_in_r_bypass_regNext_31_2_data_6;
  reg                 io_in_r_bypass_regNext_31_2_load_store_6;
  reg                 io_in_r_bypass_regNext_31_2_df_is_ws_6;
  reg                 io_in_r_bypass_regNext_31_2_stall_6;
  reg        [15:0]   io_in_r_bypass_regNext_31_3_data_6;
  reg                 io_in_r_bypass_regNext_31_3_load_store_6;
  reg                 io_in_r_bypass_regNext_31_3_df_is_ws_6;
  reg                 io_in_r_bypass_regNext_31_3_stall_6;
  reg        [15:0]   io_in_r_bypass_regNext_0_0_data_7;
  reg                 io_in_r_bypass_regNext_0_0_load_store_7;
  reg                 io_in_r_bypass_regNext_0_0_df_is_ws_7;
  reg                 io_in_r_bypass_regNext_0_0_stall_7;
  reg        [15:0]   io_in_r_bypass_regNext_0_1_data_7;
  reg                 io_in_r_bypass_regNext_0_1_load_store_7;
  reg                 io_in_r_bypass_regNext_0_1_df_is_ws_7;
  reg                 io_in_r_bypass_regNext_0_1_stall_7;
  reg        [15:0]   io_in_r_bypass_regNext_0_2_data_7;
  reg                 io_in_r_bypass_regNext_0_2_load_store_7;
  reg                 io_in_r_bypass_regNext_0_2_df_is_ws_7;
  reg                 io_in_r_bypass_regNext_0_2_stall_7;
  reg        [15:0]   io_in_r_bypass_regNext_0_3_data_7;
  reg                 io_in_r_bypass_regNext_0_3_load_store_7;
  reg                 io_in_r_bypass_regNext_0_3_df_is_ws_7;
  reg                 io_in_r_bypass_regNext_0_3_stall_7;
  reg        [15:0]   io_in_r_bypass_regNext_1_0_data_7;
  reg                 io_in_r_bypass_regNext_1_0_load_store_7;
  reg                 io_in_r_bypass_regNext_1_0_df_is_ws_7;
  reg                 io_in_r_bypass_regNext_1_0_stall_7;
  reg        [15:0]   io_in_r_bypass_regNext_1_1_data_7;
  reg                 io_in_r_bypass_regNext_1_1_load_store_7;
  reg                 io_in_r_bypass_regNext_1_1_df_is_ws_7;
  reg                 io_in_r_bypass_regNext_1_1_stall_7;
  reg        [15:0]   io_in_r_bypass_regNext_1_2_data_7;
  reg                 io_in_r_bypass_regNext_1_2_load_store_7;
  reg                 io_in_r_bypass_regNext_1_2_df_is_ws_7;
  reg                 io_in_r_bypass_regNext_1_2_stall_7;
  reg        [15:0]   io_in_r_bypass_regNext_1_3_data_7;
  reg                 io_in_r_bypass_regNext_1_3_load_store_7;
  reg                 io_in_r_bypass_regNext_1_3_df_is_ws_7;
  reg                 io_in_r_bypass_regNext_1_3_stall_7;
  reg        [15:0]   io_in_r_bypass_regNext_2_0_data_7;
  reg                 io_in_r_bypass_regNext_2_0_load_store_7;
  reg                 io_in_r_bypass_regNext_2_0_df_is_ws_7;
  reg                 io_in_r_bypass_regNext_2_0_stall_7;
  reg        [15:0]   io_in_r_bypass_regNext_2_1_data_7;
  reg                 io_in_r_bypass_regNext_2_1_load_store_7;
  reg                 io_in_r_bypass_regNext_2_1_df_is_ws_7;
  reg                 io_in_r_bypass_regNext_2_1_stall_7;
  reg        [15:0]   io_in_r_bypass_regNext_2_2_data_7;
  reg                 io_in_r_bypass_regNext_2_2_load_store_7;
  reg                 io_in_r_bypass_regNext_2_2_df_is_ws_7;
  reg                 io_in_r_bypass_regNext_2_2_stall_7;
  reg        [15:0]   io_in_r_bypass_regNext_2_3_data_7;
  reg                 io_in_r_bypass_regNext_2_3_load_store_7;
  reg                 io_in_r_bypass_regNext_2_3_df_is_ws_7;
  reg                 io_in_r_bypass_regNext_2_3_stall_7;
  reg        [15:0]   io_in_r_bypass_regNext_3_0_data_7;
  reg                 io_in_r_bypass_regNext_3_0_load_store_7;
  reg                 io_in_r_bypass_regNext_3_0_df_is_ws_7;
  reg                 io_in_r_bypass_regNext_3_0_stall_7;
  reg        [15:0]   io_in_r_bypass_regNext_3_1_data_7;
  reg                 io_in_r_bypass_regNext_3_1_load_store_7;
  reg                 io_in_r_bypass_regNext_3_1_df_is_ws_7;
  reg                 io_in_r_bypass_regNext_3_1_stall_7;
  reg        [15:0]   io_in_r_bypass_regNext_3_2_data_7;
  reg                 io_in_r_bypass_regNext_3_2_load_store_7;
  reg                 io_in_r_bypass_regNext_3_2_df_is_ws_7;
  reg                 io_in_r_bypass_regNext_3_2_stall_7;
  reg        [15:0]   io_in_r_bypass_regNext_3_3_data_7;
  reg                 io_in_r_bypass_regNext_3_3_load_store_7;
  reg                 io_in_r_bypass_regNext_3_3_df_is_ws_7;
  reg                 io_in_r_bypass_regNext_3_3_stall_7;
  reg        [15:0]   io_in_r_bypass_regNext_4_0_data_7;
  reg                 io_in_r_bypass_regNext_4_0_load_store_7;
  reg                 io_in_r_bypass_regNext_4_0_df_is_ws_7;
  reg                 io_in_r_bypass_regNext_4_0_stall_7;
  reg        [15:0]   io_in_r_bypass_regNext_4_1_data_7;
  reg                 io_in_r_bypass_regNext_4_1_load_store_7;
  reg                 io_in_r_bypass_regNext_4_1_df_is_ws_7;
  reg                 io_in_r_bypass_regNext_4_1_stall_7;
  reg        [15:0]   io_in_r_bypass_regNext_4_2_data_7;
  reg                 io_in_r_bypass_regNext_4_2_load_store_7;
  reg                 io_in_r_bypass_regNext_4_2_df_is_ws_7;
  reg                 io_in_r_bypass_regNext_4_2_stall_7;
  reg        [15:0]   io_in_r_bypass_regNext_4_3_data_7;
  reg                 io_in_r_bypass_regNext_4_3_load_store_7;
  reg                 io_in_r_bypass_regNext_4_3_df_is_ws_7;
  reg                 io_in_r_bypass_regNext_4_3_stall_7;
  reg        [15:0]   io_in_r_bypass_regNext_5_0_data_7;
  reg                 io_in_r_bypass_regNext_5_0_load_store_7;
  reg                 io_in_r_bypass_regNext_5_0_df_is_ws_7;
  reg                 io_in_r_bypass_regNext_5_0_stall_7;
  reg        [15:0]   io_in_r_bypass_regNext_5_1_data_7;
  reg                 io_in_r_bypass_regNext_5_1_load_store_7;
  reg                 io_in_r_bypass_regNext_5_1_df_is_ws_7;
  reg                 io_in_r_bypass_regNext_5_1_stall_7;
  reg        [15:0]   io_in_r_bypass_regNext_5_2_data_7;
  reg                 io_in_r_bypass_regNext_5_2_load_store_7;
  reg                 io_in_r_bypass_regNext_5_2_df_is_ws_7;
  reg                 io_in_r_bypass_regNext_5_2_stall_7;
  reg        [15:0]   io_in_r_bypass_regNext_5_3_data_7;
  reg                 io_in_r_bypass_regNext_5_3_load_store_7;
  reg                 io_in_r_bypass_regNext_5_3_df_is_ws_7;
  reg                 io_in_r_bypass_regNext_5_3_stall_7;
  reg        [15:0]   io_in_r_bypass_regNext_6_0_data_7;
  reg                 io_in_r_bypass_regNext_6_0_load_store_7;
  reg                 io_in_r_bypass_regNext_6_0_df_is_ws_7;
  reg                 io_in_r_bypass_regNext_6_0_stall_7;
  reg        [15:0]   io_in_r_bypass_regNext_6_1_data_7;
  reg                 io_in_r_bypass_regNext_6_1_load_store_7;
  reg                 io_in_r_bypass_regNext_6_1_df_is_ws_7;
  reg                 io_in_r_bypass_regNext_6_1_stall_7;
  reg        [15:0]   io_in_r_bypass_regNext_6_2_data_7;
  reg                 io_in_r_bypass_regNext_6_2_load_store_7;
  reg                 io_in_r_bypass_regNext_6_2_df_is_ws_7;
  reg                 io_in_r_bypass_regNext_6_2_stall_7;
  reg        [15:0]   io_in_r_bypass_regNext_6_3_data_7;
  reg                 io_in_r_bypass_regNext_6_3_load_store_7;
  reg                 io_in_r_bypass_regNext_6_3_df_is_ws_7;
  reg                 io_in_r_bypass_regNext_6_3_stall_7;
  reg        [15:0]   io_in_r_bypass_regNext_7_0_data_7;
  reg                 io_in_r_bypass_regNext_7_0_load_store_7;
  reg                 io_in_r_bypass_regNext_7_0_df_is_ws_7;
  reg                 io_in_r_bypass_regNext_7_0_stall_7;
  reg        [15:0]   io_in_r_bypass_regNext_7_1_data_7;
  reg                 io_in_r_bypass_regNext_7_1_load_store_7;
  reg                 io_in_r_bypass_regNext_7_1_df_is_ws_7;
  reg                 io_in_r_bypass_regNext_7_1_stall_7;
  reg        [15:0]   io_in_r_bypass_regNext_7_2_data_7;
  reg                 io_in_r_bypass_regNext_7_2_load_store_7;
  reg                 io_in_r_bypass_regNext_7_2_df_is_ws_7;
  reg                 io_in_r_bypass_regNext_7_2_stall_7;
  reg        [15:0]   io_in_r_bypass_regNext_7_3_data_7;
  reg                 io_in_r_bypass_regNext_7_3_load_store_7;
  reg                 io_in_r_bypass_regNext_7_3_df_is_ws_7;
  reg                 io_in_r_bypass_regNext_7_3_stall_7;
  reg        [15:0]   io_in_r_bypass_regNext_8_0_data_7;
  reg                 io_in_r_bypass_regNext_8_0_load_store_7;
  reg                 io_in_r_bypass_regNext_8_0_df_is_ws_7;
  reg                 io_in_r_bypass_regNext_8_0_stall_7;
  reg        [15:0]   io_in_r_bypass_regNext_8_1_data_7;
  reg                 io_in_r_bypass_regNext_8_1_load_store_7;
  reg                 io_in_r_bypass_regNext_8_1_df_is_ws_7;
  reg                 io_in_r_bypass_regNext_8_1_stall_7;
  reg        [15:0]   io_in_r_bypass_regNext_8_2_data_7;
  reg                 io_in_r_bypass_regNext_8_2_load_store_7;
  reg                 io_in_r_bypass_regNext_8_2_df_is_ws_7;
  reg                 io_in_r_bypass_regNext_8_2_stall_7;
  reg        [15:0]   io_in_r_bypass_regNext_8_3_data_7;
  reg                 io_in_r_bypass_regNext_8_3_load_store_7;
  reg                 io_in_r_bypass_regNext_8_3_df_is_ws_7;
  reg                 io_in_r_bypass_regNext_8_3_stall_7;
  reg        [15:0]   io_in_r_bypass_regNext_9_0_data_7;
  reg                 io_in_r_bypass_regNext_9_0_load_store_7;
  reg                 io_in_r_bypass_regNext_9_0_df_is_ws_7;
  reg                 io_in_r_bypass_regNext_9_0_stall_7;
  reg        [15:0]   io_in_r_bypass_regNext_9_1_data_7;
  reg                 io_in_r_bypass_regNext_9_1_load_store_7;
  reg                 io_in_r_bypass_regNext_9_1_df_is_ws_7;
  reg                 io_in_r_bypass_regNext_9_1_stall_7;
  reg        [15:0]   io_in_r_bypass_regNext_9_2_data_7;
  reg                 io_in_r_bypass_regNext_9_2_load_store_7;
  reg                 io_in_r_bypass_regNext_9_2_df_is_ws_7;
  reg                 io_in_r_bypass_regNext_9_2_stall_7;
  reg        [15:0]   io_in_r_bypass_regNext_9_3_data_7;
  reg                 io_in_r_bypass_regNext_9_3_load_store_7;
  reg                 io_in_r_bypass_regNext_9_3_df_is_ws_7;
  reg                 io_in_r_bypass_regNext_9_3_stall_7;
  reg        [15:0]   io_in_r_bypass_regNext_10_0_data_7;
  reg                 io_in_r_bypass_regNext_10_0_load_store_7;
  reg                 io_in_r_bypass_regNext_10_0_df_is_ws_7;
  reg                 io_in_r_bypass_regNext_10_0_stall_7;
  reg        [15:0]   io_in_r_bypass_regNext_10_1_data_7;
  reg                 io_in_r_bypass_regNext_10_1_load_store_7;
  reg                 io_in_r_bypass_regNext_10_1_df_is_ws_7;
  reg                 io_in_r_bypass_regNext_10_1_stall_7;
  reg        [15:0]   io_in_r_bypass_regNext_10_2_data_7;
  reg                 io_in_r_bypass_regNext_10_2_load_store_7;
  reg                 io_in_r_bypass_regNext_10_2_df_is_ws_7;
  reg                 io_in_r_bypass_regNext_10_2_stall_7;
  reg        [15:0]   io_in_r_bypass_regNext_10_3_data_7;
  reg                 io_in_r_bypass_regNext_10_3_load_store_7;
  reg                 io_in_r_bypass_regNext_10_3_df_is_ws_7;
  reg                 io_in_r_bypass_regNext_10_3_stall_7;
  reg        [15:0]   io_in_r_bypass_regNext_11_0_data_7;
  reg                 io_in_r_bypass_regNext_11_0_load_store_7;
  reg                 io_in_r_bypass_regNext_11_0_df_is_ws_7;
  reg                 io_in_r_bypass_regNext_11_0_stall_7;
  reg        [15:0]   io_in_r_bypass_regNext_11_1_data_7;
  reg                 io_in_r_bypass_regNext_11_1_load_store_7;
  reg                 io_in_r_bypass_regNext_11_1_df_is_ws_7;
  reg                 io_in_r_bypass_regNext_11_1_stall_7;
  reg        [15:0]   io_in_r_bypass_regNext_11_2_data_7;
  reg                 io_in_r_bypass_regNext_11_2_load_store_7;
  reg                 io_in_r_bypass_regNext_11_2_df_is_ws_7;
  reg                 io_in_r_bypass_regNext_11_2_stall_7;
  reg        [15:0]   io_in_r_bypass_regNext_11_3_data_7;
  reg                 io_in_r_bypass_regNext_11_3_load_store_7;
  reg                 io_in_r_bypass_regNext_11_3_df_is_ws_7;
  reg                 io_in_r_bypass_regNext_11_3_stall_7;
  reg        [15:0]   io_in_r_bypass_regNext_12_0_data_7;
  reg                 io_in_r_bypass_regNext_12_0_load_store_7;
  reg                 io_in_r_bypass_regNext_12_0_df_is_ws_7;
  reg                 io_in_r_bypass_regNext_12_0_stall_7;
  reg        [15:0]   io_in_r_bypass_regNext_12_1_data_7;
  reg                 io_in_r_bypass_regNext_12_1_load_store_7;
  reg                 io_in_r_bypass_regNext_12_1_df_is_ws_7;
  reg                 io_in_r_bypass_regNext_12_1_stall_7;
  reg        [15:0]   io_in_r_bypass_regNext_12_2_data_7;
  reg                 io_in_r_bypass_regNext_12_2_load_store_7;
  reg                 io_in_r_bypass_regNext_12_2_df_is_ws_7;
  reg                 io_in_r_bypass_regNext_12_2_stall_7;
  reg        [15:0]   io_in_r_bypass_regNext_12_3_data_7;
  reg                 io_in_r_bypass_regNext_12_3_load_store_7;
  reg                 io_in_r_bypass_regNext_12_3_df_is_ws_7;
  reg                 io_in_r_bypass_regNext_12_3_stall_7;
  reg        [15:0]   io_in_r_bypass_regNext_13_0_data_7;
  reg                 io_in_r_bypass_regNext_13_0_load_store_7;
  reg                 io_in_r_bypass_regNext_13_0_df_is_ws_7;
  reg                 io_in_r_bypass_regNext_13_0_stall_7;
  reg        [15:0]   io_in_r_bypass_regNext_13_1_data_7;
  reg                 io_in_r_bypass_regNext_13_1_load_store_7;
  reg                 io_in_r_bypass_regNext_13_1_df_is_ws_7;
  reg                 io_in_r_bypass_regNext_13_1_stall_7;
  reg        [15:0]   io_in_r_bypass_regNext_13_2_data_7;
  reg                 io_in_r_bypass_regNext_13_2_load_store_7;
  reg                 io_in_r_bypass_regNext_13_2_df_is_ws_7;
  reg                 io_in_r_bypass_regNext_13_2_stall_7;
  reg        [15:0]   io_in_r_bypass_regNext_13_3_data_7;
  reg                 io_in_r_bypass_regNext_13_3_load_store_7;
  reg                 io_in_r_bypass_regNext_13_3_df_is_ws_7;
  reg                 io_in_r_bypass_regNext_13_3_stall_7;
  reg        [15:0]   io_in_r_bypass_regNext_14_0_data_7;
  reg                 io_in_r_bypass_regNext_14_0_load_store_7;
  reg                 io_in_r_bypass_regNext_14_0_df_is_ws_7;
  reg                 io_in_r_bypass_regNext_14_0_stall_7;
  reg        [15:0]   io_in_r_bypass_regNext_14_1_data_7;
  reg                 io_in_r_bypass_regNext_14_1_load_store_7;
  reg                 io_in_r_bypass_regNext_14_1_df_is_ws_7;
  reg                 io_in_r_bypass_regNext_14_1_stall_7;
  reg        [15:0]   io_in_r_bypass_regNext_14_2_data_7;
  reg                 io_in_r_bypass_regNext_14_2_load_store_7;
  reg                 io_in_r_bypass_regNext_14_2_df_is_ws_7;
  reg                 io_in_r_bypass_regNext_14_2_stall_7;
  reg        [15:0]   io_in_r_bypass_regNext_14_3_data_7;
  reg                 io_in_r_bypass_regNext_14_3_load_store_7;
  reg                 io_in_r_bypass_regNext_14_3_df_is_ws_7;
  reg                 io_in_r_bypass_regNext_14_3_stall_7;
  reg        [15:0]   io_in_r_bypass_regNext_15_0_data_7;
  reg                 io_in_r_bypass_regNext_15_0_load_store_7;
  reg                 io_in_r_bypass_regNext_15_0_df_is_ws_7;
  reg                 io_in_r_bypass_regNext_15_0_stall_7;
  reg        [15:0]   io_in_r_bypass_regNext_15_1_data_7;
  reg                 io_in_r_bypass_regNext_15_1_load_store_7;
  reg                 io_in_r_bypass_regNext_15_1_df_is_ws_7;
  reg                 io_in_r_bypass_regNext_15_1_stall_7;
  reg        [15:0]   io_in_r_bypass_regNext_15_2_data_7;
  reg                 io_in_r_bypass_regNext_15_2_load_store_7;
  reg                 io_in_r_bypass_regNext_15_2_df_is_ws_7;
  reg                 io_in_r_bypass_regNext_15_2_stall_7;
  reg        [15:0]   io_in_r_bypass_regNext_15_3_data_7;
  reg                 io_in_r_bypass_regNext_15_3_load_store_7;
  reg                 io_in_r_bypass_regNext_15_3_df_is_ws_7;
  reg                 io_in_r_bypass_regNext_15_3_stall_7;
  reg        [15:0]   io_in_r_bypass_regNext_16_0_data_7;
  reg                 io_in_r_bypass_regNext_16_0_load_store_7;
  reg                 io_in_r_bypass_regNext_16_0_df_is_ws_7;
  reg                 io_in_r_bypass_regNext_16_0_stall_7;
  reg        [15:0]   io_in_r_bypass_regNext_16_1_data_7;
  reg                 io_in_r_bypass_regNext_16_1_load_store_7;
  reg                 io_in_r_bypass_regNext_16_1_df_is_ws_7;
  reg                 io_in_r_bypass_regNext_16_1_stall_7;
  reg        [15:0]   io_in_r_bypass_regNext_16_2_data_7;
  reg                 io_in_r_bypass_regNext_16_2_load_store_7;
  reg                 io_in_r_bypass_regNext_16_2_df_is_ws_7;
  reg                 io_in_r_bypass_regNext_16_2_stall_7;
  reg        [15:0]   io_in_r_bypass_regNext_16_3_data_7;
  reg                 io_in_r_bypass_regNext_16_3_load_store_7;
  reg                 io_in_r_bypass_regNext_16_3_df_is_ws_7;
  reg                 io_in_r_bypass_regNext_16_3_stall_7;
  reg        [15:0]   io_in_r_bypass_regNext_17_0_data_7;
  reg                 io_in_r_bypass_regNext_17_0_load_store_7;
  reg                 io_in_r_bypass_regNext_17_0_df_is_ws_7;
  reg                 io_in_r_bypass_regNext_17_0_stall_7;
  reg        [15:0]   io_in_r_bypass_regNext_17_1_data_7;
  reg                 io_in_r_bypass_regNext_17_1_load_store_7;
  reg                 io_in_r_bypass_regNext_17_1_df_is_ws_7;
  reg                 io_in_r_bypass_regNext_17_1_stall_7;
  reg        [15:0]   io_in_r_bypass_regNext_17_2_data_7;
  reg                 io_in_r_bypass_regNext_17_2_load_store_7;
  reg                 io_in_r_bypass_regNext_17_2_df_is_ws_7;
  reg                 io_in_r_bypass_regNext_17_2_stall_7;
  reg        [15:0]   io_in_r_bypass_regNext_17_3_data_7;
  reg                 io_in_r_bypass_regNext_17_3_load_store_7;
  reg                 io_in_r_bypass_regNext_17_3_df_is_ws_7;
  reg                 io_in_r_bypass_regNext_17_3_stall_7;
  reg        [15:0]   io_in_r_bypass_regNext_18_0_data_7;
  reg                 io_in_r_bypass_regNext_18_0_load_store_7;
  reg                 io_in_r_bypass_regNext_18_0_df_is_ws_7;
  reg                 io_in_r_bypass_regNext_18_0_stall_7;
  reg        [15:0]   io_in_r_bypass_regNext_18_1_data_7;
  reg                 io_in_r_bypass_regNext_18_1_load_store_7;
  reg                 io_in_r_bypass_regNext_18_1_df_is_ws_7;
  reg                 io_in_r_bypass_regNext_18_1_stall_7;
  reg        [15:0]   io_in_r_bypass_regNext_18_2_data_7;
  reg                 io_in_r_bypass_regNext_18_2_load_store_7;
  reg                 io_in_r_bypass_regNext_18_2_df_is_ws_7;
  reg                 io_in_r_bypass_regNext_18_2_stall_7;
  reg        [15:0]   io_in_r_bypass_regNext_18_3_data_7;
  reg                 io_in_r_bypass_regNext_18_3_load_store_7;
  reg                 io_in_r_bypass_regNext_18_3_df_is_ws_7;
  reg                 io_in_r_bypass_regNext_18_3_stall_7;
  reg        [15:0]   io_in_r_bypass_regNext_19_0_data_7;
  reg                 io_in_r_bypass_regNext_19_0_load_store_7;
  reg                 io_in_r_bypass_regNext_19_0_df_is_ws_7;
  reg                 io_in_r_bypass_regNext_19_0_stall_7;
  reg        [15:0]   io_in_r_bypass_regNext_19_1_data_7;
  reg                 io_in_r_bypass_regNext_19_1_load_store_7;
  reg                 io_in_r_bypass_regNext_19_1_df_is_ws_7;
  reg                 io_in_r_bypass_regNext_19_1_stall_7;
  reg        [15:0]   io_in_r_bypass_regNext_19_2_data_7;
  reg                 io_in_r_bypass_regNext_19_2_load_store_7;
  reg                 io_in_r_bypass_regNext_19_2_df_is_ws_7;
  reg                 io_in_r_bypass_regNext_19_2_stall_7;
  reg        [15:0]   io_in_r_bypass_regNext_19_3_data_7;
  reg                 io_in_r_bypass_regNext_19_3_load_store_7;
  reg                 io_in_r_bypass_regNext_19_3_df_is_ws_7;
  reg                 io_in_r_bypass_regNext_19_3_stall_7;
  reg        [15:0]   io_in_r_bypass_regNext_20_0_data_7;
  reg                 io_in_r_bypass_regNext_20_0_load_store_7;
  reg                 io_in_r_bypass_regNext_20_0_df_is_ws_7;
  reg                 io_in_r_bypass_regNext_20_0_stall_7;
  reg        [15:0]   io_in_r_bypass_regNext_20_1_data_7;
  reg                 io_in_r_bypass_regNext_20_1_load_store_7;
  reg                 io_in_r_bypass_regNext_20_1_df_is_ws_7;
  reg                 io_in_r_bypass_regNext_20_1_stall_7;
  reg        [15:0]   io_in_r_bypass_regNext_20_2_data_7;
  reg                 io_in_r_bypass_regNext_20_2_load_store_7;
  reg                 io_in_r_bypass_regNext_20_2_df_is_ws_7;
  reg                 io_in_r_bypass_regNext_20_2_stall_7;
  reg        [15:0]   io_in_r_bypass_regNext_20_3_data_7;
  reg                 io_in_r_bypass_regNext_20_3_load_store_7;
  reg                 io_in_r_bypass_regNext_20_3_df_is_ws_7;
  reg                 io_in_r_bypass_regNext_20_3_stall_7;
  reg        [15:0]   io_in_r_bypass_regNext_21_0_data_7;
  reg                 io_in_r_bypass_regNext_21_0_load_store_7;
  reg                 io_in_r_bypass_regNext_21_0_df_is_ws_7;
  reg                 io_in_r_bypass_regNext_21_0_stall_7;
  reg        [15:0]   io_in_r_bypass_regNext_21_1_data_7;
  reg                 io_in_r_bypass_regNext_21_1_load_store_7;
  reg                 io_in_r_bypass_regNext_21_1_df_is_ws_7;
  reg                 io_in_r_bypass_regNext_21_1_stall_7;
  reg        [15:0]   io_in_r_bypass_regNext_21_2_data_7;
  reg                 io_in_r_bypass_regNext_21_2_load_store_7;
  reg                 io_in_r_bypass_regNext_21_2_df_is_ws_7;
  reg                 io_in_r_bypass_regNext_21_2_stall_7;
  reg        [15:0]   io_in_r_bypass_regNext_21_3_data_7;
  reg                 io_in_r_bypass_regNext_21_3_load_store_7;
  reg                 io_in_r_bypass_regNext_21_3_df_is_ws_7;
  reg                 io_in_r_bypass_regNext_21_3_stall_7;
  reg        [15:0]   io_in_r_bypass_regNext_22_0_data_7;
  reg                 io_in_r_bypass_regNext_22_0_load_store_7;
  reg                 io_in_r_bypass_regNext_22_0_df_is_ws_7;
  reg                 io_in_r_bypass_regNext_22_0_stall_7;
  reg        [15:0]   io_in_r_bypass_regNext_22_1_data_7;
  reg                 io_in_r_bypass_regNext_22_1_load_store_7;
  reg                 io_in_r_bypass_regNext_22_1_df_is_ws_7;
  reg                 io_in_r_bypass_regNext_22_1_stall_7;
  reg        [15:0]   io_in_r_bypass_regNext_22_2_data_7;
  reg                 io_in_r_bypass_regNext_22_2_load_store_7;
  reg                 io_in_r_bypass_regNext_22_2_df_is_ws_7;
  reg                 io_in_r_bypass_regNext_22_2_stall_7;
  reg        [15:0]   io_in_r_bypass_regNext_22_3_data_7;
  reg                 io_in_r_bypass_regNext_22_3_load_store_7;
  reg                 io_in_r_bypass_regNext_22_3_df_is_ws_7;
  reg                 io_in_r_bypass_regNext_22_3_stall_7;
  reg        [15:0]   io_in_r_bypass_regNext_23_0_data_7;
  reg                 io_in_r_bypass_regNext_23_0_load_store_7;
  reg                 io_in_r_bypass_regNext_23_0_df_is_ws_7;
  reg                 io_in_r_bypass_regNext_23_0_stall_7;
  reg        [15:0]   io_in_r_bypass_regNext_23_1_data_7;
  reg                 io_in_r_bypass_regNext_23_1_load_store_7;
  reg                 io_in_r_bypass_regNext_23_1_df_is_ws_7;
  reg                 io_in_r_bypass_regNext_23_1_stall_7;
  reg        [15:0]   io_in_r_bypass_regNext_23_2_data_7;
  reg                 io_in_r_bypass_regNext_23_2_load_store_7;
  reg                 io_in_r_bypass_regNext_23_2_df_is_ws_7;
  reg                 io_in_r_bypass_regNext_23_2_stall_7;
  reg        [15:0]   io_in_r_bypass_regNext_23_3_data_7;
  reg                 io_in_r_bypass_regNext_23_3_load_store_7;
  reg                 io_in_r_bypass_regNext_23_3_df_is_ws_7;
  reg                 io_in_r_bypass_regNext_23_3_stall_7;
  reg        [15:0]   io_in_r_bypass_regNext_24_0_data_7;
  reg                 io_in_r_bypass_regNext_24_0_load_store_7;
  reg                 io_in_r_bypass_regNext_24_0_df_is_ws_7;
  reg                 io_in_r_bypass_regNext_24_0_stall_7;
  reg        [15:0]   io_in_r_bypass_regNext_24_1_data_7;
  reg                 io_in_r_bypass_regNext_24_1_load_store_7;
  reg                 io_in_r_bypass_regNext_24_1_df_is_ws_7;
  reg                 io_in_r_bypass_regNext_24_1_stall_7;
  reg        [15:0]   io_in_r_bypass_regNext_24_2_data_7;
  reg                 io_in_r_bypass_regNext_24_2_load_store_7;
  reg                 io_in_r_bypass_regNext_24_2_df_is_ws_7;
  reg                 io_in_r_bypass_regNext_24_2_stall_7;
  reg        [15:0]   io_in_r_bypass_regNext_24_3_data_7;
  reg                 io_in_r_bypass_regNext_24_3_load_store_7;
  reg                 io_in_r_bypass_regNext_24_3_df_is_ws_7;
  reg                 io_in_r_bypass_regNext_24_3_stall_7;
  reg        [15:0]   io_in_r_bypass_regNext_25_0_data_7;
  reg                 io_in_r_bypass_regNext_25_0_load_store_7;
  reg                 io_in_r_bypass_regNext_25_0_df_is_ws_7;
  reg                 io_in_r_bypass_regNext_25_0_stall_7;
  reg        [15:0]   io_in_r_bypass_regNext_25_1_data_7;
  reg                 io_in_r_bypass_regNext_25_1_load_store_7;
  reg                 io_in_r_bypass_regNext_25_1_df_is_ws_7;
  reg                 io_in_r_bypass_regNext_25_1_stall_7;
  reg        [15:0]   io_in_r_bypass_regNext_25_2_data_7;
  reg                 io_in_r_bypass_regNext_25_2_load_store_7;
  reg                 io_in_r_bypass_regNext_25_2_df_is_ws_7;
  reg                 io_in_r_bypass_regNext_25_2_stall_7;
  reg        [15:0]   io_in_r_bypass_regNext_25_3_data_7;
  reg                 io_in_r_bypass_regNext_25_3_load_store_7;
  reg                 io_in_r_bypass_regNext_25_3_df_is_ws_7;
  reg                 io_in_r_bypass_regNext_25_3_stall_7;
  reg        [15:0]   io_in_r_bypass_regNext_26_0_data_7;
  reg                 io_in_r_bypass_regNext_26_0_load_store_7;
  reg                 io_in_r_bypass_regNext_26_0_df_is_ws_7;
  reg                 io_in_r_bypass_regNext_26_0_stall_7;
  reg        [15:0]   io_in_r_bypass_regNext_26_1_data_7;
  reg                 io_in_r_bypass_regNext_26_1_load_store_7;
  reg                 io_in_r_bypass_regNext_26_1_df_is_ws_7;
  reg                 io_in_r_bypass_regNext_26_1_stall_7;
  reg        [15:0]   io_in_r_bypass_regNext_26_2_data_7;
  reg                 io_in_r_bypass_regNext_26_2_load_store_7;
  reg                 io_in_r_bypass_regNext_26_2_df_is_ws_7;
  reg                 io_in_r_bypass_regNext_26_2_stall_7;
  reg        [15:0]   io_in_r_bypass_regNext_26_3_data_7;
  reg                 io_in_r_bypass_regNext_26_3_load_store_7;
  reg                 io_in_r_bypass_regNext_26_3_df_is_ws_7;
  reg                 io_in_r_bypass_regNext_26_3_stall_7;
  reg        [15:0]   io_in_r_bypass_regNext_27_0_data_7;
  reg                 io_in_r_bypass_regNext_27_0_load_store_7;
  reg                 io_in_r_bypass_regNext_27_0_df_is_ws_7;
  reg                 io_in_r_bypass_regNext_27_0_stall_7;
  reg        [15:0]   io_in_r_bypass_regNext_27_1_data_7;
  reg                 io_in_r_bypass_regNext_27_1_load_store_7;
  reg                 io_in_r_bypass_regNext_27_1_df_is_ws_7;
  reg                 io_in_r_bypass_regNext_27_1_stall_7;
  reg        [15:0]   io_in_r_bypass_regNext_27_2_data_7;
  reg                 io_in_r_bypass_regNext_27_2_load_store_7;
  reg                 io_in_r_bypass_regNext_27_2_df_is_ws_7;
  reg                 io_in_r_bypass_regNext_27_2_stall_7;
  reg        [15:0]   io_in_r_bypass_regNext_27_3_data_7;
  reg                 io_in_r_bypass_regNext_27_3_load_store_7;
  reg                 io_in_r_bypass_regNext_27_3_df_is_ws_7;
  reg                 io_in_r_bypass_regNext_27_3_stall_7;
  reg        [15:0]   io_in_r_bypass_regNext_28_0_data_7;
  reg                 io_in_r_bypass_regNext_28_0_load_store_7;
  reg                 io_in_r_bypass_regNext_28_0_df_is_ws_7;
  reg                 io_in_r_bypass_regNext_28_0_stall_7;
  reg        [15:0]   io_in_r_bypass_regNext_28_1_data_7;
  reg                 io_in_r_bypass_regNext_28_1_load_store_7;
  reg                 io_in_r_bypass_regNext_28_1_df_is_ws_7;
  reg                 io_in_r_bypass_regNext_28_1_stall_7;
  reg        [15:0]   io_in_r_bypass_regNext_28_2_data_7;
  reg                 io_in_r_bypass_regNext_28_2_load_store_7;
  reg                 io_in_r_bypass_regNext_28_2_df_is_ws_7;
  reg                 io_in_r_bypass_regNext_28_2_stall_7;
  reg        [15:0]   io_in_r_bypass_regNext_28_3_data_7;
  reg                 io_in_r_bypass_regNext_28_3_load_store_7;
  reg                 io_in_r_bypass_regNext_28_3_df_is_ws_7;
  reg                 io_in_r_bypass_regNext_28_3_stall_7;
  reg        [15:0]   io_in_r_bypass_regNext_29_0_data_7;
  reg                 io_in_r_bypass_regNext_29_0_load_store_7;
  reg                 io_in_r_bypass_regNext_29_0_df_is_ws_7;
  reg                 io_in_r_bypass_regNext_29_0_stall_7;
  reg        [15:0]   io_in_r_bypass_regNext_29_1_data_7;
  reg                 io_in_r_bypass_regNext_29_1_load_store_7;
  reg                 io_in_r_bypass_regNext_29_1_df_is_ws_7;
  reg                 io_in_r_bypass_regNext_29_1_stall_7;
  reg        [15:0]   io_in_r_bypass_regNext_29_2_data_7;
  reg                 io_in_r_bypass_regNext_29_2_load_store_7;
  reg                 io_in_r_bypass_regNext_29_2_df_is_ws_7;
  reg                 io_in_r_bypass_regNext_29_2_stall_7;
  reg        [15:0]   io_in_r_bypass_regNext_29_3_data_7;
  reg                 io_in_r_bypass_regNext_29_3_load_store_7;
  reg                 io_in_r_bypass_regNext_29_3_df_is_ws_7;
  reg                 io_in_r_bypass_regNext_29_3_stall_7;
  reg        [15:0]   io_in_r_bypass_regNext_30_0_data_7;
  reg                 io_in_r_bypass_regNext_30_0_load_store_7;
  reg                 io_in_r_bypass_regNext_30_0_df_is_ws_7;
  reg                 io_in_r_bypass_regNext_30_0_stall_7;
  reg        [15:0]   io_in_r_bypass_regNext_30_1_data_7;
  reg                 io_in_r_bypass_regNext_30_1_load_store_7;
  reg                 io_in_r_bypass_regNext_30_1_df_is_ws_7;
  reg                 io_in_r_bypass_regNext_30_1_stall_7;
  reg        [15:0]   io_in_r_bypass_regNext_30_2_data_7;
  reg                 io_in_r_bypass_regNext_30_2_load_store_7;
  reg                 io_in_r_bypass_regNext_30_2_df_is_ws_7;
  reg                 io_in_r_bypass_regNext_30_2_stall_7;
  reg        [15:0]   io_in_r_bypass_regNext_30_3_data_7;
  reg                 io_in_r_bypass_regNext_30_3_load_store_7;
  reg                 io_in_r_bypass_regNext_30_3_df_is_ws_7;
  reg                 io_in_r_bypass_regNext_30_3_stall_7;
  reg        [15:0]   io_in_r_bypass_regNext_31_0_data_7;
  reg                 io_in_r_bypass_regNext_31_0_load_store_7;
  reg                 io_in_r_bypass_regNext_31_0_df_is_ws_7;
  reg                 io_in_r_bypass_regNext_31_0_stall_7;
  reg        [15:0]   io_in_r_bypass_regNext_31_1_data_7;
  reg                 io_in_r_bypass_regNext_31_1_load_store_7;
  reg                 io_in_r_bypass_regNext_31_1_df_is_ws_7;
  reg                 io_in_r_bypass_regNext_31_1_stall_7;
  reg        [15:0]   io_in_r_bypass_regNext_31_2_data_7;
  reg                 io_in_r_bypass_regNext_31_2_load_store_7;
  reg                 io_in_r_bypass_regNext_31_2_df_is_ws_7;
  reg                 io_in_r_bypass_regNext_31_2_stall_7;
  reg        [15:0]   io_in_r_bypass_regNext_31_3_data_7;
  reg                 io_in_r_bypass_regNext_31_3_load_store_7;
  reg                 io_in_r_bypass_regNext_31_3_df_is_ws_7;
  reg                 io_in_r_bypass_regNext_31_3_stall_7;
  reg        [15:0]   io_in_r_bypass_regNext_0_0_data_8;
  reg                 io_in_r_bypass_regNext_0_0_load_store_8;
  reg                 io_in_r_bypass_regNext_0_0_df_is_ws_8;
  reg                 io_in_r_bypass_regNext_0_0_stall_8;
  reg        [15:0]   io_in_r_bypass_regNext_0_1_data_8;
  reg                 io_in_r_bypass_regNext_0_1_load_store_8;
  reg                 io_in_r_bypass_regNext_0_1_df_is_ws_8;
  reg                 io_in_r_bypass_regNext_0_1_stall_8;
  reg        [15:0]   io_in_r_bypass_regNext_0_2_data_8;
  reg                 io_in_r_bypass_regNext_0_2_load_store_8;
  reg                 io_in_r_bypass_regNext_0_2_df_is_ws_8;
  reg                 io_in_r_bypass_regNext_0_2_stall_8;
  reg        [15:0]   io_in_r_bypass_regNext_0_3_data_8;
  reg                 io_in_r_bypass_regNext_0_3_load_store_8;
  reg                 io_in_r_bypass_regNext_0_3_df_is_ws_8;
  reg                 io_in_r_bypass_regNext_0_3_stall_8;
  reg        [15:0]   io_in_r_bypass_regNext_1_0_data_8;
  reg                 io_in_r_bypass_regNext_1_0_load_store_8;
  reg                 io_in_r_bypass_regNext_1_0_df_is_ws_8;
  reg                 io_in_r_bypass_regNext_1_0_stall_8;
  reg        [15:0]   io_in_r_bypass_regNext_1_1_data_8;
  reg                 io_in_r_bypass_regNext_1_1_load_store_8;
  reg                 io_in_r_bypass_regNext_1_1_df_is_ws_8;
  reg                 io_in_r_bypass_regNext_1_1_stall_8;
  reg        [15:0]   io_in_r_bypass_regNext_1_2_data_8;
  reg                 io_in_r_bypass_regNext_1_2_load_store_8;
  reg                 io_in_r_bypass_regNext_1_2_df_is_ws_8;
  reg                 io_in_r_bypass_regNext_1_2_stall_8;
  reg        [15:0]   io_in_r_bypass_regNext_1_3_data_8;
  reg                 io_in_r_bypass_regNext_1_3_load_store_8;
  reg                 io_in_r_bypass_regNext_1_3_df_is_ws_8;
  reg                 io_in_r_bypass_regNext_1_3_stall_8;
  reg        [15:0]   io_in_r_bypass_regNext_2_0_data_8;
  reg                 io_in_r_bypass_regNext_2_0_load_store_8;
  reg                 io_in_r_bypass_regNext_2_0_df_is_ws_8;
  reg                 io_in_r_bypass_regNext_2_0_stall_8;
  reg        [15:0]   io_in_r_bypass_regNext_2_1_data_8;
  reg                 io_in_r_bypass_regNext_2_1_load_store_8;
  reg                 io_in_r_bypass_regNext_2_1_df_is_ws_8;
  reg                 io_in_r_bypass_regNext_2_1_stall_8;
  reg        [15:0]   io_in_r_bypass_regNext_2_2_data_8;
  reg                 io_in_r_bypass_regNext_2_2_load_store_8;
  reg                 io_in_r_bypass_regNext_2_2_df_is_ws_8;
  reg                 io_in_r_bypass_regNext_2_2_stall_8;
  reg        [15:0]   io_in_r_bypass_regNext_2_3_data_8;
  reg                 io_in_r_bypass_regNext_2_3_load_store_8;
  reg                 io_in_r_bypass_regNext_2_3_df_is_ws_8;
  reg                 io_in_r_bypass_regNext_2_3_stall_8;
  reg        [15:0]   io_in_r_bypass_regNext_3_0_data_8;
  reg                 io_in_r_bypass_regNext_3_0_load_store_8;
  reg                 io_in_r_bypass_regNext_3_0_df_is_ws_8;
  reg                 io_in_r_bypass_regNext_3_0_stall_8;
  reg        [15:0]   io_in_r_bypass_regNext_3_1_data_8;
  reg                 io_in_r_bypass_regNext_3_1_load_store_8;
  reg                 io_in_r_bypass_regNext_3_1_df_is_ws_8;
  reg                 io_in_r_bypass_regNext_3_1_stall_8;
  reg        [15:0]   io_in_r_bypass_regNext_3_2_data_8;
  reg                 io_in_r_bypass_regNext_3_2_load_store_8;
  reg                 io_in_r_bypass_regNext_3_2_df_is_ws_8;
  reg                 io_in_r_bypass_regNext_3_2_stall_8;
  reg        [15:0]   io_in_r_bypass_regNext_3_3_data_8;
  reg                 io_in_r_bypass_regNext_3_3_load_store_8;
  reg                 io_in_r_bypass_regNext_3_3_df_is_ws_8;
  reg                 io_in_r_bypass_regNext_3_3_stall_8;
  reg        [15:0]   io_in_r_bypass_regNext_4_0_data_8;
  reg                 io_in_r_bypass_regNext_4_0_load_store_8;
  reg                 io_in_r_bypass_regNext_4_0_df_is_ws_8;
  reg                 io_in_r_bypass_regNext_4_0_stall_8;
  reg        [15:0]   io_in_r_bypass_regNext_4_1_data_8;
  reg                 io_in_r_bypass_regNext_4_1_load_store_8;
  reg                 io_in_r_bypass_regNext_4_1_df_is_ws_8;
  reg                 io_in_r_bypass_regNext_4_1_stall_8;
  reg        [15:0]   io_in_r_bypass_regNext_4_2_data_8;
  reg                 io_in_r_bypass_regNext_4_2_load_store_8;
  reg                 io_in_r_bypass_regNext_4_2_df_is_ws_8;
  reg                 io_in_r_bypass_regNext_4_2_stall_8;
  reg        [15:0]   io_in_r_bypass_regNext_4_3_data_8;
  reg                 io_in_r_bypass_regNext_4_3_load_store_8;
  reg                 io_in_r_bypass_regNext_4_3_df_is_ws_8;
  reg                 io_in_r_bypass_regNext_4_3_stall_8;
  reg        [15:0]   io_in_r_bypass_regNext_5_0_data_8;
  reg                 io_in_r_bypass_regNext_5_0_load_store_8;
  reg                 io_in_r_bypass_regNext_5_0_df_is_ws_8;
  reg                 io_in_r_bypass_regNext_5_0_stall_8;
  reg        [15:0]   io_in_r_bypass_regNext_5_1_data_8;
  reg                 io_in_r_bypass_regNext_5_1_load_store_8;
  reg                 io_in_r_bypass_regNext_5_1_df_is_ws_8;
  reg                 io_in_r_bypass_regNext_5_1_stall_8;
  reg        [15:0]   io_in_r_bypass_regNext_5_2_data_8;
  reg                 io_in_r_bypass_regNext_5_2_load_store_8;
  reg                 io_in_r_bypass_regNext_5_2_df_is_ws_8;
  reg                 io_in_r_bypass_regNext_5_2_stall_8;
  reg        [15:0]   io_in_r_bypass_regNext_5_3_data_8;
  reg                 io_in_r_bypass_regNext_5_3_load_store_8;
  reg                 io_in_r_bypass_regNext_5_3_df_is_ws_8;
  reg                 io_in_r_bypass_regNext_5_3_stall_8;
  reg        [15:0]   io_in_r_bypass_regNext_6_0_data_8;
  reg                 io_in_r_bypass_regNext_6_0_load_store_8;
  reg                 io_in_r_bypass_regNext_6_0_df_is_ws_8;
  reg                 io_in_r_bypass_regNext_6_0_stall_8;
  reg        [15:0]   io_in_r_bypass_regNext_6_1_data_8;
  reg                 io_in_r_bypass_regNext_6_1_load_store_8;
  reg                 io_in_r_bypass_regNext_6_1_df_is_ws_8;
  reg                 io_in_r_bypass_regNext_6_1_stall_8;
  reg        [15:0]   io_in_r_bypass_regNext_6_2_data_8;
  reg                 io_in_r_bypass_regNext_6_2_load_store_8;
  reg                 io_in_r_bypass_regNext_6_2_df_is_ws_8;
  reg                 io_in_r_bypass_regNext_6_2_stall_8;
  reg        [15:0]   io_in_r_bypass_regNext_6_3_data_8;
  reg                 io_in_r_bypass_regNext_6_3_load_store_8;
  reg                 io_in_r_bypass_regNext_6_3_df_is_ws_8;
  reg                 io_in_r_bypass_regNext_6_3_stall_8;
  reg        [15:0]   io_in_r_bypass_regNext_7_0_data_8;
  reg                 io_in_r_bypass_regNext_7_0_load_store_8;
  reg                 io_in_r_bypass_regNext_7_0_df_is_ws_8;
  reg                 io_in_r_bypass_regNext_7_0_stall_8;
  reg        [15:0]   io_in_r_bypass_regNext_7_1_data_8;
  reg                 io_in_r_bypass_regNext_7_1_load_store_8;
  reg                 io_in_r_bypass_regNext_7_1_df_is_ws_8;
  reg                 io_in_r_bypass_regNext_7_1_stall_8;
  reg        [15:0]   io_in_r_bypass_regNext_7_2_data_8;
  reg                 io_in_r_bypass_regNext_7_2_load_store_8;
  reg                 io_in_r_bypass_regNext_7_2_df_is_ws_8;
  reg                 io_in_r_bypass_regNext_7_2_stall_8;
  reg        [15:0]   io_in_r_bypass_regNext_7_3_data_8;
  reg                 io_in_r_bypass_regNext_7_3_load_store_8;
  reg                 io_in_r_bypass_regNext_7_3_df_is_ws_8;
  reg                 io_in_r_bypass_regNext_7_3_stall_8;
  reg        [15:0]   io_in_r_bypass_regNext_8_0_data_8;
  reg                 io_in_r_bypass_regNext_8_0_load_store_8;
  reg                 io_in_r_bypass_regNext_8_0_df_is_ws_8;
  reg                 io_in_r_bypass_regNext_8_0_stall_8;
  reg        [15:0]   io_in_r_bypass_regNext_8_1_data_8;
  reg                 io_in_r_bypass_regNext_8_1_load_store_8;
  reg                 io_in_r_bypass_regNext_8_1_df_is_ws_8;
  reg                 io_in_r_bypass_regNext_8_1_stall_8;
  reg        [15:0]   io_in_r_bypass_regNext_8_2_data_8;
  reg                 io_in_r_bypass_regNext_8_2_load_store_8;
  reg                 io_in_r_bypass_regNext_8_2_df_is_ws_8;
  reg                 io_in_r_bypass_regNext_8_2_stall_8;
  reg        [15:0]   io_in_r_bypass_regNext_8_3_data_8;
  reg                 io_in_r_bypass_regNext_8_3_load_store_8;
  reg                 io_in_r_bypass_regNext_8_3_df_is_ws_8;
  reg                 io_in_r_bypass_regNext_8_3_stall_8;
  reg        [15:0]   io_in_r_bypass_regNext_9_0_data_8;
  reg                 io_in_r_bypass_regNext_9_0_load_store_8;
  reg                 io_in_r_bypass_regNext_9_0_df_is_ws_8;
  reg                 io_in_r_bypass_regNext_9_0_stall_8;
  reg        [15:0]   io_in_r_bypass_regNext_9_1_data_8;
  reg                 io_in_r_bypass_regNext_9_1_load_store_8;
  reg                 io_in_r_bypass_regNext_9_1_df_is_ws_8;
  reg                 io_in_r_bypass_regNext_9_1_stall_8;
  reg        [15:0]   io_in_r_bypass_regNext_9_2_data_8;
  reg                 io_in_r_bypass_regNext_9_2_load_store_8;
  reg                 io_in_r_bypass_regNext_9_2_df_is_ws_8;
  reg                 io_in_r_bypass_regNext_9_2_stall_8;
  reg        [15:0]   io_in_r_bypass_regNext_9_3_data_8;
  reg                 io_in_r_bypass_regNext_9_3_load_store_8;
  reg                 io_in_r_bypass_regNext_9_3_df_is_ws_8;
  reg                 io_in_r_bypass_regNext_9_3_stall_8;
  reg        [15:0]   io_in_r_bypass_regNext_10_0_data_8;
  reg                 io_in_r_bypass_regNext_10_0_load_store_8;
  reg                 io_in_r_bypass_regNext_10_0_df_is_ws_8;
  reg                 io_in_r_bypass_regNext_10_0_stall_8;
  reg        [15:0]   io_in_r_bypass_regNext_10_1_data_8;
  reg                 io_in_r_bypass_regNext_10_1_load_store_8;
  reg                 io_in_r_bypass_regNext_10_1_df_is_ws_8;
  reg                 io_in_r_bypass_regNext_10_1_stall_8;
  reg        [15:0]   io_in_r_bypass_regNext_10_2_data_8;
  reg                 io_in_r_bypass_regNext_10_2_load_store_8;
  reg                 io_in_r_bypass_regNext_10_2_df_is_ws_8;
  reg                 io_in_r_bypass_regNext_10_2_stall_8;
  reg        [15:0]   io_in_r_bypass_regNext_10_3_data_8;
  reg                 io_in_r_bypass_regNext_10_3_load_store_8;
  reg                 io_in_r_bypass_regNext_10_3_df_is_ws_8;
  reg                 io_in_r_bypass_regNext_10_3_stall_8;
  reg        [15:0]   io_in_r_bypass_regNext_11_0_data_8;
  reg                 io_in_r_bypass_regNext_11_0_load_store_8;
  reg                 io_in_r_bypass_regNext_11_0_df_is_ws_8;
  reg                 io_in_r_bypass_regNext_11_0_stall_8;
  reg        [15:0]   io_in_r_bypass_regNext_11_1_data_8;
  reg                 io_in_r_bypass_regNext_11_1_load_store_8;
  reg                 io_in_r_bypass_regNext_11_1_df_is_ws_8;
  reg                 io_in_r_bypass_regNext_11_1_stall_8;
  reg        [15:0]   io_in_r_bypass_regNext_11_2_data_8;
  reg                 io_in_r_bypass_regNext_11_2_load_store_8;
  reg                 io_in_r_bypass_regNext_11_2_df_is_ws_8;
  reg                 io_in_r_bypass_regNext_11_2_stall_8;
  reg        [15:0]   io_in_r_bypass_regNext_11_3_data_8;
  reg                 io_in_r_bypass_regNext_11_3_load_store_8;
  reg                 io_in_r_bypass_regNext_11_3_df_is_ws_8;
  reg                 io_in_r_bypass_regNext_11_3_stall_8;
  reg        [15:0]   io_in_r_bypass_regNext_12_0_data_8;
  reg                 io_in_r_bypass_regNext_12_0_load_store_8;
  reg                 io_in_r_bypass_regNext_12_0_df_is_ws_8;
  reg                 io_in_r_bypass_regNext_12_0_stall_8;
  reg        [15:0]   io_in_r_bypass_regNext_12_1_data_8;
  reg                 io_in_r_bypass_regNext_12_1_load_store_8;
  reg                 io_in_r_bypass_regNext_12_1_df_is_ws_8;
  reg                 io_in_r_bypass_regNext_12_1_stall_8;
  reg        [15:0]   io_in_r_bypass_regNext_12_2_data_8;
  reg                 io_in_r_bypass_regNext_12_2_load_store_8;
  reg                 io_in_r_bypass_regNext_12_2_df_is_ws_8;
  reg                 io_in_r_bypass_regNext_12_2_stall_8;
  reg        [15:0]   io_in_r_bypass_regNext_12_3_data_8;
  reg                 io_in_r_bypass_regNext_12_3_load_store_8;
  reg                 io_in_r_bypass_regNext_12_3_df_is_ws_8;
  reg                 io_in_r_bypass_regNext_12_3_stall_8;
  reg        [15:0]   io_in_r_bypass_regNext_13_0_data_8;
  reg                 io_in_r_bypass_regNext_13_0_load_store_8;
  reg                 io_in_r_bypass_regNext_13_0_df_is_ws_8;
  reg                 io_in_r_bypass_regNext_13_0_stall_8;
  reg        [15:0]   io_in_r_bypass_regNext_13_1_data_8;
  reg                 io_in_r_bypass_regNext_13_1_load_store_8;
  reg                 io_in_r_bypass_regNext_13_1_df_is_ws_8;
  reg                 io_in_r_bypass_regNext_13_1_stall_8;
  reg        [15:0]   io_in_r_bypass_regNext_13_2_data_8;
  reg                 io_in_r_bypass_regNext_13_2_load_store_8;
  reg                 io_in_r_bypass_regNext_13_2_df_is_ws_8;
  reg                 io_in_r_bypass_regNext_13_2_stall_8;
  reg        [15:0]   io_in_r_bypass_regNext_13_3_data_8;
  reg                 io_in_r_bypass_regNext_13_3_load_store_8;
  reg                 io_in_r_bypass_regNext_13_3_df_is_ws_8;
  reg                 io_in_r_bypass_regNext_13_3_stall_8;
  reg        [15:0]   io_in_r_bypass_regNext_14_0_data_8;
  reg                 io_in_r_bypass_regNext_14_0_load_store_8;
  reg                 io_in_r_bypass_regNext_14_0_df_is_ws_8;
  reg                 io_in_r_bypass_regNext_14_0_stall_8;
  reg        [15:0]   io_in_r_bypass_regNext_14_1_data_8;
  reg                 io_in_r_bypass_regNext_14_1_load_store_8;
  reg                 io_in_r_bypass_regNext_14_1_df_is_ws_8;
  reg                 io_in_r_bypass_regNext_14_1_stall_8;
  reg        [15:0]   io_in_r_bypass_regNext_14_2_data_8;
  reg                 io_in_r_bypass_regNext_14_2_load_store_8;
  reg                 io_in_r_bypass_regNext_14_2_df_is_ws_8;
  reg                 io_in_r_bypass_regNext_14_2_stall_8;
  reg        [15:0]   io_in_r_bypass_regNext_14_3_data_8;
  reg                 io_in_r_bypass_regNext_14_3_load_store_8;
  reg                 io_in_r_bypass_regNext_14_3_df_is_ws_8;
  reg                 io_in_r_bypass_regNext_14_3_stall_8;
  reg        [15:0]   io_in_r_bypass_regNext_15_0_data_8;
  reg                 io_in_r_bypass_regNext_15_0_load_store_8;
  reg                 io_in_r_bypass_regNext_15_0_df_is_ws_8;
  reg                 io_in_r_bypass_regNext_15_0_stall_8;
  reg        [15:0]   io_in_r_bypass_regNext_15_1_data_8;
  reg                 io_in_r_bypass_regNext_15_1_load_store_8;
  reg                 io_in_r_bypass_regNext_15_1_df_is_ws_8;
  reg                 io_in_r_bypass_regNext_15_1_stall_8;
  reg        [15:0]   io_in_r_bypass_regNext_15_2_data_8;
  reg                 io_in_r_bypass_regNext_15_2_load_store_8;
  reg                 io_in_r_bypass_regNext_15_2_df_is_ws_8;
  reg                 io_in_r_bypass_regNext_15_2_stall_8;
  reg        [15:0]   io_in_r_bypass_regNext_15_3_data_8;
  reg                 io_in_r_bypass_regNext_15_3_load_store_8;
  reg                 io_in_r_bypass_regNext_15_3_df_is_ws_8;
  reg                 io_in_r_bypass_regNext_15_3_stall_8;
  reg        [15:0]   io_in_r_bypass_regNext_16_0_data_8;
  reg                 io_in_r_bypass_regNext_16_0_load_store_8;
  reg                 io_in_r_bypass_regNext_16_0_df_is_ws_8;
  reg                 io_in_r_bypass_regNext_16_0_stall_8;
  reg        [15:0]   io_in_r_bypass_regNext_16_1_data_8;
  reg                 io_in_r_bypass_regNext_16_1_load_store_8;
  reg                 io_in_r_bypass_regNext_16_1_df_is_ws_8;
  reg                 io_in_r_bypass_regNext_16_1_stall_8;
  reg        [15:0]   io_in_r_bypass_regNext_16_2_data_8;
  reg                 io_in_r_bypass_regNext_16_2_load_store_8;
  reg                 io_in_r_bypass_regNext_16_2_df_is_ws_8;
  reg                 io_in_r_bypass_regNext_16_2_stall_8;
  reg        [15:0]   io_in_r_bypass_regNext_16_3_data_8;
  reg                 io_in_r_bypass_regNext_16_3_load_store_8;
  reg                 io_in_r_bypass_regNext_16_3_df_is_ws_8;
  reg                 io_in_r_bypass_regNext_16_3_stall_8;
  reg        [15:0]   io_in_r_bypass_regNext_17_0_data_8;
  reg                 io_in_r_bypass_regNext_17_0_load_store_8;
  reg                 io_in_r_bypass_regNext_17_0_df_is_ws_8;
  reg                 io_in_r_bypass_regNext_17_0_stall_8;
  reg        [15:0]   io_in_r_bypass_regNext_17_1_data_8;
  reg                 io_in_r_bypass_regNext_17_1_load_store_8;
  reg                 io_in_r_bypass_regNext_17_1_df_is_ws_8;
  reg                 io_in_r_bypass_regNext_17_1_stall_8;
  reg        [15:0]   io_in_r_bypass_regNext_17_2_data_8;
  reg                 io_in_r_bypass_regNext_17_2_load_store_8;
  reg                 io_in_r_bypass_regNext_17_2_df_is_ws_8;
  reg                 io_in_r_bypass_regNext_17_2_stall_8;
  reg        [15:0]   io_in_r_bypass_regNext_17_3_data_8;
  reg                 io_in_r_bypass_regNext_17_3_load_store_8;
  reg                 io_in_r_bypass_regNext_17_3_df_is_ws_8;
  reg                 io_in_r_bypass_regNext_17_3_stall_8;
  reg        [15:0]   io_in_r_bypass_regNext_18_0_data_8;
  reg                 io_in_r_bypass_regNext_18_0_load_store_8;
  reg                 io_in_r_bypass_regNext_18_0_df_is_ws_8;
  reg                 io_in_r_bypass_regNext_18_0_stall_8;
  reg        [15:0]   io_in_r_bypass_regNext_18_1_data_8;
  reg                 io_in_r_bypass_regNext_18_1_load_store_8;
  reg                 io_in_r_bypass_regNext_18_1_df_is_ws_8;
  reg                 io_in_r_bypass_regNext_18_1_stall_8;
  reg        [15:0]   io_in_r_bypass_regNext_18_2_data_8;
  reg                 io_in_r_bypass_regNext_18_2_load_store_8;
  reg                 io_in_r_bypass_regNext_18_2_df_is_ws_8;
  reg                 io_in_r_bypass_regNext_18_2_stall_8;
  reg        [15:0]   io_in_r_bypass_regNext_18_3_data_8;
  reg                 io_in_r_bypass_regNext_18_3_load_store_8;
  reg                 io_in_r_bypass_regNext_18_3_df_is_ws_8;
  reg                 io_in_r_bypass_regNext_18_3_stall_8;
  reg        [15:0]   io_in_r_bypass_regNext_19_0_data_8;
  reg                 io_in_r_bypass_regNext_19_0_load_store_8;
  reg                 io_in_r_bypass_regNext_19_0_df_is_ws_8;
  reg                 io_in_r_bypass_regNext_19_0_stall_8;
  reg        [15:0]   io_in_r_bypass_regNext_19_1_data_8;
  reg                 io_in_r_bypass_regNext_19_1_load_store_8;
  reg                 io_in_r_bypass_regNext_19_1_df_is_ws_8;
  reg                 io_in_r_bypass_regNext_19_1_stall_8;
  reg        [15:0]   io_in_r_bypass_regNext_19_2_data_8;
  reg                 io_in_r_bypass_regNext_19_2_load_store_8;
  reg                 io_in_r_bypass_regNext_19_2_df_is_ws_8;
  reg                 io_in_r_bypass_regNext_19_2_stall_8;
  reg        [15:0]   io_in_r_bypass_regNext_19_3_data_8;
  reg                 io_in_r_bypass_regNext_19_3_load_store_8;
  reg                 io_in_r_bypass_regNext_19_3_df_is_ws_8;
  reg                 io_in_r_bypass_regNext_19_3_stall_8;
  reg        [15:0]   io_in_r_bypass_regNext_20_0_data_8;
  reg                 io_in_r_bypass_regNext_20_0_load_store_8;
  reg                 io_in_r_bypass_regNext_20_0_df_is_ws_8;
  reg                 io_in_r_bypass_regNext_20_0_stall_8;
  reg        [15:0]   io_in_r_bypass_regNext_20_1_data_8;
  reg                 io_in_r_bypass_regNext_20_1_load_store_8;
  reg                 io_in_r_bypass_regNext_20_1_df_is_ws_8;
  reg                 io_in_r_bypass_regNext_20_1_stall_8;
  reg        [15:0]   io_in_r_bypass_regNext_20_2_data_8;
  reg                 io_in_r_bypass_regNext_20_2_load_store_8;
  reg                 io_in_r_bypass_regNext_20_2_df_is_ws_8;
  reg                 io_in_r_bypass_regNext_20_2_stall_8;
  reg        [15:0]   io_in_r_bypass_regNext_20_3_data_8;
  reg                 io_in_r_bypass_regNext_20_3_load_store_8;
  reg                 io_in_r_bypass_regNext_20_3_df_is_ws_8;
  reg                 io_in_r_bypass_regNext_20_3_stall_8;
  reg        [15:0]   io_in_r_bypass_regNext_21_0_data_8;
  reg                 io_in_r_bypass_regNext_21_0_load_store_8;
  reg                 io_in_r_bypass_regNext_21_0_df_is_ws_8;
  reg                 io_in_r_bypass_regNext_21_0_stall_8;
  reg        [15:0]   io_in_r_bypass_regNext_21_1_data_8;
  reg                 io_in_r_bypass_regNext_21_1_load_store_8;
  reg                 io_in_r_bypass_regNext_21_1_df_is_ws_8;
  reg                 io_in_r_bypass_regNext_21_1_stall_8;
  reg        [15:0]   io_in_r_bypass_regNext_21_2_data_8;
  reg                 io_in_r_bypass_regNext_21_2_load_store_8;
  reg                 io_in_r_bypass_regNext_21_2_df_is_ws_8;
  reg                 io_in_r_bypass_regNext_21_2_stall_8;
  reg        [15:0]   io_in_r_bypass_regNext_21_3_data_8;
  reg                 io_in_r_bypass_regNext_21_3_load_store_8;
  reg                 io_in_r_bypass_regNext_21_3_df_is_ws_8;
  reg                 io_in_r_bypass_regNext_21_3_stall_8;
  reg        [15:0]   io_in_r_bypass_regNext_22_0_data_8;
  reg                 io_in_r_bypass_regNext_22_0_load_store_8;
  reg                 io_in_r_bypass_regNext_22_0_df_is_ws_8;
  reg                 io_in_r_bypass_regNext_22_0_stall_8;
  reg        [15:0]   io_in_r_bypass_regNext_22_1_data_8;
  reg                 io_in_r_bypass_regNext_22_1_load_store_8;
  reg                 io_in_r_bypass_regNext_22_1_df_is_ws_8;
  reg                 io_in_r_bypass_regNext_22_1_stall_8;
  reg        [15:0]   io_in_r_bypass_regNext_22_2_data_8;
  reg                 io_in_r_bypass_regNext_22_2_load_store_8;
  reg                 io_in_r_bypass_regNext_22_2_df_is_ws_8;
  reg                 io_in_r_bypass_regNext_22_2_stall_8;
  reg        [15:0]   io_in_r_bypass_regNext_22_3_data_8;
  reg                 io_in_r_bypass_regNext_22_3_load_store_8;
  reg                 io_in_r_bypass_regNext_22_3_df_is_ws_8;
  reg                 io_in_r_bypass_regNext_22_3_stall_8;
  reg        [15:0]   io_in_r_bypass_regNext_23_0_data_8;
  reg                 io_in_r_bypass_regNext_23_0_load_store_8;
  reg                 io_in_r_bypass_regNext_23_0_df_is_ws_8;
  reg                 io_in_r_bypass_regNext_23_0_stall_8;
  reg        [15:0]   io_in_r_bypass_regNext_23_1_data_8;
  reg                 io_in_r_bypass_regNext_23_1_load_store_8;
  reg                 io_in_r_bypass_regNext_23_1_df_is_ws_8;
  reg                 io_in_r_bypass_regNext_23_1_stall_8;
  reg        [15:0]   io_in_r_bypass_regNext_23_2_data_8;
  reg                 io_in_r_bypass_regNext_23_2_load_store_8;
  reg                 io_in_r_bypass_regNext_23_2_df_is_ws_8;
  reg                 io_in_r_bypass_regNext_23_2_stall_8;
  reg        [15:0]   io_in_r_bypass_regNext_23_3_data_8;
  reg                 io_in_r_bypass_regNext_23_3_load_store_8;
  reg                 io_in_r_bypass_regNext_23_3_df_is_ws_8;
  reg                 io_in_r_bypass_regNext_23_3_stall_8;
  reg        [15:0]   io_in_r_bypass_regNext_24_0_data_8;
  reg                 io_in_r_bypass_regNext_24_0_load_store_8;
  reg                 io_in_r_bypass_regNext_24_0_df_is_ws_8;
  reg                 io_in_r_bypass_regNext_24_0_stall_8;
  reg        [15:0]   io_in_r_bypass_regNext_24_1_data_8;
  reg                 io_in_r_bypass_regNext_24_1_load_store_8;
  reg                 io_in_r_bypass_regNext_24_1_df_is_ws_8;
  reg                 io_in_r_bypass_regNext_24_1_stall_8;
  reg        [15:0]   io_in_r_bypass_regNext_24_2_data_8;
  reg                 io_in_r_bypass_regNext_24_2_load_store_8;
  reg                 io_in_r_bypass_regNext_24_2_df_is_ws_8;
  reg                 io_in_r_bypass_regNext_24_2_stall_8;
  reg        [15:0]   io_in_r_bypass_regNext_24_3_data_8;
  reg                 io_in_r_bypass_regNext_24_3_load_store_8;
  reg                 io_in_r_bypass_regNext_24_3_df_is_ws_8;
  reg                 io_in_r_bypass_regNext_24_3_stall_8;
  reg        [15:0]   io_in_r_bypass_regNext_25_0_data_8;
  reg                 io_in_r_bypass_regNext_25_0_load_store_8;
  reg                 io_in_r_bypass_regNext_25_0_df_is_ws_8;
  reg                 io_in_r_bypass_regNext_25_0_stall_8;
  reg        [15:0]   io_in_r_bypass_regNext_25_1_data_8;
  reg                 io_in_r_bypass_regNext_25_1_load_store_8;
  reg                 io_in_r_bypass_regNext_25_1_df_is_ws_8;
  reg                 io_in_r_bypass_regNext_25_1_stall_8;
  reg        [15:0]   io_in_r_bypass_regNext_25_2_data_8;
  reg                 io_in_r_bypass_regNext_25_2_load_store_8;
  reg                 io_in_r_bypass_regNext_25_2_df_is_ws_8;
  reg                 io_in_r_bypass_regNext_25_2_stall_8;
  reg        [15:0]   io_in_r_bypass_regNext_25_3_data_8;
  reg                 io_in_r_bypass_regNext_25_3_load_store_8;
  reg                 io_in_r_bypass_regNext_25_3_df_is_ws_8;
  reg                 io_in_r_bypass_regNext_25_3_stall_8;
  reg        [15:0]   io_in_r_bypass_regNext_26_0_data_8;
  reg                 io_in_r_bypass_regNext_26_0_load_store_8;
  reg                 io_in_r_bypass_regNext_26_0_df_is_ws_8;
  reg                 io_in_r_bypass_regNext_26_0_stall_8;
  reg        [15:0]   io_in_r_bypass_regNext_26_1_data_8;
  reg                 io_in_r_bypass_regNext_26_1_load_store_8;
  reg                 io_in_r_bypass_regNext_26_1_df_is_ws_8;
  reg                 io_in_r_bypass_regNext_26_1_stall_8;
  reg        [15:0]   io_in_r_bypass_regNext_26_2_data_8;
  reg                 io_in_r_bypass_regNext_26_2_load_store_8;
  reg                 io_in_r_bypass_regNext_26_2_df_is_ws_8;
  reg                 io_in_r_bypass_regNext_26_2_stall_8;
  reg        [15:0]   io_in_r_bypass_regNext_26_3_data_8;
  reg                 io_in_r_bypass_regNext_26_3_load_store_8;
  reg                 io_in_r_bypass_regNext_26_3_df_is_ws_8;
  reg                 io_in_r_bypass_regNext_26_3_stall_8;
  reg        [15:0]   io_in_r_bypass_regNext_27_0_data_8;
  reg                 io_in_r_bypass_regNext_27_0_load_store_8;
  reg                 io_in_r_bypass_regNext_27_0_df_is_ws_8;
  reg                 io_in_r_bypass_regNext_27_0_stall_8;
  reg        [15:0]   io_in_r_bypass_regNext_27_1_data_8;
  reg                 io_in_r_bypass_regNext_27_1_load_store_8;
  reg                 io_in_r_bypass_regNext_27_1_df_is_ws_8;
  reg                 io_in_r_bypass_regNext_27_1_stall_8;
  reg        [15:0]   io_in_r_bypass_regNext_27_2_data_8;
  reg                 io_in_r_bypass_regNext_27_2_load_store_8;
  reg                 io_in_r_bypass_regNext_27_2_df_is_ws_8;
  reg                 io_in_r_bypass_regNext_27_2_stall_8;
  reg        [15:0]   io_in_r_bypass_regNext_27_3_data_8;
  reg                 io_in_r_bypass_regNext_27_3_load_store_8;
  reg                 io_in_r_bypass_regNext_27_3_df_is_ws_8;
  reg                 io_in_r_bypass_regNext_27_3_stall_8;
  reg        [15:0]   io_in_r_bypass_regNext_28_0_data_8;
  reg                 io_in_r_bypass_regNext_28_0_load_store_8;
  reg                 io_in_r_bypass_regNext_28_0_df_is_ws_8;
  reg                 io_in_r_bypass_regNext_28_0_stall_8;
  reg        [15:0]   io_in_r_bypass_regNext_28_1_data_8;
  reg                 io_in_r_bypass_regNext_28_1_load_store_8;
  reg                 io_in_r_bypass_regNext_28_1_df_is_ws_8;
  reg                 io_in_r_bypass_regNext_28_1_stall_8;
  reg        [15:0]   io_in_r_bypass_regNext_28_2_data_8;
  reg                 io_in_r_bypass_regNext_28_2_load_store_8;
  reg                 io_in_r_bypass_regNext_28_2_df_is_ws_8;
  reg                 io_in_r_bypass_regNext_28_2_stall_8;
  reg        [15:0]   io_in_r_bypass_regNext_28_3_data_8;
  reg                 io_in_r_bypass_regNext_28_3_load_store_8;
  reg                 io_in_r_bypass_regNext_28_3_df_is_ws_8;
  reg                 io_in_r_bypass_regNext_28_3_stall_8;
  reg        [15:0]   io_in_r_bypass_regNext_29_0_data_8;
  reg                 io_in_r_bypass_regNext_29_0_load_store_8;
  reg                 io_in_r_bypass_regNext_29_0_df_is_ws_8;
  reg                 io_in_r_bypass_regNext_29_0_stall_8;
  reg        [15:0]   io_in_r_bypass_regNext_29_1_data_8;
  reg                 io_in_r_bypass_regNext_29_1_load_store_8;
  reg                 io_in_r_bypass_regNext_29_1_df_is_ws_8;
  reg                 io_in_r_bypass_regNext_29_1_stall_8;
  reg        [15:0]   io_in_r_bypass_regNext_29_2_data_8;
  reg                 io_in_r_bypass_regNext_29_2_load_store_8;
  reg                 io_in_r_bypass_regNext_29_2_df_is_ws_8;
  reg                 io_in_r_bypass_regNext_29_2_stall_8;
  reg        [15:0]   io_in_r_bypass_regNext_29_3_data_8;
  reg                 io_in_r_bypass_regNext_29_3_load_store_8;
  reg                 io_in_r_bypass_regNext_29_3_df_is_ws_8;
  reg                 io_in_r_bypass_regNext_29_3_stall_8;
  reg        [15:0]   io_in_r_bypass_regNext_30_0_data_8;
  reg                 io_in_r_bypass_regNext_30_0_load_store_8;
  reg                 io_in_r_bypass_regNext_30_0_df_is_ws_8;
  reg                 io_in_r_bypass_regNext_30_0_stall_8;
  reg        [15:0]   io_in_r_bypass_regNext_30_1_data_8;
  reg                 io_in_r_bypass_regNext_30_1_load_store_8;
  reg                 io_in_r_bypass_regNext_30_1_df_is_ws_8;
  reg                 io_in_r_bypass_regNext_30_1_stall_8;
  reg        [15:0]   io_in_r_bypass_regNext_30_2_data_8;
  reg                 io_in_r_bypass_regNext_30_2_load_store_8;
  reg                 io_in_r_bypass_regNext_30_2_df_is_ws_8;
  reg                 io_in_r_bypass_regNext_30_2_stall_8;
  reg        [15:0]   io_in_r_bypass_regNext_30_3_data_8;
  reg                 io_in_r_bypass_regNext_30_3_load_store_8;
  reg                 io_in_r_bypass_regNext_30_3_df_is_ws_8;
  reg                 io_in_r_bypass_regNext_30_3_stall_8;
  reg        [15:0]   io_in_r_bypass_regNext_31_0_data_8;
  reg                 io_in_r_bypass_regNext_31_0_load_store_8;
  reg                 io_in_r_bypass_regNext_31_0_df_is_ws_8;
  reg                 io_in_r_bypass_regNext_31_0_stall_8;
  reg        [15:0]   io_in_r_bypass_regNext_31_1_data_8;
  reg                 io_in_r_bypass_regNext_31_1_load_store_8;
  reg                 io_in_r_bypass_regNext_31_1_df_is_ws_8;
  reg                 io_in_r_bypass_regNext_31_1_stall_8;
  reg        [15:0]   io_in_r_bypass_regNext_31_2_data_8;
  reg                 io_in_r_bypass_regNext_31_2_load_store_8;
  reg                 io_in_r_bypass_regNext_31_2_df_is_ws_8;
  reg                 io_in_r_bypass_regNext_31_2_stall_8;
  reg        [15:0]   io_in_r_bypass_regNext_31_3_data_8;
  reg                 io_in_r_bypass_regNext_31_3_load_store_8;
  reg                 io_in_r_bypass_regNext_31_3_df_is_ws_8;
  reg                 io_in_r_bypass_regNext_31_3_stall_8;
  reg        [15:0]   io_in_r_bypass_regNext_0_0_data_9;
  reg                 io_in_r_bypass_regNext_0_0_load_store_9;
  reg                 io_in_r_bypass_regNext_0_0_df_is_ws_9;
  reg                 io_in_r_bypass_regNext_0_0_stall_9;
  reg        [15:0]   io_in_r_bypass_regNext_0_1_data_9;
  reg                 io_in_r_bypass_regNext_0_1_load_store_9;
  reg                 io_in_r_bypass_regNext_0_1_df_is_ws_9;
  reg                 io_in_r_bypass_regNext_0_1_stall_9;
  reg        [15:0]   io_in_r_bypass_regNext_0_2_data_9;
  reg                 io_in_r_bypass_regNext_0_2_load_store_9;
  reg                 io_in_r_bypass_regNext_0_2_df_is_ws_9;
  reg                 io_in_r_bypass_regNext_0_2_stall_9;
  reg        [15:0]   io_in_r_bypass_regNext_0_3_data_9;
  reg                 io_in_r_bypass_regNext_0_3_load_store_9;
  reg                 io_in_r_bypass_regNext_0_3_df_is_ws_9;
  reg                 io_in_r_bypass_regNext_0_3_stall_9;
  reg        [15:0]   io_in_r_bypass_regNext_1_0_data_9;
  reg                 io_in_r_bypass_regNext_1_0_load_store_9;
  reg                 io_in_r_bypass_regNext_1_0_df_is_ws_9;
  reg                 io_in_r_bypass_regNext_1_0_stall_9;
  reg        [15:0]   io_in_r_bypass_regNext_1_1_data_9;
  reg                 io_in_r_bypass_regNext_1_1_load_store_9;
  reg                 io_in_r_bypass_regNext_1_1_df_is_ws_9;
  reg                 io_in_r_bypass_regNext_1_1_stall_9;
  reg        [15:0]   io_in_r_bypass_regNext_1_2_data_9;
  reg                 io_in_r_bypass_regNext_1_2_load_store_9;
  reg                 io_in_r_bypass_regNext_1_2_df_is_ws_9;
  reg                 io_in_r_bypass_regNext_1_2_stall_9;
  reg        [15:0]   io_in_r_bypass_regNext_1_3_data_9;
  reg                 io_in_r_bypass_regNext_1_3_load_store_9;
  reg                 io_in_r_bypass_regNext_1_3_df_is_ws_9;
  reg                 io_in_r_bypass_regNext_1_3_stall_9;
  reg        [15:0]   io_in_r_bypass_regNext_2_0_data_9;
  reg                 io_in_r_bypass_regNext_2_0_load_store_9;
  reg                 io_in_r_bypass_regNext_2_0_df_is_ws_9;
  reg                 io_in_r_bypass_regNext_2_0_stall_9;
  reg        [15:0]   io_in_r_bypass_regNext_2_1_data_9;
  reg                 io_in_r_bypass_regNext_2_1_load_store_9;
  reg                 io_in_r_bypass_regNext_2_1_df_is_ws_9;
  reg                 io_in_r_bypass_regNext_2_1_stall_9;
  reg        [15:0]   io_in_r_bypass_regNext_2_2_data_9;
  reg                 io_in_r_bypass_regNext_2_2_load_store_9;
  reg                 io_in_r_bypass_regNext_2_2_df_is_ws_9;
  reg                 io_in_r_bypass_regNext_2_2_stall_9;
  reg        [15:0]   io_in_r_bypass_regNext_2_3_data_9;
  reg                 io_in_r_bypass_regNext_2_3_load_store_9;
  reg                 io_in_r_bypass_regNext_2_3_df_is_ws_9;
  reg                 io_in_r_bypass_regNext_2_3_stall_9;
  reg        [15:0]   io_in_r_bypass_regNext_3_0_data_9;
  reg                 io_in_r_bypass_regNext_3_0_load_store_9;
  reg                 io_in_r_bypass_regNext_3_0_df_is_ws_9;
  reg                 io_in_r_bypass_regNext_3_0_stall_9;
  reg        [15:0]   io_in_r_bypass_regNext_3_1_data_9;
  reg                 io_in_r_bypass_regNext_3_1_load_store_9;
  reg                 io_in_r_bypass_regNext_3_1_df_is_ws_9;
  reg                 io_in_r_bypass_regNext_3_1_stall_9;
  reg        [15:0]   io_in_r_bypass_regNext_3_2_data_9;
  reg                 io_in_r_bypass_regNext_3_2_load_store_9;
  reg                 io_in_r_bypass_regNext_3_2_df_is_ws_9;
  reg                 io_in_r_bypass_regNext_3_2_stall_9;
  reg        [15:0]   io_in_r_bypass_regNext_3_3_data_9;
  reg                 io_in_r_bypass_regNext_3_3_load_store_9;
  reg                 io_in_r_bypass_regNext_3_3_df_is_ws_9;
  reg                 io_in_r_bypass_regNext_3_3_stall_9;
  reg        [15:0]   io_in_r_bypass_regNext_4_0_data_9;
  reg                 io_in_r_bypass_regNext_4_0_load_store_9;
  reg                 io_in_r_bypass_regNext_4_0_df_is_ws_9;
  reg                 io_in_r_bypass_regNext_4_0_stall_9;
  reg        [15:0]   io_in_r_bypass_regNext_4_1_data_9;
  reg                 io_in_r_bypass_regNext_4_1_load_store_9;
  reg                 io_in_r_bypass_regNext_4_1_df_is_ws_9;
  reg                 io_in_r_bypass_regNext_4_1_stall_9;
  reg        [15:0]   io_in_r_bypass_regNext_4_2_data_9;
  reg                 io_in_r_bypass_regNext_4_2_load_store_9;
  reg                 io_in_r_bypass_regNext_4_2_df_is_ws_9;
  reg                 io_in_r_bypass_regNext_4_2_stall_9;
  reg        [15:0]   io_in_r_bypass_regNext_4_3_data_9;
  reg                 io_in_r_bypass_regNext_4_3_load_store_9;
  reg                 io_in_r_bypass_regNext_4_3_df_is_ws_9;
  reg                 io_in_r_bypass_regNext_4_3_stall_9;
  reg        [15:0]   io_in_r_bypass_regNext_5_0_data_9;
  reg                 io_in_r_bypass_regNext_5_0_load_store_9;
  reg                 io_in_r_bypass_regNext_5_0_df_is_ws_9;
  reg                 io_in_r_bypass_regNext_5_0_stall_9;
  reg        [15:0]   io_in_r_bypass_regNext_5_1_data_9;
  reg                 io_in_r_bypass_regNext_5_1_load_store_9;
  reg                 io_in_r_bypass_regNext_5_1_df_is_ws_9;
  reg                 io_in_r_bypass_regNext_5_1_stall_9;
  reg        [15:0]   io_in_r_bypass_regNext_5_2_data_9;
  reg                 io_in_r_bypass_regNext_5_2_load_store_9;
  reg                 io_in_r_bypass_regNext_5_2_df_is_ws_9;
  reg                 io_in_r_bypass_regNext_5_2_stall_9;
  reg        [15:0]   io_in_r_bypass_regNext_5_3_data_9;
  reg                 io_in_r_bypass_regNext_5_3_load_store_9;
  reg                 io_in_r_bypass_regNext_5_3_df_is_ws_9;
  reg                 io_in_r_bypass_regNext_5_3_stall_9;
  reg        [15:0]   io_in_r_bypass_regNext_6_0_data_9;
  reg                 io_in_r_bypass_regNext_6_0_load_store_9;
  reg                 io_in_r_bypass_regNext_6_0_df_is_ws_9;
  reg                 io_in_r_bypass_regNext_6_0_stall_9;
  reg        [15:0]   io_in_r_bypass_regNext_6_1_data_9;
  reg                 io_in_r_bypass_regNext_6_1_load_store_9;
  reg                 io_in_r_bypass_regNext_6_1_df_is_ws_9;
  reg                 io_in_r_bypass_regNext_6_1_stall_9;
  reg        [15:0]   io_in_r_bypass_regNext_6_2_data_9;
  reg                 io_in_r_bypass_regNext_6_2_load_store_9;
  reg                 io_in_r_bypass_regNext_6_2_df_is_ws_9;
  reg                 io_in_r_bypass_regNext_6_2_stall_9;
  reg        [15:0]   io_in_r_bypass_regNext_6_3_data_9;
  reg                 io_in_r_bypass_regNext_6_3_load_store_9;
  reg                 io_in_r_bypass_regNext_6_3_df_is_ws_9;
  reg                 io_in_r_bypass_regNext_6_3_stall_9;
  reg        [15:0]   io_in_r_bypass_regNext_7_0_data_9;
  reg                 io_in_r_bypass_regNext_7_0_load_store_9;
  reg                 io_in_r_bypass_regNext_7_0_df_is_ws_9;
  reg                 io_in_r_bypass_regNext_7_0_stall_9;
  reg        [15:0]   io_in_r_bypass_regNext_7_1_data_9;
  reg                 io_in_r_bypass_regNext_7_1_load_store_9;
  reg                 io_in_r_bypass_regNext_7_1_df_is_ws_9;
  reg                 io_in_r_bypass_regNext_7_1_stall_9;
  reg        [15:0]   io_in_r_bypass_regNext_7_2_data_9;
  reg                 io_in_r_bypass_regNext_7_2_load_store_9;
  reg                 io_in_r_bypass_regNext_7_2_df_is_ws_9;
  reg                 io_in_r_bypass_regNext_7_2_stall_9;
  reg        [15:0]   io_in_r_bypass_regNext_7_3_data_9;
  reg                 io_in_r_bypass_regNext_7_3_load_store_9;
  reg                 io_in_r_bypass_regNext_7_3_df_is_ws_9;
  reg                 io_in_r_bypass_regNext_7_3_stall_9;
  reg        [15:0]   io_in_r_bypass_regNext_8_0_data_9;
  reg                 io_in_r_bypass_regNext_8_0_load_store_9;
  reg                 io_in_r_bypass_regNext_8_0_df_is_ws_9;
  reg                 io_in_r_bypass_regNext_8_0_stall_9;
  reg        [15:0]   io_in_r_bypass_regNext_8_1_data_9;
  reg                 io_in_r_bypass_regNext_8_1_load_store_9;
  reg                 io_in_r_bypass_regNext_8_1_df_is_ws_9;
  reg                 io_in_r_bypass_regNext_8_1_stall_9;
  reg        [15:0]   io_in_r_bypass_regNext_8_2_data_9;
  reg                 io_in_r_bypass_regNext_8_2_load_store_9;
  reg                 io_in_r_bypass_regNext_8_2_df_is_ws_9;
  reg                 io_in_r_bypass_regNext_8_2_stall_9;
  reg        [15:0]   io_in_r_bypass_regNext_8_3_data_9;
  reg                 io_in_r_bypass_regNext_8_3_load_store_9;
  reg                 io_in_r_bypass_regNext_8_3_df_is_ws_9;
  reg                 io_in_r_bypass_regNext_8_3_stall_9;
  reg        [15:0]   io_in_r_bypass_regNext_9_0_data_9;
  reg                 io_in_r_bypass_regNext_9_0_load_store_9;
  reg                 io_in_r_bypass_regNext_9_0_df_is_ws_9;
  reg                 io_in_r_bypass_regNext_9_0_stall_9;
  reg        [15:0]   io_in_r_bypass_regNext_9_1_data_9;
  reg                 io_in_r_bypass_regNext_9_1_load_store_9;
  reg                 io_in_r_bypass_regNext_9_1_df_is_ws_9;
  reg                 io_in_r_bypass_regNext_9_1_stall_9;
  reg        [15:0]   io_in_r_bypass_regNext_9_2_data_9;
  reg                 io_in_r_bypass_regNext_9_2_load_store_9;
  reg                 io_in_r_bypass_regNext_9_2_df_is_ws_9;
  reg                 io_in_r_bypass_regNext_9_2_stall_9;
  reg        [15:0]   io_in_r_bypass_regNext_9_3_data_9;
  reg                 io_in_r_bypass_regNext_9_3_load_store_9;
  reg                 io_in_r_bypass_regNext_9_3_df_is_ws_9;
  reg                 io_in_r_bypass_regNext_9_3_stall_9;
  reg        [15:0]   io_in_r_bypass_regNext_10_0_data_9;
  reg                 io_in_r_bypass_regNext_10_0_load_store_9;
  reg                 io_in_r_bypass_regNext_10_0_df_is_ws_9;
  reg                 io_in_r_bypass_regNext_10_0_stall_9;
  reg        [15:0]   io_in_r_bypass_regNext_10_1_data_9;
  reg                 io_in_r_bypass_regNext_10_1_load_store_9;
  reg                 io_in_r_bypass_regNext_10_1_df_is_ws_9;
  reg                 io_in_r_bypass_regNext_10_1_stall_9;
  reg        [15:0]   io_in_r_bypass_regNext_10_2_data_9;
  reg                 io_in_r_bypass_regNext_10_2_load_store_9;
  reg                 io_in_r_bypass_regNext_10_2_df_is_ws_9;
  reg                 io_in_r_bypass_regNext_10_2_stall_9;
  reg        [15:0]   io_in_r_bypass_regNext_10_3_data_9;
  reg                 io_in_r_bypass_regNext_10_3_load_store_9;
  reg                 io_in_r_bypass_regNext_10_3_df_is_ws_9;
  reg                 io_in_r_bypass_regNext_10_3_stall_9;
  reg        [15:0]   io_in_r_bypass_regNext_11_0_data_9;
  reg                 io_in_r_bypass_regNext_11_0_load_store_9;
  reg                 io_in_r_bypass_regNext_11_0_df_is_ws_9;
  reg                 io_in_r_bypass_regNext_11_0_stall_9;
  reg        [15:0]   io_in_r_bypass_regNext_11_1_data_9;
  reg                 io_in_r_bypass_regNext_11_1_load_store_9;
  reg                 io_in_r_bypass_regNext_11_1_df_is_ws_9;
  reg                 io_in_r_bypass_regNext_11_1_stall_9;
  reg        [15:0]   io_in_r_bypass_regNext_11_2_data_9;
  reg                 io_in_r_bypass_regNext_11_2_load_store_9;
  reg                 io_in_r_bypass_regNext_11_2_df_is_ws_9;
  reg                 io_in_r_bypass_regNext_11_2_stall_9;
  reg        [15:0]   io_in_r_bypass_regNext_11_3_data_9;
  reg                 io_in_r_bypass_regNext_11_3_load_store_9;
  reg                 io_in_r_bypass_regNext_11_3_df_is_ws_9;
  reg                 io_in_r_bypass_regNext_11_3_stall_9;
  reg        [15:0]   io_in_r_bypass_regNext_12_0_data_9;
  reg                 io_in_r_bypass_regNext_12_0_load_store_9;
  reg                 io_in_r_bypass_regNext_12_0_df_is_ws_9;
  reg                 io_in_r_bypass_regNext_12_0_stall_9;
  reg        [15:0]   io_in_r_bypass_regNext_12_1_data_9;
  reg                 io_in_r_bypass_regNext_12_1_load_store_9;
  reg                 io_in_r_bypass_regNext_12_1_df_is_ws_9;
  reg                 io_in_r_bypass_regNext_12_1_stall_9;
  reg        [15:0]   io_in_r_bypass_regNext_12_2_data_9;
  reg                 io_in_r_bypass_regNext_12_2_load_store_9;
  reg                 io_in_r_bypass_regNext_12_2_df_is_ws_9;
  reg                 io_in_r_bypass_regNext_12_2_stall_9;
  reg        [15:0]   io_in_r_bypass_regNext_12_3_data_9;
  reg                 io_in_r_bypass_regNext_12_3_load_store_9;
  reg                 io_in_r_bypass_regNext_12_3_df_is_ws_9;
  reg                 io_in_r_bypass_regNext_12_3_stall_9;
  reg        [15:0]   io_in_r_bypass_regNext_13_0_data_9;
  reg                 io_in_r_bypass_regNext_13_0_load_store_9;
  reg                 io_in_r_bypass_regNext_13_0_df_is_ws_9;
  reg                 io_in_r_bypass_regNext_13_0_stall_9;
  reg        [15:0]   io_in_r_bypass_regNext_13_1_data_9;
  reg                 io_in_r_bypass_regNext_13_1_load_store_9;
  reg                 io_in_r_bypass_regNext_13_1_df_is_ws_9;
  reg                 io_in_r_bypass_regNext_13_1_stall_9;
  reg        [15:0]   io_in_r_bypass_regNext_13_2_data_9;
  reg                 io_in_r_bypass_regNext_13_2_load_store_9;
  reg                 io_in_r_bypass_regNext_13_2_df_is_ws_9;
  reg                 io_in_r_bypass_regNext_13_2_stall_9;
  reg        [15:0]   io_in_r_bypass_regNext_13_3_data_9;
  reg                 io_in_r_bypass_regNext_13_3_load_store_9;
  reg                 io_in_r_bypass_regNext_13_3_df_is_ws_9;
  reg                 io_in_r_bypass_regNext_13_3_stall_9;
  reg        [15:0]   io_in_r_bypass_regNext_14_0_data_9;
  reg                 io_in_r_bypass_regNext_14_0_load_store_9;
  reg                 io_in_r_bypass_regNext_14_0_df_is_ws_9;
  reg                 io_in_r_bypass_regNext_14_0_stall_9;
  reg        [15:0]   io_in_r_bypass_regNext_14_1_data_9;
  reg                 io_in_r_bypass_regNext_14_1_load_store_9;
  reg                 io_in_r_bypass_regNext_14_1_df_is_ws_9;
  reg                 io_in_r_bypass_regNext_14_1_stall_9;
  reg        [15:0]   io_in_r_bypass_regNext_14_2_data_9;
  reg                 io_in_r_bypass_regNext_14_2_load_store_9;
  reg                 io_in_r_bypass_regNext_14_2_df_is_ws_9;
  reg                 io_in_r_bypass_regNext_14_2_stall_9;
  reg        [15:0]   io_in_r_bypass_regNext_14_3_data_9;
  reg                 io_in_r_bypass_regNext_14_3_load_store_9;
  reg                 io_in_r_bypass_regNext_14_3_df_is_ws_9;
  reg                 io_in_r_bypass_regNext_14_3_stall_9;
  reg        [15:0]   io_in_r_bypass_regNext_15_0_data_9;
  reg                 io_in_r_bypass_regNext_15_0_load_store_9;
  reg                 io_in_r_bypass_regNext_15_0_df_is_ws_9;
  reg                 io_in_r_bypass_regNext_15_0_stall_9;
  reg        [15:0]   io_in_r_bypass_regNext_15_1_data_9;
  reg                 io_in_r_bypass_regNext_15_1_load_store_9;
  reg                 io_in_r_bypass_regNext_15_1_df_is_ws_9;
  reg                 io_in_r_bypass_regNext_15_1_stall_9;
  reg        [15:0]   io_in_r_bypass_regNext_15_2_data_9;
  reg                 io_in_r_bypass_regNext_15_2_load_store_9;
  reg                 io_in_r_bypass_regNext_15_2_df_is_ws_9;
  reg                 io_in_r_bypass_regNext_15_2_stall_9;
  reg        [15:0]   io_in_r_bypass_regNext_15_3_data_9;
  reg                 io_in_r_bypass_regNext_15_3_load_store_9;
  reg                 io_in_r_bypass_regNext_15_3_df_is_ws_9;
  reg                 io_in_r_bypass_regNext_15_3_stall_9;
  reg        [15:0]   io_in_r_bypass_regNext_16_0_data_9;
  reg                 io_in_r_bypass_regNext_16_0_load_store_9;
  reg                 io_in_r_bypass_regNext_16_0_df_is_ws_9;
  reg                 io_in_r_bypass_regNext_16_0_stall_9;
  reg        [15:0]   io_in_r_bypass_regNext_16_1_data_9;
  reg                 io_in_r_bypass_regNext_16_1_load_store_9;
  reg                 io_in_r_bypass_regNext_16_1_df_is_ws_9;
  reg                 io_in_r_bypass_regNext_16_1_stall_9;
  reg        [15:0]   io_in_r_bypass_regNext_16_2_data_9;
  reg                 io_in_r_bypass_regNext_16_2_load_store_9;
  reg                 io_in_r_bypass_regNext_16_2_df_is_ws_9;
  reg                 io_in_r_bypass_regNext_16_2_stall_9;
  reg        [15:0]   io_in_r_bypass_regNext_16_3_data_9;
  reg                 io_in_r_bypass_regNext_16_3_load_store_9;
  reg                 io_in_r_bypass_regNext_16_3_df_is_ws_9;
  reg                 io_in_r_bypass_regNext_16_3_stall_9;
  reg        [15:0]   io_in_r_bypass_regNext_17_0_data_9;
  reg                 io_in_r_bypass_regNext_17_0_load_store_9;
  reg                 io_in_r_bypass_regNext_17_0_df_is_ws_9;
  reg                 io_in_r_bypass_regNext_17_0_stall_9;
  reg        [15:0]   io_in_r_bypass_regNext_17_1_data_9;
  reg                 io_in_r_bypass_regNext_17_1_load_store_9;
  reg                 io_in_r_bypass_regNext_17_1_df_is_ws_9;
  reg                 io_in_r_bypass_regNext_17_1_stall_9;
  reg        [15:0]   io_in_r_bypass_regNext_17_2_data_9;
  reg                 io_in_r_bypass_regNext_17_2_load_store_9;
  reg                 io_in_r_bypass_regNext_17_2_df_is_ws_9;
  reg                 io_in_r_bypass_regNext_17_2_stall_9;
  reg        [15:0]   io_in_r_bypass_regNext_17_3_data_9;
  reg                 io_in_r_bypass_regNext_17_3_load_store_9;
  reg                 io_in_r_bypass_regNext_17_3_df_is_ws_9;
  reg                 io_in_r_bypass_regNext_17_3_stall_9;
  reg        [15:0]   io_in_r_bypass_regNext_18_0_data_9;
  reg                 io_in_r_bypass_regNext_18_0_load_store_9;
  reg                 io_in_r_bypass_regNext_18_0_df_is_ws_9;
  reg                 io_in_r_bypass_regNext_18_0_stall_9;
  reg        [15:0]   io_in_r_bypass_regNext_18_1_data_9;
  reg                 io_in_r_bypass_regNext_18_1_load_store_9;
  reg                 io_in_r_bypass_regNext_18_1_df_is_ws_9;
  reg                 io_in_r_bypass_regNext_18_1_stall_9;
  reg        [15:0]   io_in_r_bypass_regNext_18_2_data_9;
  reg                 io_in_r_bypass_regNext_18_2_load_store_9;
  reg                 io_in_r_bypass_regNext_18_2_df_is_ws_9;
  reg                 io_in_r_bypass_regNext_18_2_stall_9;
  reg        [15:0]   io_in_r_bypass_regNext_18_3_data_9;
  reg                 io_in_r_bypass_regNext_18_3_load_store_9;
  reg                 io_in_r_bypass_regNext_18_3_df_is_ws_9;
  reg                 io_in_r_bypass_regNext_18_3_stall_9;
  reg        [15:0]   io_in_r_bypass_regNext_19_0_data_9;
  reg                 io_in_r_bypass_regNext_19_0_load_store_9;
  reg                 io_in_r_bypass_regNext_19_0_df_is_ws_9;
  reg                 io_in_r_bypass_regNext_19_0_stall_9;
  reg        [15:0]   io_in_r_bypass_regNext_19_1_data_9;
  reg                 io_in_r_bypass_regNext_19_1_load_store_9;
  reg                 io_in_r_bypass_regNext_19_1_df_is_ws_9;
  reg                 io_in_r_bypass_regNext_19_1_stall_9;
  reg        [15:0]   io_in_r_bypass_regNext_19_2_data_9;
  reg                 io_in_r_bypass_regNext_19_2_load_store_9;
  reg                 io_in_r_bypass_regNext_19_2_df_is_ws_9;
  reg                 io_in_r_bypass_regNext_19_2_stall_9;
  reg        [15:0]   io_in_r_bypass_regNext_19_3_data_9;
  reg                 io_in_r_bypass_regNext_19_3_load_store_9;
  reg                 io_in_r_bypass_regNext_19_3_df_is_ws_9;
  reg                 io_in_r_bypass_regNext_19_3_stall_9;
  reg        [15:0]   io_in_r_bypass_regNext_20_0_data_9;
  reg                 io_in_r_bypass_regNext_20_0_load_store_9;
  reg                 io_in_r_bypass_regNext_20_0_df_is_ws_9;
  reg                 io_in_r_bypass_regNext_20_0_stall_9;
  reg        [15:0]   io_in_r_bypass_regNext_20_1_data_9;
  reg                 io_in_r_bypass_regNext_20_1_load_store_9;
  reg                 io_in_r_bypass_regNext_20_1_df_is_ws_9;
  reg                 io_in_r_bypass_regNext_20_1_stall_9;
  reg        [15:0]   io_in_r_bypass_regNext_20_2_data_9;
  reg                 io_in_r_bypass_regNext_20_2_load_store_9;
  reg                 io_in_r_bypass_regNext_20_2_df_is_ws_9;
  reg                 io_in_r_bypass_regNext_20_2_stall_9;
  reg        [15:0]   io_in_r_bypass_regNext_20_3_data_9;
  reg                 io_in_r_bypass_regNext_20_3_load_store_9;
  reg                 io_in_r_bypass_regNext_20_3_df_is_ws_9;
  reg                 io_in_r_bypass_regNext_20_3_stall_9;
  reg        [15:0]   io_in_r_bypass_regNext_21_0_data_9;
  reg                 io_in_r_bypass_regNext_21_0_load_store_9;
  reg                 io_in_r_bypass_regNext_21_0_df_is_ws_9;
  reg                 io_in_r_bypass_regNext_21_0_stall_9;
  reg        [15:0]   io_in_r_bypass_regNext_21_1_data_9;
  reg                 io_in_r_bypass_regNext_21_1_load_store_9;
  reg                 io_in_r_bypass_regNext_21_1_df_is_ws_9;
  reg                 io_in_r_bypass_regNext_21_1_stall_9;
  reg        [15:0]   io_in_r_bypass_regNext_21_2_data_9;
  reg                 io_in_r_bypass_regNext_21_2_load_store_9;
  reg                 io_in_r_bypass_regNext_21_2_df_is_ws_9;
  reg                 io_in_r_bypass_regNext_21_2_stall_9;
  reg        [15:0]   io_in_r_bypass_regNext_21_3_data_9;
  reg                 io_in_r_bypass_regNext_21_3_load_store_9;
  reg                 io_in_r_bypass_regNext_21_3_df_is_ws_9;
  reg                 io_in_r_bypass_regNext_21_3_stall_9;
  reg        [15:0]   io_in_r_bypass_regNext_22_0_data_9;
  reg                 io_in_r_bypass_regNext_22_0_load_store_9;
  reg                 io_in_r_bypass_regNext_22_0_df_is_ws_9;
  reg                 io_in_r_bypass_regNext_22_0_stall_9;
  reg        [15:0]   io_in_r_bypass_regNext_22_1_data_9;
  reg                 io_in_r_bypass_regNext_22_1_load_store_9;
  reg                 io_in_r_bypass_regNext_22_1_df_is_ws_9;
  reg                 io_in_r_bypass_regNext_22_1_stall_9;
  reg        [15:0]   io_in_r_bypass_regNext_22_2_data_9;
  reg                 io_in_r_bypass_regNext_22_2_load_store_9;
  reg                 io_in_r_bypass_regNext_22_2_df_is_ws_9;
  reg                 io_in_r_bypass_regNext_22_2_stall_9;
  reg        [15:0]   io_in_r_bypass_regNext_22_3_data_9;
  reg                 io_in_r_bypass_regNext_22_3_load_store_9;
  reg                 io_in_r_bypass_regNext_22_3_df_is_ws_9;
  reg                 io_in_r_bypass_regNext_22_3_stall_9;
  reg        [15:0]   io_in_r_bypass_regNext_23_0_data_9;
  reg                 io_in_r_bypass_regNext_23_0_load_store_9;
  reg                 io_in_r_bypass_regNext_23_0_df_is_ws_9;
  reg                 io_in_r_bypass_regNext_23_0_stall_9;
  reg        [15:0]   io_in_r_bypass_regNext_23_1_data_9;
  reg                 io_in_r_bypass_regNext_23_1_load_store_9;
  reg                 io_in_r_bypass_regNext_23_1_df_is_ws_9;
  reg                 io_in_r_bypass_regNext_23_1_stall_9;
  reg        [15:0]   io_in_r_bypass_regNext_23_2_data_9;
  reg                 io_in_r_bypass_regNext_23_2_load_store_9;
  reg                 io_in_r_bypass_regNext_23_2_df_is_ws_9;
  reg                 io_in_r_bypass_regNext_23_2_stall_9;
  reg        [15:0]   io_in_r_bypass_regNext_23_3_data_9;
  reg                 io_in_r_bypass_regNext_23_3_load_store_9;
  reg                 io_in_r_bypass_regNext_23_3_df_is_ws_9;
  reg                 io_in_r_bypass_regNext_23_3_stall_9;
  reg        [15:0]   io_in_r_bypass_regNext_24_0_data_9;
  reg                 io_in_r_bypass_regNext_24_0_load_store_9;
  reg                 io_in_r_bypass_regNext_24_0_df_is_ws_9;
  reg                 io_in_r_bypass_regNext_24_0_stall_9;
  reg        [15:0]   io_in_r_bypass_regNext_24_1_data_9;
  reg                 io_in_r_bypass_regNext_24_1_load_store_9;
  reg                 io_in_r_bypass_regNext_24_1_df_is_ws_9;
  reg                 io_in_r_bypass_regNext_24_1_stall_9;
  reg        [15:0]   io_in_r_bypass_regNext_24_2_data_9;
  reg                 io_in_r_bypass_regNext_24_2_load_store_9;
  reg                 io_in_r_bypass_regNext_24_2_df_is_ws_9;
  reg                 io_in_r_bypass_regNext_24_2_stall_9;
  reg        [15:0]   io_in_r_bypass_regNext_24_3_data_9;
  reg                 io_in_r_bypass_regNext_24_3_load_store_9;
  reg                 io_in_r_bypass_regNext_24_3_df_is_ws_9;
  reg                 io_in_r_bypass_regNext_24_3_stall_9;
  reg        [15:0]   io_in_r_bypass_regNext_25_0_data_9;
  reg                 io_in_r_bypass_regNext_25_0_load_store_9;
  reg                 io_in_r_bypass_regNext_25_0_df_is_ws_9;
  reg                 io_in_r_bypass_regNext_25_0_stall_9;
  reg        [15:0]   io_in_r_bypass_regNext_25_1_data_9;
  reg                 io_in_r_bypass_regNext_25_1_load_store_9;
  reg                 io_in_r_bypass_regNext_25_1_df_is_ws_9;
  reg                 io_in_r_bypass_regNext_25_1_stall_9;
  reg        [15:0]   io_in_r_bypass_regNext_25_2_data_9;
  reg                 io_in_r_bypass_regNext_25_2_load_store_9;
  reg                 io_in_r_bypass_regNext_25_2_df_is_ws_9;
  reg                 io_in_r_bypass_regNext_25_2_stall_9;
  reg        [15:0]   io_in_r_bypass_regNext_25_3_data_9;
  reg                 io_in_r_bypass_regNext_25_3_load_store_9;
  reg                 io_in_r_bypass_regNext_25_3_df_is_ws_9;
  reg                 io_in_r_bypass_regNext_25_3_stall_9;
  reg        [15:0]   io_in_r_bypass_regNext_26_0_data_9;
  reg                 io_in_r_bypass_regNext_26_0_load_store_9;
  reg                 io_in_r_bypass_regNext_26_0_df_is_ws_9;
  reg                 io_in_r_bypass_regNext_26_0_stall_9;
  reg        [15:0]   io_in_r_bypass_regNext_26_1_data_9;
  reg                 io_in_r_bypass_regNext_26_1_load_store_9;
  reg                 io_in_r_bypass_regNext_26_1_df_is_ws_9;
  reg                 io_in_r_bypass_regNext_26_1_stall_9;
  reg        [15:0]   io_in_r_bypass_regNext_26_2_data_9;
  reg                 io_in_r_bypass_regNext_26_2_load_store_9;
  reg                 io_in_r_bypass_regNext_26_2_df_is_ws_9;
  reg                 io_in_r_bypass_regNext_26_2_stall_9;
  reg        [15:0]   io_in_r_bypass_regNext_26_3_data_9;
  reg                 io_in_r_bypass_regNext_26_3_load_store_9;
  reg                 io_in_r_bypass_regNext_26_3_df_is_ws_9;
  reg                 io_in_r_bypass_regNext_26_3_stall_9;
  reg        [15:0]   io_in_r_bypass_regNext_27_0_data_9;
  reg                 io_in_r_bypass_regNext_27_0_load_store_9;
  reg                 io_in_r_bypass_regNext_27_0_df_is_ws_9;
  reg                 io_in_r_bypass_regNext_27_0_stall_9;
  reg        [15:0]   io_in_r_bypass_regNext_27_1_data_9;
  reg                 io_in_r_bypass_regNext_27_1_load_store_9;
  reg                 io_in_r_bypass_regNext_27_1_df_is_ws_9;
  reg                 io_in_r_bypass_regNext_27_1_stall_9;
  reg        [15:0]   io_in_r_bypass_regNext_27_2_data_9;
  reg                 io_in_r_bypass_regNext_27_2_load_store_9;
  reg                 io_in_r_bypass_regNext_27_2_df_is_ws_9;
  reg                 io_in_r_bypass_regNext_27_2_stall_9;
  reg        [15:0]   io_in_r_bypass_regNext_27_3_data_9;
  reg                 io_in_r_bypass_regNext_27_3_load_store_9;
  reg                 io_in_r_bypass_regNext_27_3_df_is_ws_9;
  reg                 io_in_r_bypass_regNext_27_3_stall_9;
  reg        [15:0]   io_in_r_bypass_regNext_28_0_data_9;
  reg                 io_in_r_bypass_regNext_28_0_load_store_9;
  reg                 io_in_r_bypass_regNext_28_0_df_is_ws_9;
  reg                 io_in_r_bypass_regNext_28_0_stall_9;
  reg        [15:0]   io_in_r_bypass_regNext_28_1_data_9;
  reg                 io_in_r_bypass_regNext_28_1_load_store_9;
  reg                 io_in_r_bypass_regNext_28_1_df_is_ws_9;
  reg                 io_in_r_bypass_regNext_28_1_stall_9;
  reg        [15:0]   io_in_r_bypass_regNext_28_2_data_9;
  reg                 io_in_r_bypass_regNext_28_2_load_store_9;
  reg                 io_in_r_bypass_regNext_28_2_df_is_ws_9;
  reg                 io_in_r_bypass_regNext_28_2_stall_9;
  reg        [15:0]   io_in_r_bypass_regNext_28_3_data_9;
  reg                 io_in_r_bypass_regNext_28_3_load_store_9;
  reg                 io_in_r_bypass_regNext_28_3_df_is_ws_9;
  reg                 io_in_r_bypass_regNext_28_3_stall_9;
  reg        [15:0]   io_in_r_bypass_regNext_29_0_data_9;
  reg                 io_in_r_bypass_regNext_29_0_load_store_9;
  reg                 io_in_r_bypass_regNext_29_0_df_is_ws_9;
  reg                 io_in_r_bypass_regNext_29_0_stall_9;
  reg        [15:0]   io_in_r_bypass_regNext_29_1_data_9;
  reg                 io_in_r_bypass_regNext_29_1_load_store_9;
  reg                 io_in_r_bypass_regNext_29_1_df_is_ws_9;
  reg                 io_in_r_bypass_regNext_29_1_stall_9;
  reg        [15:0]   io_in_r_bypass_regNext_29_2_data_9;
  reg                 io_in_r_bypass_regNext_29_2_load_store_9;
  reg                 io_in_r_bypass_regNext_29_2_df_is_ws_9;
  reg                 io_in_r_bypass_regNext_29_2_stall_9;
  reg        [15:0]   io_in_r_bypass_regNext_29_3_data_9;
  reg                 io_in_r_bypass_regNext_29_3_load_store_9;
  reg                 io_in_r_bypass_regNext_29_3_df_is_ws_9;
  reg                 io_in_r_bypass_regNext_29_3_stall_9;
  reg        [15:0]   io_in_r_bypass_regNext_30_0_data_9;
  reg                 io_in_r_bypass_regNext_30_0_load_store_9;
  reg                 io_in_r_bypass_regNext_30_0_df_is_ws_9;
  reg                 io_in_r_bypass_regNext_30_0_stall_9;
  reg        [15:0]   io_in_r_bypass_regNext_30_1_data_9;
  reg                 io_in_r_bypass_regNext_30_1_load_store_9;
  reg                 io_in_r_bypass_regNext_30_1_df_is_ws_9;
  reg                 io_in_r_bypass_regNext_30_1_stall_9;
  reg        [15:0]   io_in_r_bypass_regNext_30_2_data_9;
  reg                 io_in_r_bypass_regNext_30_2_load_store_9;
  reg                 io_in_r_bypass_regNext_30_2_df_is_ws_9;
  reg                 io_in_r_bypass_regNext_30_2_stall_9;
  reg        [15:0]   io_in_r_bypass_regNext_30_3_data_9;
  reg                 io_in_r_bypass_regNext_30_3_load_store_9;
  reg                 io_in_r_bypass_regNext_30_3_df_is_ws_9;
  reg                 io_in_r_bypass_regNext_30_3_stall_9;
  reg        [15:0]   io_in_r_bypass_regNext_31_0_data_9;
  reg                 io_in_r_bypass_regNext_31_0_load_store_9;
  reg                 io_in_r_bypass_regNext_31_0_df_is_ws_9;
  reg                 io_in_r_bypass_regNext_31_0_stall_9;
  reg        [15:0]   io_in_r_bypass_regNext_31_1_data_9;
  reg                 io_in_r_bypass_regNext_31_1_load_store_9;
  reg                 io_in_r_bypass_regNext_31_1_df_is_ws_9;
  reg                 io_in_r_bypass_regNext_31_1_stall_9;
  reg        [15:0]   io_in_r_bypass_regNext_31_2_data_9;
  reg                 io_in_r_bypass_regNext_31_2_load_store_9;
  reg                 io_in_r_bypass_regNext_31_2_df_is_ws_9;
  reg                 io_in_r_bypass_regNext_31_2_stall_9;
  reg        [15:0]   io_in_r_bypass_regNext_31_3_data_9;
  reg                 io_in_r_bypass_regNext_31_3_load_store_9;
  reg                 io_in_r_bypass_regNext_31_3_df_is_ws_9;
  reg                 io_in_r_bypass_regNext_31_3_stall_9;
  reg        [15:0]   io_in_r_bypass_regNext_0_0_data_10;
  reg                 io_in_r_bypass_regNext_0_0_load_store_10;
  reg                 io_in_r_bypass_regNext_0_0_df_is_ws_10;
  reg                 io_in_r_bypass_regNext_0_0_stall_10;
  reg        [15:0]   io_in_r_bypass_regNext_0_1_data_10;
  reg                 io_in_r_bypass_regNext_0_1_load_store_10;
  reg                 io_in_r_bypass_regNext_0_1_df_is_ws_10;
  reg                 io_in_r_bypass_regNext_0_1_stall_10;
  reg        [15:0]   io_in_r_bypass_regNext_0_2_data_10;
  reg                 io_in_r_bypass_regNext_0_2_load_store_10;
  reg                 io_in_r_bypass_regNext_0_2_df_is_ws_10;
  reg                 io_in_r_bypass_regNext_0_2_stall_10;
  reg        [15:0]   io_in_r_bypass_regNext_0_3_data_10;
  reg                 io_in_r_bypass_regNext_0_3_load_store_10;
  reg                 io_in_r_bypass_regNext_0_3_df_is_ws_10;
  reg                 io_in_r_bypass_regNext_0_3_stall_10;
  reg        [15:0]   io_in_r_bypass_regNext_1_0_data_10;
  reg                 io_in_r_bypass_regNext_1_0_load_store_10;
  reg                 io_in_r_bypass_regNext_1_0_df_is_ws_10;
  reg                 io_in_r_bypass_regNext_1_0_stall_10;
  reg        [15:0]   io_in_r_bypass_regNext_1_1_data_10;
  reg                 io_in_r_bypass_regNext_1_1_load_store_10;
  reg                 io_in_r_bypass_regNext_1_1_df_is_ws_10;
  reg                 io_in_r_bypass_regNext_1_1_stall_10;
  reg        [15:0]   io_in_r_bypass_regNext_1_2_data_10;
  reg                 io_in_r_bypass_regNext_1_2_load_store_10;
  reg                 io_in_r_bypass_regNext_1_2_df_is_ws_10;
  reg                 io_in_r_bypass_regNext_1_2_stall_10;
  reg        [15:0]   io_in_r_bypass_regNext_1_3_data_10;
  reg                 io_in_r_bypass_regNext_1_3_load_store_10;
  reg                 io_in_r_bypass_regNext_1_3_df_is_ws_10;
  reg                 io_in_r_bypass_regNext_1_3_stall_10;
  reg        [15:0]   io_in_r_bypass_regNext_2_0_data_10;
  reg                 io_in_r_bypass_regNext_2_0_load_store_10;
  reg                 io_in_r_bypass_regNext_2_0_df_is_ws_10;
  reg                 io_in_r_bypass_regNext_2_0_stall_10;
  reg        [15:0]   io_in_r_bypass_regNext_2_1_data_10;
  reg                 io_in_r_bypass_regNext_2_1_load_store_10;
  reg                 io_in_r_bypass_regNext_2_1_df_is_ws_10;
  reg                 io_in_r_bypass_regNext_2_1_stall_10;
  reg        [15:0]   io_in_r_bypass_regNext_2_2_data_10;
  reg                 io_in_r_bypass_regNext_2_2_load_store_10;
  reg                 io_in_r_bypass_regNext_2_2_df_is_ws_10;
  reg                 io_in_r_bypass_regNext_2_2_stall_10;
  reg        [15:0]   io_in_r_bypass_regNext_2_3_data_10;
  reg                 io_in_r_bypass_regNext_2_3_load_store_10;
  reg                 io_in_r_bypass_regNext_2_3_df_is_ws_10;
  reg                 io_in_r_bypass_regNext_2_3_stall_10;
  reg        [15:0]   io_in_r_bypass_regNext_3_0_data_10;
  reg                 io_in_r_bypass_regNext_3_0_load_store_10;
  reg                 io_in_r_bypass_regNext_3_0_df_is_ws_10;
  reg                 io_in_r_bypass_regNext_3_0_stall_10;
  reg        [15:0]   io_in_r_bypass_regNext_3_1_data_10;
  reg                 io_in_r_bypass_regNext_3_1_load_store_10;
  reg                 io_in_r_bypass_regNext_3_1_df_is_ws_10;
  reg                 io_in_r_bypass_regNext_3_1_stall_10;
  reg        [15:0]   io_in_r_bypass_regNext_3_2_data_10;
  reg                 io_in_r_bypass_regNext_3_2_load_store_10;
  reg                 io_in_r_bypass_regNext_3_2_df_is_ws_10;
  reg                 io_in_r_bypass_regNext_3_2_stall_10;
  reg        [15:0]   io_in_r_bypass_regNext_3_3_data_10;
  reg                 io_in_r_bypass_regNext_3_3_load_store_10;
  reg                 io_in_r_bypass_regNext_3_3_df_is_ws_10;
  reg                 io_in_r_bypass_regNext_3_3_stall_10;
  reg        [15:0]   io_in_r_bypass_regNext_4_0_data_10;
  reg                 io_in_r_bypass_regNext_4_0_load_store_10;
  reg                 io_in_r_bypass_regNext_4_0_df_is_ws_10;
  reg                 io_in_r_bypass_regNext_4_0_stall_10;
  reg        [15:0]   io_in_r_bypass_regNext_4_1_data_10;
  reg                 io_in_r_bypass_regNext_4_1_load_store_10;
  reg                 io_in_r_bypass_regNext_4_1_df_is_ws_10;
  reg                 io_in_r_bypass_regNext_4_1_stall_10;
  reg        [15:0]   io_in_r_bypass_regNext_4_2_data_10;
  reg                 io_in_r_bypass_regNext_4_2_load_store_10;
  reg                 io_in_r_bypass_regNext_4_2_df_is_ws_10;
  reg                 io_in_r_bypass_regNext_4_2_stall_10;
  reg        [15:0]   io_in_r_bypass_regNext_4_3_data_10;
  reg                 io_in_r_bypass_regNext_4_3_load_store_10;
  reg                 io_in_r_bypass_regNext_4_3_df_is_ws_10;
  reg                 io_in_r_bypass_regNext_4_3_stall_10;
  reg        [15:0]   io_in_r_bypass_regNext_5_0_data_10;
  reg                 io_in_r_bypass_regNext_5_0_load_store_10;
  reg                 io_in_r_bypass_regNext_5_0_df_is_ws_10;
  reg                 io_in_r_bypass_regNext_5_0_stall_10;
  reg        [15:0]   io_in_r_bypass_regNext_5_1_data_10;
  reg                 io_in_r_bypass_regNext_5_1_load_store_10;
  reg                 io_in_r_bypass_regNext_5_1_df_is_ws_10;
  reg                 io_in_r_bypass_regNext_5_1_stall_10;
  reg        [15:0]   io_in_r_bypass_regNext_5_2_data_10;
  reg                 io_in_r_bypass_regNext_5_2_load_store_10;
  reg                 io_in_r_bypass_regNext_5_2_df_is_ws_10;
  reg                 io_in_r_bypass_regNext_5_2_stall_10;
  reg        [15:0]   io_in_r_bypass_regNext_5_3_data_10;
  reg                 io_in_r_bypass_regNext_5_3_load_store_10;
  reg                 io_in_r_bypass_regNext_5_3_df_is_ws_10;
  reg                 io_in_r_bypass_regNext_5_3_stall_10;
  reg        [15:0]   io_in_r_bypass_regNext_6_0_data_10;
  reg                 io_in_r_bypass_regNext_6_0_load_store_10;
  reg                 io_in_r_bypass_regNext_6_0_df_is_ws_10;
  reg                 io_in_r_bypass_regNext_6_0_stall_10;
  reg        [15:0]   io_in_r_bypass_regNext_6_1_data_10;
  reg                 io_in_r_bypass_regNext_6_1_load_store_10;
  reg                 io_in_r_bypass_regNext_6_1_df_is_ws_10;
  reg                 io_in_r_bypass_regNext_6_1_stall_10;
  reg        [15:0]   io_in_r_bypass_regNext_6_2_data_10;
  reg                 io_in_r_bypass_regNext_6_2_load_store_10;
  reg                 io_in_r_bypass_regNext_6_2_df_is_ws_10;
  reg                 io_in_r_bypass_regNext_6_2_stall_10;
  reg        [15:0]   io_in_r_bypass_regNext_6_3_data_10;
  reg                 io_in_r_bypass_regNext_6_3_load_store_10;
  reg                 io_in_r_bypass_regNext_6_3_df_is_ws_10;
  reg                 io_in_r_bypass_regNext_6_3_stall_10;
  reg        [15:0]   io_in_r_bypass_regNext_7_0_data_10;
  reg                 io_in_r_bypass_regNext_7_0_load_store_10;
  reg                 io_in_r_bypass_regNext_7_0_df_is_ws_10;
  reg                 io_in_r_bypass_regNext_7_0_stall_10;
  reg        [15:0]   io_in_r_bypass_regNext_7_1_data_10;
  reg                 io_in_r_bypass_regNext_7_1_load_store_10;
  reg                 io_in_r_bypass_regNext_7_1_df_is_ws_10;
  reg                 io_in_r_bypass_regNext_7_1_stall_10;
  reg        [15:0]   io_in_r_bypass_regNext_7_2_data_10;
  reg                 io_in_r_bypass_regNext_7_2_load_store_10;
  reg                 io_in_r_bypass_regNext_7_2_df_is_ws_10;
  reg                 io_in_r_bypass_regNext_7_2_stall_10;
  reg        [15:0]   io_in_r_bypass_regNext_7_3_data_10;
  reg                 io_in_r_bypass_regNext_7_3_load_store_10;
  reg                 io_in_r_bypass_regNext_7_3_df_is_ws_10;
  reg                 io_in_r_bypass_regNext_7_3_stall_10;
  reg        [15:0]   io_in_r_bypass_regNext_8_0_data_10;
  reg                 io_in_r_bypass_regNext_8_0_load_store_10;
  reg                 io_in_r_bypass_regNext_8_0_df_is_ws_10;
  reg                 io_in_r_bypass_regNext_8_0_stall_10;
  reg        [15:0]   io_in_r_bypass_regNext_8_1_data_10;
  reg                 io_in_r_bypass_regNext_8_1_load_store_10;
  reg                 io_in_r_bypass_regNext_8_1_df_is_ws_10;
  reg                 io_in_r_bypass_regNext_8_1_stall_10;
  reg        [15:0]   io_in_r_bypass_regNext_8_2_data_10;
  reg                 io_in_r_bypass_regNext_8_2_load_store_10;
  reg                 io_in_r_bypass_regNext_8_2_df_is_ws_10;
  reg                 io_in_r_bypass_regNext_8_2_stall_10;
  reg        [15:0]   io_in_r_bypass_regNext_8_3_data_10;
  reg                 io_in_r_bypass_regNext_8_3_load_store_10;
  reg                 io_in_r_bypass_regNext_8_3_df_is_ws_10;
  reg                 io_in_r_bypass_regNext_8_3_stall_10;
  reg        [15:0]   io_in_r_bypass_regNext_9_0_data_10;
  reg                 io_in_r_bypass_regNext_9_0_load_store_10;
  reg                 io_in_r_bypass_regNext_9_0_df_is_ws_10;
  reg                 io_in_r_bypass_regNext_9_0_stall_10;
  reg        [15:0]   io_in_r_bypass_regNext_9_1_data_10;
  reg                 io_in_r_bypass_regNext_9_1_load_store_10;
  reg                 io_in_r_bypass_regNext_9_1_df_is_ws_10;
  reg                 io_in_r_bypass_regNext_9_1_stall_10;
  reg        [15:0]   io_in_r_bypass_regNext_9_2_data_10;
  reg                 io_in_r_bypass_regNext_9_2_load_store_10;
  reg                 io_in_r_bypass_regNext_9_2_df_is_ws_10;
  reg                 io_in_r_bypass_regNext_9_2_stall_10;
  reg        [15:0]   io_in_r_bypass_regNext_9_3_data_10;
  reg                 io_in_r_bypass_regNext_9_3_load_store_10;
  reg                 io_in_r_bypass_regNext_9_3_df_is_ws_10;
  reg                 io_in_r_bypass_regNext_9_3_stall_10;
  reg        [15:0]   io_in_r_bypass_regNext_10_0_data_10;
  reg                 io_in_r_bypass_regNext_10_0_load_store_10;
  reg                 io_in_r_bypass_regNext_10_0_df_is_ws_10;
  reg                 io_in_r_bypass_regNext_10_0_stall_10;
  reg        [15:0]   io_in_r_bypass_regNext_10_1_data_10;
  reg                 io_in_r_bypass_regNext_10_1_load_store_10;
  reg                 io_in_r_bypass_regNext_10_1_df_is_ws_10;
  reg                 io_in_r_bypass_regNext_10_1_stall_10;
  reg        [15:0]   io_in_r_bypass_regNext_10_2_data_10;
  reg                 io_in_r_bypass_regNext_10_2_load_store_10;
  reg                 io_in_r_bypass_regNext_10_2_df_is_ws_10;
  reg                 io_in_r_bypass_regNext_10_2_stall_10;
  reg        [15:0]   io_in_r_bypass_regNext_10_3_data_10;
  reg                 io_in_r_bypass_regNext_10_3_load_store_10;
  reg                 io_in_r_bypass_regNext_10_3_df_is_ws_10;
  reg                 io_in_r_bypass_regNext_10_3_stall_10;
  reg        [15:0]   io_in_r_bypass_regNext_11_0_data_10;
  reg                 io_in_r_bypass_regNext_11_0_load_store_10;
  reg                 io_in_r_bypass_regNext_11_0_df_is_ws_10;
  reg                 io_in_r_bypass_regNext_11_0_stall_10;
  reg        [15:0]   io_in_r_bypass_regNext_11_1_data_10;
  reg                 io_in_r_bypass_regNext_11_1_load_store_10;
  reg                 io_in_r_bypass_regNext_11_1_df_is_ws_10;
  reg                 io_in_r_bypass_regNext_11_1_stall_10;
  reg        [15:0]   io_in_r_bypass_regNext_11_2_data_10;
  reg                 io_in_r_bypass_regNext_11_2_load_store_10;
  reg                 io_in_r_bypass_regNext_11_2_df_is_ws_10;
  reg                 io_in_r_bypass_regNext_11_2_stall_10;
  reg        [15:0]   io_in_r_bypass_regNext_11_3_data_10;
  reg                 io_in_r_bypass_regNext_11_3_load_store_10;
  reg                 io_in_r_bypass_regNext_11_3_df_is_ws_10;
  reg                 io_in_r_bypass_regNext_11_3_stall_10;
  reg        [15:0]   io_in_r_bypass_regNext_12_0_data_10;
  reg                 io_in_r_bypass_regNext_12_0_load_store_10;
  reg                 io_in_r_bypass_regNext_12_0_df_is_ws_10;
  reg                 io_in_r_bypass_regNext_12_0_stall_10;
  reg        [15:0]   io_in_r_bypass_regNext_12_1_data_10;
  reg                 io_in_r_bypass_regNext_12_1_load_store_10;
  reg                 io_in_r_bypass_regNext_12_1_df_is_ws_10;
  reg                 io_in_r_bypass_regNext_12_1_stall_10;
  reg        [15:0]   io_in_r_bypass_regNext_12_2_data_10;
  reg                 io_in_r_bypass_regNext_12_2_load_store_10;
  reg                 io_in_r_bypass_regNext_12_2_df_is_ws_10;
  reg                 io_in_r_bypass_regNext_12_2_stall_10;
  reg        [15:0]   io_in_r_bypass_regNext_12_3_data_10;
  reg                 io_in_r_bypass_regNext_12_3_load_store_10;
  reg                 io_in_r_bypass_regNext_12_3_df_is_ws_10;
  reg                 io_in_r_bypass_regNext_12_3_stall_10;
  reg        [15:0]   io_in_r_bypass_regNext_13_0_data_10;
  reg                 io_in_r_bypass_regNext_13_0_load_store_10;
  reg                 io_in_r_bypass_regNext_13_0_df_is_ws_10;
  reg                 io_in_r_bypass_regNext_13_0_stall_10;
  reg        [15:0]   io_in_r_bypass_regNext_13_1_data_10;
  reg                 io_in_r_bypass_regNext_13_1_load_store_10;
  reg                 io_in_r_bypass_regNext_13_1_df_is_ws_10;
  reg                 io_in_r_bypass_regNext_13_1_stall_10;
  reg        [15:0]   io_in_r_bypass_regNext_13_2_data_10;
  reg                 io_in_r_bypass_regNext_13_2_load_store_10;
  reg                 io_in_r_bypass_regNext_13_2_df_is_ws_10;
  reg                 io_in_r_bypass_regNext_13_2_stall_10;
  reg        [15:0]   io_in_r_bypass_regNext_13_3_data_10;
  reg                 io_in_r_bypass_regNext_13_3_load_store_10;
  reg                 io_in_r_bypass_regNext_13_3_df_is_ws_10;
  reg                 io_in_r_bypass_regNext_13_3_stall_10;
  reg        [15:0]   io_in_r_bypass_regNext_14_0_data_10;
  reg                 io_in_r_bypass_regNext_14_0_load_store_10;
  reg                 io_in_r_bypass_regNext_14_0_df_is_ws_10;
  reg                 io_in_r_bypass_regNext_14_0_stall_10;
  reg        [15:0]   io_in_r_bypass_regNext_14_1_data_10;
  reg                 io_in_r_bypass_regNext_14_1_load_store_10;
  reg                 io_in_r_bypass_regNext_14_1_df_is_ws_10;
  reg                 io_in_r_bypass_regNext_14_1_stall_10;
  reg        [15:0]   io_in_r_bypass_regNext_14_2_data_10;
  reg                 io_in_r_bypass_regNext_14_2_load_store_10;
  reg                 io_in_r_bypass_regNext_14_2_df_is_ws_10;
  reg                 io_in_r_bypass_regNext_14_2_stall_10;
  reg        [15:0]   io_in_r_bypass_regNext_14_3_data_10;
  reg                 io_in_r_bypass_regNext_14_3_load_store_10;
  reg                 io_in_r_bypass_regNext_14_3_df_is_ws_10;
  reg                 io_in_r_bypass_regNext_14_3_stall_10;
  reg        [15:0]   io_in_r_bypass_regNext_15_0_data_10;
  reg                 io_in_r_bypass_regNext_15_0_load_store_10;
  reg                 io_in_r_bypass_regNext_15_0_df_is_ws_10;
  reg                 io_in_r_bypass_regNext_15_0_stall_10;
  reg        [15:0]   io_in_r_bypass_regNext_15_1_data_10;
  reg                 io_in_r_bypass_regNext_15_1_load_store_10;
  reg                 io_in_r_bypass_regNext_15_1_df_is_ws_10;
  reg                 io_in_r_bypass_regNext_15_1_stall_10;
  reg        [15:0]   io_in_r_bypass_regNext_15_2_data_10;
  reg                 io_in_r_bypass_regNext_15_2_load_store_10;
  reg                 io_in_r_bypass_regNext_15_2_df_is_ws_10;
  reg                 io_in_r_bypass_regNext_15_2_stall_10;
  reg        [15:0]   io_in_r_bypass_regNext_15_3_data_10;
  reg                 io_in_r_bypass_regNext_15_3_load_store_10;
  reg                 io_in_r_bypass_regNext_15_3_df_is_ws_10;
  reg                 io_in_r_bypass_regNext_15_3_stall_10;
  reg        [15:0]   io_in_r_bypass_regNext_16_0_data_10;
  reg                 io_in_r_bypass_regNext_16_0_load_store_10;
  reg                 io_in_r_bypass_regNext_16_0_df_is_ws_10;
  reg                 io_in_r_bypass_regNext_16_0_stall_10;
  reg        [15:0]   io_in_r_bypass_regNext_16_1_data_10;
  reg                 io_in_r_bypass_regNext_16_1_load_store_10;
  reg                 io_in_r_bypass_regNext_16_1_df_is_ws_10;
  reg                 io_in_r_bypass_regNext_16_1_stall_10;
  reg        [15:0]   io_in_r_bypass_regNext_16_2_data_10;
  reg                 io_in_r_bypass_regNext_16_2_load_store_10;
  reg                 io_in_r_bypass_regNext_16_2_df_is_ws_10;
  reg                 io_in_r_bypass_regNext_16_2_stall_10;
  reg        [15:0]   io_in_r_bypass_regNext_16_3_data_10;
  reg                 io_in_r_bypass_regNext_16_3_load_store_10;
  reg                 io_in_r_bypass_regNext_16_3_df_is_ws_10;
  reg                 io_in_r_bypass_regNext_16_3_stall_10;
  reg        [15:0]   io_in_r_bypass_regNext_17_0_data_10;
  reg                 io_in_r_bypass_regNext_17_0_load_store_10;
  reg                 io_in_r_bypass_regNext_17_0_df_is_ws_10;
  reg                 io_in_r_bypass_regNext_17_0_stall_10;
  reg        [15:0]   io_in_r_bypass_regNext_17_1_data_10;
  reg                 io_in_r_bypass_regNext_17_1_load_store_10;
  reg                 io_in_r_bypass_regNext_17_1_df_is_ws_10;
  reg                 io_in_r_bypass_regNext_17_1_stall_10;
  reg        [15:0]   io_in_r_bypass_regNext_17_2_data_10;
  reg                 io_in_r_bypass_regNext_17_2_load_store_10;
  reg                 io_in_r_bypass_regNext_17_2_df_is_ws_10;
  reg                 io_in_r_bypass_regNext_17_2_stall_10;
  reg        [15:0]   io_in_r_bypass_regNext_17_3_data_10;
  reg                 io_in_r_bypass_regNext_17_3_load_store_10;
  reg                 io_in_r_bypass_regNext_17_3_df_is_ws_10;
  reg                 io_in_r_bypass_regNext_17_3_stall_10;
  reg        [15:0]   io_in_r_bypass_regNext_18_0_data_10;
  reg                 io_in_r_bypass_regNext_18_0_load_store_10;
  reg                 io_in_r_bypass_regNext_18_0_df_is_ws_10;
  reg                 io_in_r_bypass_regNext_18_0_stall_10;
  reg        [15:0]   io_in_r_bypass_regNext_18_1_data_10;
  reg                 io_in_r_bypass_regNext_18_1_load_store_10;
  reg                 io_in_r_bypass_regNext_18_1_df_is_ws_10;
  reg                 io_in_r_bypass_regNext_18_1_stall_10;
  reg        [15:0]   io_in_r_bypass_regNext_18_2_data_10;
  reg                 io_in_r_bypass_regNext_18_2_load_store_10;
  reg                 io_in_r_bypass_regNext_18_2_df_is_ws_10;
  reg                 io_in_r_bypass_regNext_18_2_stall_10;
  reg        [15:0]   io_in_r_bypass_regNext_18_3_data_10;
  reg                 io_in_r_bypass_regNext_18_3_load_store_10;
  reg                 io_in_r_bypass_regNext_18_3_df_is_ws_10;
  reg                 io_in_r_bypass_regNext_18_3_stall_10;
  reg        [15:0]   io_in_r_bypass_regNext_19_0_data_10;
  reg                 io_in_r_bypass_regNext_19_0_load_store_10;
  reg                 io_in_r_bypass_regNext_19_0_df_is_ws_10;
  reg                 io_in_r_bypass_regNext_19_0_stall_10;
  reg        [15:0]   io_in_r_bypass_regNext_19_1_data_10;
  reg                 io_in_r_bypass_regNext_19_1_load_store_10;
  reg                 io_in_r_bypass_regNext_19_1_df_is_ws_10;
  reg                 io_in_r_bypass_regNext_19_1_stall_10;
  reg        [15:0]   io_in_r_bypass_regNext_19_2_data_10;
  reg                 io_in_r_bypass_regNext_19_2_load_store_10;
  reg                 io_in_r_bypass_regNext_19_2_df_is_ws_10;
  reg                 io_in_r_bypass_regNext_19_2_stall_10;
  reg        [15:0]   io_in_r_bypass_regNext_19_3_data_10;
  reg                 io_in_r_bypass_regNext_19_3_load_store_10;
  reg                 io_in_r_bypass_regNext_19_3_df_is_ws_10;
  reg                 io_in_r_bypass_regNext_19_3_stall_10;
  reg        [15:0]   io_in_r_bypass_regNext_20_0_data_10;
  reg                 io_in_r_bypass_regNext_20_0_load_store_10;
  reg                 io_in_r_bypass_regNext_20_0_df_is_ws_10;
  reg                 io_in_r_bypass_regNext_20_0_stall_10;
  reg        [15:0]   io_in_r_bypass_regNext_20_1_data_10;
  reg                 io_in_r_bypass_regNext_20_1_load_store_10;
  reg                 io_in_r_bypass_regNext_20_1_df_is_ws_10;
  reg                 io_in_r_bypass_regNext_20_1_stall_10;
  reg        [15:0]   io_in_r_bypass_regNext_20_2_data_10;
  reg                 io_in_r_bypass_regNext_20_2_load_store_10;
  reg                 io_in_r_bypass_regNext_20_2_df_is_ws_10;
  reg                 io_in_r_bypass_regNext_20_2_stall_10;
  reg        [15:0]   io_in_r_bypass_regNext_20_3_data_10;
  reg                 io_in_r_bypass_regNext_20_3_load_store_10;
  reg                 io_in_r_bypass_regNext_20_3_df_is_ws_10;
  reg                 io_in_r_bypass_regNext_20_3_stall_10;
  reg        [15:0]   io_in_r_bypass_regNext_21_0_data_10;
  reg                 io_in_r_bypass_regNext_21_0_load_store_10;
  reg                 io_in_r_bypass_regNext_21_0_df_is_ws_10;
  reg                 io_in_r_bypass_regNext_21_0_stall_10;
  reg        [15:0]   io_in_r_bypass_regNext_21_1_data_10;
  reg                 io_in_r_bypass_regNext_21_1_load_store_10;
  reg                 io_in_r_bypass_regNext_21_1_df_is_ws_10;
  reg                 io_in_r_bypass_regNext_21_1_stall_10;
  reg        [15:0]   io_in_r_bypass_regNext_21_2_data_10;
  reg                 io_in_r_bypass_regNext_21_2_load_store_10;
  reg                 io_in_r_bypass_regNext_21_2_df_is_ws_10;
  reg                 io_in_r_bypass_regNext_21_2_stall_10;
  reg        [15:0]   io_in_r_bypass_regNext_21_3_data_10;
  reg                 io_in_r_bypass_regNext_21_3_load_store_10;
  reg                 io_in_r_bypass_regNext_21_3_df_is_ws_10;
  reg                 io_in_r_bypass_regNext_21_3_stall_10;
  reg        [15:0]   io_in_r_bypass_regNext_22_0_data_10;
  reg                 io_in_r_bypass_regNext_22_0_load_store_10;
  reg                 io_in_r_bypass_regNext_22_0_df_is_ws_10;
  reg                 io_in_r_bypass_regNext_22_0_stall_10;
  reg        [15:0]   io_in_r_bypass_regNext_22_1_data_10;
  reg                 io_in_r_bypass_regNext_22_1_load_store_10;
  reg                 io_in_r_bypass_regNext_22_1_df_is_ws_10;
  reg                 io_in_r_bypass_regNext_22_1_stall_10;
  reg        [15:0]   io_in_r_bypass_regNext_22_2_data_10;
  reg                 io_in_r_bypass_regNext_22_2_load_store_10;
  reg                 io_in_r_bypass_regNext_22_2_df_is_ws_10;
  reg                 io_in_r_bypass_regNext_22_2_stall_10;
  reg        [15:0]   io_in_r_bypass_regNext_22_3_data_10;
  reg                 io_in_r_bypass_regNext_22_3_load_store_10;
  reg                 io_in_r_bypass_regNext_22_3_df_is_ws_10;
  reg                 io_in_r_bypass_regNext_22_3_stall_10;
  reg        [15:0]   io_in_r_bypass_regNext_23_0_data_10;
  reg                 io_in_r_bypass_regNext_23_0_load_store_10;
  reg                 io_in_r_bypass_regNext_23_0_df_is_ws_10;
  reg                 io_in_r_bypass_regNext_23_0_stall_10;
  reg        [15:0]   io_in_r_bypass_regNext_23_1_data_10;
  reg                 io_in_r_bypass_regNext_23_1_load_store_10;
  reg                 io_in_r_bypass_regNext_23_1_df_is_ws_10;
  reg                 io_in_r_bypass_regNext_23_1_stall_10;
  reg        [15:0]   io_in_r_bypass_regNext_23_2_data_10;
  reg                 io_in_r_bypass_regNext_23_2_load_store_10;
  reg                 io_in_r_bypass_regNext_23_2_df_is_ws_10;
  reg                 io_in_r_bypass_regNext_23_2_stall_10;
  reg        [15:0]   io_in_r_bypass_regNext_23_3_data_10;
  reg                 io_in_r_bypass_regNext_23_3_load_store_10;
  reg                 io_in_r_bypass_regNext_23_3_df_is_ws_10;
  reg                 io_in_r_bypass_regNext_23_3_stall_10;
  reg        [15:0]   io_in_r_bypass_regNext_24_0_data_10;
  reg                 io_in_r_bypass_regNext_24_0_load_store_10;
  reg                 io_in_r_bypass_regNext_24_0_df_is_ws_10;
  reg                 io_in_r_bypass_regNext_24_0_stall_10;
  reg        [15:0]   io_in_r_bypass_regNext_24_1_data_10;
  reg                 io_in_r_bypass_regNext_24_1_load_store_10;
  reg                 io_in_r_bypass_regNext_24_1_df_is_ws_10;
  reg                 io_in_r_bypass_regNext_24_1_stall_10;
  reg        [15:0]   io_in_r_bypass_regNext_24_2_data_10;
  reg                 io_in_r_bypass_regNext_24_2_load_store_10;
  reg                 io_in_r_bypass_regNext_24_2_df_is_ws_10;
  reg                 io_in_r_bypass_regNext_24_2_stall_10;
  reg        [15:0]   io_in_r_bypass_regNext_24_3_data_10;
  reg                 io_in_r_bypass_regNext_24_3_load_store_10;
  reg                 io_in_r_bypass_regNext_24_3_df_is_ws_10;
  reg                 io_in_r_bypass_regNext_24_3_stall_10;
  reg        [15:0]   io_in_r_bypass_regNext_25_0_data_10;
  reg                 io_in_r_bypass_regNext_25_0_load_store_10;
  reg                 io_in_r_bypass_regNext_25_0_df_is_ws_10;
  reg                 io_in_r_bypass_regNext_25_0_stall_10;
  reg        [15:0]   io_in_r_bypass_regNext_25_1_data_10;
  reg                 io_in_r_bypass_regNext_25_1_load_store_10;
  reg                 io_in_r_bypass_regNext_25_1_df_is_ws_10;
  reg                 io_in_r_bypass_regNext_25_1_stall_10;
  reg        [15:0]   io_in_r_bypass_regNext_25_2_data_10;
  reg                 io_in_r_bypass_regNext_25_2_load_store_10;
  reg                 io_in_r_bypass_regNext_25_2_df_is_ws_10;
  reg                 io_in_r_bypass_regNext_25_2_stall_10;
  reg        [15:0]   io_in_r_bypass_regNext_25_3_data_10;
  reg                 io_in_r_bypass_regNext_25_3_load_store_10;
  reg                 io_in_r_bypass_regNext_25_3_df_is_ws_10;
  reg                 io_in_r_bypass_regNext_25_3_stall_10;
  reg        [15:0]   io_in_r_bypass_regNext_26_0_data_10;
  reg                 io_in_r_bypass_regNext_26_0_load_store_10;
  reg                 io_in_r_bypass_regNext_26_0_df_is_ws_10;
  reg                 io_in_r_bypass_regNext_26_0_stall_10;
  reg        [15:0]   io_in_r_bypass_regNext_26_1_data_10;
  reg                 io_in_r_bypass_regNext_26_1_load_store_10;
  reg                 io_in_r_bypass_regNext_26_1_df_is_ws_10;
  reg                 io_in_r_bypass_regNext_26_1_stall_10;
  reg        [15:0]   io_in_r_bypass_regNext_26_2_data_10;
  reg                 io_in_r_bypass_regNext_26_2_load_store_10;
  reg                 io_in_r_bypass_regNext_26_2_df_is_ws_10;
  reg                 io_in_r_bypass_regNext_26_2_stall_10;
  reg        [15:0]   io_in_r_bypass_regNext_26_3_data_10;
  reg                 io_in_r_bypass_regNext_26_3_load_store_10;
  reg                 io_in_r_bypass_regNext_26_3_df_is_ws_10;
  reg                 io_in_r_bypass_regNext_26_3_stall_10;
  reg        [15:0]   io_in_r_bypass_regNext_27_0_data_10;
  reg                 io_in_r_bypass_regNext_27_0_load_store_10;
  reg                 io_in_r_bypass_regNext_27_0_df_is_ws_10;
  reg                 io_in_r_bypass_regNext_27_0_stall_10;
  reg        [15:0]   io_in_r_bypass_regNext_27_1_data_10;
  reg                 io_in_r_bypass_regNext_27_1_load_store_10;
  reg                 io_in_r_bypass_regNext_27_1_df_is_ws_10;
  reg                 io_in_r_bypass_regNext_27_1_stall_10;
  reg        [15:0]   io_in_r_bypass_regNext_27_2_data_10;
  reg                 io_in_r_bypass_regNext_27_2_load_store_10;
  reg                 io_in_r_bypass_regNext_27_2_df_is_ws_10;
  reg                 io_in_r_bypass_regNext_27_2_stall_10;
  reg        [15:0]   io_in_r_bypass_regNext_27_3_data_10;
  reg                 io_in_r_bypass_regNext_27_3_load_store_10;
  reg                 io_in_r_bypass_regNext_27_3_df_is_ws_10;
  reg                 io_in_r_bypass_regNext_27_3_stall_10;
  reg        [15:0]   io_in_r_bypass_regNext_28_0_data_10;
  reg                 io_in_r_bypass_regNext_28_0_load_store_10;
  reg                 io_in_r_bypass_regNext_28_0_df_is_ws_10;
  reg                 io_in_r_bypass_regNext_28_0_stall_10;
  reg        [15:0]   io_in_r_bypass_regNext_28_1_data_10;
  reg                 io_in_r_bypass_regNext_28_1_load_store_10;
  reg                 io_in_r_bypass_regNext_28_1_df_is_ws_10;
  reg                 io_in_r_bypass_regNext_28_1_stall_10;
  reg        [15:0]   io_in_r_bypass_regNext_28_2_data_10;
  reg                 io_in_r_bypass_regNext_28_2_load_store_10;
  reg                 io_in_r_bypass_regNext_28_2_df_is_ws_10;
  reg                 io_in_r_bypass_regNext_28_2_stall_10;
  reg        [15:0]   io_in_r_bypass_regNext_28_3_data_10;
  reg                 io_in_r_bypass_regNext_28_3_load_store_10;
  reg                 io_in_r_bypass_regNext_28_3_df_is_ws_10;
  reg                 io_in_r_bypass_regNext_28_3_stall_10;
  reg        [15:0]   io_in_r_bypass_regNext_29_0_data_10;
  reg                 io_in_r_bypass_regNext_29_0_load_store_10;
  reg                 io_in_r_bypass_regNext_29_0_df_is_ws_10;
  reg                 io_in_r_bypass_regNext_29_0_stall_10;
  reg        [15:0]   io_in_r_bypass_regNext_29_1_data_10;
  reg                 io_in_r_bypass_regNext_29_1_load_store_10;
  reg                 io_in_r_bypass_regNext_29_1_df_is_ws_10;
  reg                 io_in_r_bypass_regNext_29_1_stall_10;
  reg        [15:0]   io_in_r_bypass_regNext_29_2_data_10;
  reg                 io_in_r_bypass_regNext_29_2_load_store_10;
  reg                 io_in_r_bypass_regNext_29_2_df_is_ws_10;
  reg                 io_in_r_bypass_regNext_29_2_stall_10;
  reg        [15:0]   io_in_r_bypass_regNext_29_3_data_10;
  reg                 io_in_r_bypass_regNext_29_3_load_store_10;
  reg                 io_in_r_bypass_regNext_29_3_df_is_ws_10;
  reg                 io_in_r_bypass_regNext_29_3_stall_10;
  reg        [15:0]   io_in_r_bypass_regNext_30_0_data_10;
  reg                 io_in_r_bypass_regNext_30_0_load_store_10;
  reg                 io_in_r_bypass_regNext_30_0_df_is_ws_10;
  reg                 io_in_r_bypass_regNext_30_0_stall_10;
  reg        [15:0]   io_in_r_bypass_regNext_30_1_data_10;
  reg                 io_in_r_bypass_regNext_30_1_load_store_10;
  reg                 io_in_r_bypass_regNext_30_1_df_is_ws_10;
  reg                 io_in_r_bypass_regNext_30_1_stall_10;
  reg        [15:0]   io_in_r_bypass_regNext_30_2_data_10;
  reg                 io_in_r_bypass_regNext_30_2_load_store_10;
  reg                 io_in_r_bypass_regNext_30_2_df_is_ws_10;
  reg                 io_in_r_bypass_regNext_30_2_stall_10;
  reg        [15:0]   io_in_r_bypass_regNext_30_3_data_10;
  reg                 io_in_r_bypass_regNext_30_3_load_store_10;
  reg                 io_in_r_bypass_regNext_30_3_df_is_ws_10;
  reg                 io_in_r_bypass_regNext_30_3_stall_10;
  reg        [15:0]   io_in_r_bypass_regNext_31_0_data_10;
  reg                 io_in_r_bypass_regNext_31_0_load_store_10;
  reg                 io_in_r_bypass_regNext_31_0_df_is_ws_10;
  reg                 io_in_r_bypass_regNext_31_0_stall_10;
  reg        [15:0]   io_in_r_bypass_regNext_31_1_data_10;
  reg                 io_in_r_bypass_regNext_31_1_load_store_10;
  reg                 io_in_r_bypass_regNext_31_1_df_is_ws_10;
  reg                 io_in_r_bypass_regNext_31_1_stall_10;
  reg        [15:0]   io_in_r_bypass_regNext_31_2_data_10;
  reg                 io_in_r_bypass_regNext_31_2_load_store_10;
  reg                 io_in_r_bypass_regNext_31_2_df_is_ws_10;
  reg                 io_in_r_bypass_regNext_31_2_stall_10;
  reg        [15:0]   io_in_r_bypass_regNext_31_3_data_10;
  reg                 io_in_r_bypass_regNext_31_3_load_store_10;
  reg                 io_in_r_bypass_regNext_31_3_df_is_ws_10;
  reg                 io_in_r_bypass_regNext_31_3_stall_10;
  reg        [15:0]   io_in_r_bypass_regNext_0_0_data_11;
  reg                 io_in_r_bypass_regNext_0_0_load_store_11;
  reg                 io_in_r_bypass_regNext_0_0_df_is_ws_11;
  reg                 io_in_r_bypass_regNext_0_0_stall_11;
  reg        [15:0]   io_in_r_bypass_regNext_0_1_data_11;
  reg                 io_in_r_bypass_regNext_0_1_load_store_11;
  reg                 io_in_r_bypass_regNext_0_1_df_is_ws_11;
  reg                 io_in_r_bypass_regNext_0_1_stall_11;
  reg        [15:0]   io_in_r_bypass_regNext_0_2_data_11;
  reg                 io_in_r_bypass_regNext_0_2_load_store_11;
  reg                 io_in_r_bypass_regNext_0_2_df_is_ws_11;
  reg                 io_in_r_bypass_regNext_0_2_stall_11;
  reg        [15:0]   io_in_r_bypass_regNext_0_3_data_11;
  reg                 io_in_r_bypass_regNext_0_3_load_store_11;
  reg                 io_in_r_bypass_regNext_0_3_df_is_ws_11;
  reg                 io_in_r_bypass_regNext_0_3_stall_11;
  reg        [15:0]   io_in_r_bypass_regNext_1_0_data_11;
  reg                 io_in_r_bypass_regNext_1_0_load_store_11;
  reg                 io_in_r_bypass_regNext_1_0_df_is_ws_11;
  reg                 io_in_r_bypass_regNext_1_0_stall_11;
  reg        [15:0]   io_in_r_bypass_regNext_1_1_data_11;
  reg                 io_in_r_bypass_regNext_1_1_load_store_11;
  reg                 io_in_r_bypass_regNext_1_1_df_is_ws_11;
  reg                 io_in_r_bypass_regNext_1_1_stall_11;
  reg        [15:0]   io_in_r_bypass_regNext_1_2_data_11;
  reg                 io_in_r_bypass_regNext_1_2_load_store_11;
  reg                 io_in_r_bypass_regNext_1_2_df_is_ws_11;
  reg                 io_in_r_bypass_regNext_1_2_stall_11;
  reg        [15:0]   io_in_r_bypass_regNext_1_3_data_11;
  reg                 io_in_r_bypass_regNext_1_3_load_store_11;
  reg                 io_in_r_bypass_regNext_1_3_df_is_ws_11;
  reg                 io_in_r_bypass_regNext_1_3_stall_11;
  reg        [15:0]   io_in_r_bypass_regNext_2_0_data_11;
  reg                 io_in_r_bypass_regNext_2_0_load_store_11;
  reg                 io_in_r_bypass_regNext_2_0_df_is_ws_11;
  reg                 io_in_r_bypass_regNext_2_0_stall_11;
  reg        [15:0]   io_in_r_bypass_regNext_2_1_data_11;
  reg                 io_in_r_bypass_regNext_2_1_load_store_11;
  reg                 io_in_r_bypass_regNext_2_1_df_is_ws_11;
  reg                 io_in_r_bypass_regNext_2_1_stall_11;
  reg        [15:0]   io_in_r_bypass_regNext_2_2_data_11;
  reg                 io_in_r_bypass_regNext_2_2_load_store_11;
  reg                 io_in_r_bypass_regNext_2_2_df_is_ws_11;
  reg                 io_in_r_bypass_regNext_2_2_stall_11;
  reg        [15:0]   io_in_r_bypass_regNext_2_3_data_11;
  reg                 io_in_r_bypass_regNext_2_3_load_store_11;
  reg                 io_in_r_bypass_regNext_2_3_df_is_ws_11;
  reg                 io_in_r_bypass_regNext_2_3_stall_11;
  reg        [15:0]   io_in_r_bypass_regNext_3_0_data_11;
  reg                 io_in_r_bypass_regNext_3_0_load_store_11;
  reg                 io_in_r_bypass_regNext_3_0_df_is_ws_11;
  reg                 io_in_r_bypass_regNext_3_0_stall_11;
  reg        [15:0]   io_in_r_bypass_regNext_3_1_data_11;
  reg                 io_in_r_bypass_regNext_3_1_load_store_11;
  reg                 io_in_r_bypass_regNext_3_1_df_is_ws_11;
  reg                 io_in_r_bypass_regNext_3_1_stall_11;
  reg        [15:0]   io_in_r_bypass_regNext_3_2_data_11;
  reg                 io_in_r_bypass_regNext_3_2_load_store_11;
  reg                 io_in_r_bypass_regNext_3_2_df_is_ws_11;
  reg                 io_in_r_bypass_regNext_3_2_stall_11;
  reg        [15:0]   io_in_r_bypass_regNext_3_3_data_11;
  reg                 io_in_r_bypass_regNext_3_3_load_store_11;
  reg                 io_in_r_bypass_regNext_3_3_df_is_ws_11;
  reg                 io_in_r_bypass_regNext_3_3_stall_11;
  reg        [15:0]   io_in_r_bypass_regNext_4_0_data_11;
  reg                 io_in_r_bypass_regNext_4_0_load_store_11;
  reg                 io_in_r_bypass_regNext_4_0_df_is_ws_11;
  reg                 io_in_r_bypass_regNext_4_0_stall_11;
  reg        [15:0]   io_in_r_bypass_regNext_4_1_data_11;
  reg                 io_in_r_bypass_regNext_4_1_load_store_11;
  reg                 io_in_r_bypass_regNext_4_1_df_is_ws_11;
  reg                 io_in_r_bypass_regNext_4_1_stall_11;
  reg        [15:0]   io_in_r_bypass_regNext_4_2_data_11;
  reg                 io_in_r_bypass_regNext_4_2_load_store_11;
  reg                 io_in_r_bypass_regNext_4_2_df_is_ws_11;
  reg                 io_in_r_bypass_regNext_4_2_stall_11;
  reg        [15:0]   io_in_r_bypass_regNext_4_3_data_11;
  reg                 io_in_r_bypass_regNext_4_3_load_store_11;
  reg                 io_in_r_bypass_regNext_4_3_df_is_ws_11;
  reg                 io_in_r_bypass_regNext_4_3_stall_11;
  reg        [15:0]   io_in_r_bypass_regNext_5_0_data_11;
  reg                 io_in_r_bypass_regNext_5_0_load_store_11;
  reg                 io_in_r_bypass_regNext_5_0_df_is_ws_11;
  reg                 io_in_r_bypass_regNext_5_0_stall_11;
  reg        [15:0]   io_in_r_bypass_regNext_5_1_data_11;
  reg                 io_in_r_bypass_regNext_5_1_load_store_11;
  reg                 io_in_r_bypass_regNext_5_1_df_is_ws_11;
  reg                 io_in_r_bypass_regNext_5_1_stall_11;
  reg        [15:0]   io_in_r_bypass_regNext_5_2_data_11;
  reg                 io_in_r_bypass_regNext_5_2_load_store_11;
  reg                 io_in_r_bypass_regNext_5_2_df_is_ws_11;
  reg                 io_in_r_bypass_regNext_5_2_stall_11;
  reg        [15:0]   io_in_r_bypass_regNext_5_3_data_11;
  reg                 io_in_r_bypass_regNext_5_3_load_store_11;
  reg                 io_in_r_bypass_regNext_5_3_df_is_ws_11;
  reg                 io_in_r_bypass_regNext_5_3_stall_11;
  reg        [15:0]   io_in_r_bypass_regNext_6_0_data_11;
  reg                 io_in_r_bypass_regNext_6_0_load_store_11;
  reg                 io_in_r_bypass_regNext_6_0_df_is_ws_11;
  reg                 io_in_r_bypass_regNext_6_0_stall_11;
  reg        [15:0]   io_in_r_bypass_regNext_6_1_data_11;
  reg                 io_in_r_bypass_regNext_6_1_load_store_11;
  reg                 io_in_r_bypass_regNext_6_1_df_is_ws_11;
  reg                 io_in_r_bypass_regNext_6_1_stall_11;
  reg        [15:0]   io_in_r_bypass_regNext_6_2_data_11;
  reg                 io_in_r_bypass_regNext_6_2_load_store_11;
  reg                 io_in_r_bypass_regNext_6_2_df_is_ws_11;
  reg                 io_in_r_bypass_regNext_6_2_stall_11;
  reg        [15:0]   io_in_r_bypass_regNext_6_3_data_11;
  reg                 io_in_r_bypass_regNext_6_3_load_store_11;
  reg                 io_in_r_bypass_regNext_6_3_df_is_ws_11;
  reg                 io_in_r_bypass_regNext_6_3_stall_11;
  reg        [15:0]   io_in_r_bypass_regNext_7_0_data_11;
  reg                 io_in_r_bypass_regNext_7_0_load_store_11;
  reg                 io_in_r_bypass_regNext_7_0_df_is_ws_11;
  reg                 io_in_r_bypass_regNext_7_0_stall_11;
  reg        [15:0]   io_in_r_bypass_regNext_7_1_data_11;
  reg                 io_in_r_bypass_regNext_7_1_load_store_11;
  reg                 io_in_r_bypass_regNext_7_1_df_is_ws_11;
  reg                 io_in_r_bypass_regNext_7_1_stall_11;
  reg        [15:0]   io_in_r_bypass_regNext_7_2_data_11;
  reg                 io_in_r_bypass_regNext_7_2_load_store_11;
  reg                 io_in_r_bypass_regNext_7_2_df_is_ws_11;
  reg                 io_in_r_bypass_regNext_7_2_stall_11;
  reg        [15:0]   io_in_r_bypass_regNext_7_3_data_11;
  reg                 io_in_r_bypass_regNext_7_3_load_store_11;
  reg                 io_in_r_bypass_regNext_7_3_df_is_ws_11;
  reg                 io_in_r_bypass_regNext_7_3_stall_11;
  reg        [15:0]   io_in_r_bypass_regNext_8_0_data_11;
  reg                 io_in_r_bypass_regNext_8_0_load_store_11;
  reg                 io_in_r_bypass_regNext_8_0_df_is_ws_11;
  reg                 io_in_r_bypass_regNext_8_0_stall_11;
  reg        [15:0]   io_in_r_bypass_regNext_8_1_data_11;
  reg                 io_in_r_bypass_regNext_8_1_load_store_11;
  reg                 io_in_r_bypass_regNext_8_1_df_is_ws_11;
  reg                 io_in_r_bypass_regNext_8_1_stall_11;
  reg        [15:0]   io_in_r_bypass_regNext_8_2_data_11;
  reg                 io_in_r_bypass_regNext_8_2_load_store_11;
  reg                 io_in_r_bypass_regNext_8_2_df_is_ws_11;
  reg                 io_in_r_bypass_regNext_8_2_stall_11;
  reg        [15:0]   io_in_r_bypass_regNext_8_3_data_11;
  reg                 io_in_r_bypass_regNext_8_3_load_store_11;
  reg                 io_in_r_bypass_regNext_8_3_df_is_ws_11;
  reg                 io_in_r_bypass_regNext_8_3_stall_11;
  reg        [15:0]   io_in_r_bypass_regNext_9_0_data_11;
  reg                 io_in_r_bypass_regNext_9_0_load_store_11;
  reg                 io_in_r_bypass_regNext_9_0_df_is_ws_11;
  reg                 io_in_r_bypass_regNext_9_0_stall_11;
  reg        [15:0]   io_in_r_bypass_regNext_9_1_data_11;
  reg                 io_in_r_bypass_regNext_9_1_load_store_11;
  reg                 io_in_r_bypass_regNext_9_1_df_is_ws_11;
  reg                 io_in_r_bypass_regNext_9_1_stall_11;
  reg        [15:0]   io_in_r_bypass_regNext_9_2_data_11;
  reg                 io_in_r_bypass_regNext_9_2_load_store_11;
  reg                 io_in_r_bypass_regNext_9_2_df_is_ws_11;
  reg                 io_in_r_bypass_regNext_9_2_stall_11;
  reg        [15:0]   io_in_r_bypass_regNext_9_3_data_11;
  reg                 io_in_r_bypass_regNext_9_3_load_store_11;
  reg                 io_in_r_bypass_regNext_9_3_df_is_ws_11;
  reg                 io_in_r_bypass_regNext_9_3_stall_11;
  reg        [15:0]   io_in_r_bypass_regNext_10_0_data_11;
  reg                 io_in_r_bypass_regNext_10_0_load_store_11;
  reg                 io_in_r_bypass_regNext_10_0_df_is_ws_11;
  reg                 io_in_r_bypass_regNext_10_0_stall_11;
  reg        [15:0]   io_in_r_bypass_regNext_10_1_data_11;
  reg                 io_in_r_bypass_regNext_10_1_load_store_11;
  reg                 io_in_r_bypass_regNext_10_1_df_is_ws_11;
  reg                 io_in_r_bypass_regNext_10_1_stall_11;
  reg        [15:0]   io_in_r_bypass_regNext_10_2_data_11;
  reg                 io_in_r_bypass_regNext_10_2_load_store_11;
  reg                 io_in_r_bypass_regNext_10_2_df_is_ws_11;
  reg                 io_in_r_bypass_regNext_10_2_stall_11;
  reg        [15:0]   io_in_r_bypass_regNext_10_3_data_11;
  reg                 io_in_r_bypass_regNext_10_3_load_store_11;
  reg                 io_in_r_bypass_regNext_10_3_df_is_ws_11;
  reg                 io_in_r_bypass_regNext_10_3_stall_11;
  reg        [15:0]   io_in_r_bypass_regNext_11_0_data_11;
  reg                 io_in_r_bypass_regNext_11_0_load_store_11;
  reg                 io_in_r_bypass_regNext_11_0_df_is_ws_11;
  reg                 io_in_r_bypass_regNext_11_0_stall_11;
  reg        [15:0]   io_in_r_bypass_regNext_11_1_data_11;
  reg                 io_in_r_bypass_regNext_11_1_load_store_11;
  reg                 io_in_r_bypass_regNext_11_1_df_is_ws_11;
  reg                 io_in_r_bypass_regNext_11_1_stall_11;
  reg        [15:0]   io_in_r_bypass_regNext_11_2_data_11;
  reg                 io_in_r_bypass_regNext_11_2_load_store_11;
  reg                 io_in_r_bypass_regNext_11_2_df_is_ws_11;
  reg                 io_in_r_bypass_regNext_11_2_stall_11;
  reg        [15:0]   io_in_r_bypass_regNext_11_3_data_11;
  reg                 io_in_r_bypass_regNext_11_3_load_store_11;
  reg                 io_in_r_bypass_regNext_11_3_df_is_ws_11;
  reg                 io_in_r_bypass_regNext_11_3_stall_11;
  reg        [15:0]   io_in_r_bypass_regNext_12_0_data_11;
  reg                 io_in_r_bypass_regNext_12_0_load_store_11;
  reg                 io_in_r_bypass_regNext_12_0_df_is_ws_11;
  reg                 io_in_r_bypass_regNext_12_0_stall_11;
  reg        [15:0]   io_in_r_bypass_regNext_12_1_data_11;
  reg                 io_in_r_bypass_regNext_12_1_load_store_11;
  reg                 io_in_r_bypass_regNext_12_1_df_is_ws_11;
  reg                 io_in_r_bypass_regNext_12_1_stall_11;
  reg        [15:0]   io_in_r_bypass_regNext_12_2_data_11;
  reg                 io_in_r_bypass_regNext_12_2_load_store_11;
  reg                 io_in_r_bypass_regNext_12_2_df_is_ws_11;
  reg                 io_in_r_bypass_regNext_12_2_stall_11;
  reg        [15:0]   io_in_r_bypass_regNext_12_3_data_11;
  reg                 io_in_r_bypass_regNext_12_3_load_store_11;
  reg                 io_in_r_bypass_regNext_12_3_df_is_ws_11;
  reg                 io_in_r_bypass_regNext_12_3_stall_11;
  reg        [15:0]   io_in_r_bypass_regNext_13_0_data_11;
  reg                 io_in_r_bypass_regNext_13_0_load_store_11;
  reg                 io_in_r_bypass_regNext_13_0_df_is_ws_11;
  reg                 io_in_r_bypass_regNext_13_0_stall_11;
  reg        [15:0]   io_in_r_bypass_regNext_13_1_data_11;
  reg                 io_in_r_bypass_regNext_13_1_load_store_11;
  reg                 io_in_r_bypass_regNext_13_1_df_is_ws_11;
  reg                 io_in_r_bypass_regNext_13_1_stall_11;
  reg        [15:0]   io_in_r_bypass_regNext_13_2_data_11;
  reg                 io_in_r_bypass_regNext_13_2_load_store_11;
  reg                 io_in_r_bypass_regNext_13_2_df_is_ws_11;
  reg                 io_in_r_bypass_regNext_13_2_stall_11;
  reg        [15:0]   io_in_r_bypass_regNext_13_3_data_11;
  reg                 io_in_r_bypass_regNext_13_3_load_store_11;
  reg                 io_in_r_bypass_regNext_13_3_df_is_ws_11;
  reg                 io_in_r_bypass_regNext_13_3_stall_11;
  reg        [15:0]   io_in_r_bypass_regNext_14_0_data_11;
  reg                 io_in_r_bypass_regNext_14_0_load_store_11;
  reg                 io_in_r_bypass_regNext_14_0_df_is_ws_11;
  reg                 io_in_r_bypass_regNext_14_0_stall_11;
  reg        [15:0]   io_in_r_bypass_regNext_14_1_data_11;
  reg                 io_in_r_bypass_regNext_14_1_load_store_11;
  reg                 io_in_r_bypass_regNext_14_1_df_is_ws_11;
  reg                 io_in_r_bypass_regNext_14_1_stall_11;
  reg        [15:0]   io_in_r_bypass_regNext_14_2_data_11;
  reg                 io_in_r_bypass_regNext_14_2_load_store_11;
  reg                 io_in_r_bypass_regNext_14_2_df_is_ws_11;
  reg                 io_in_r_bypass_regNext_14_2_stall_11;
  reg        [15:0]   io_in_r_bypass_regNext_14_3_data_11;
  reg                 io_in_r_bypass_regNext_14_3_load_store_11;
  reg                 io_in_r_bypass_regNext_14_3_df_is_ws_11;
  reg                 io_in_r_bypass_regNext_14_3_stall_11;
  reg        [15:0]   io_in_r_bypass_regNext_15_0_data_11;
  reg                 io_in_r_bypass_regNext_15_0_load_store_11;
  reg                 io_in_r_bypass_regNext_15_0_df_is_ws_11;
  reg                 io_in_r_bypass_regNext_15_0_stall_11;
  reg        [15:0]   io_in_r_bypass_regNext_15_1_data_11;
  reg                 io_in_r_bypass_regNext_15_1_load_store_11;
  reg                 io_in_r_bypass_regNext_15_1_df_is_ws_11;
  reg                 io_in_r_bypass_regNext_15_1_stall_11;
  reg        [15:0]   io_in_r_bypass_regNext_15_2_data_11;
  reg                 io_in_r_bypass_regNext_15_2_load_store_11;
  reg                 io_in_r_bypass_regNext_15_2_df_is_ws_11;
  reg                 io_in_r_bypass_regNext_15_2_stall_11;
  reg        [15:0]   io_in_r_bypass_regNext_15_3_data_11;
  reg                 io_in_r_bypass_regNext_15_3_load_store_11;
  reg                 io_in_r_bypass_regNext_15_3_df_is_ws_11;
  reg                 io_in_r_bypass_regNext_15_3_stall_11;
  reg        [15:0]   io_in_r_bypass_regNext_16_0_data_11;
  reg                 io_in_r_bypass_regNext_16_0_load_store_11;
  reg                 io_in_r_bypass_regNext_16_0_df_is_ws_11;
  reg                 io_in_r_bypass_regNext_16_0_stall_11;
  reg        [15:0]   io_in_r_bypass_regNext_16_1_data_11;
  reg                 io_in_r_bypass_regNext_16_1_load_store_11;
  reg                 io_in_r_bypass_regNext_16_1_df_is_ws_11;
  reg                 io_in_r_bypass_regNext_16_1_stall_11;
  reg        [15:0]   io_in_r_bypass_regNext_16_2_data_11;
  reg                 io_in_r_bypass_regNext_16_2_load_store_11;
  reg                 io_in_r_bypass_regNext_16_2_df_is_ws_11;
  reg                 io_in_r_bypass_regNext_16_2_stall_11;
  reg        [15:0]   io_in_r_bypass_regNext_16_3_data_11;
  reg                 io_in_r_bypass_regNext_16_3_load_store_11;
  reg                 io_in_r_bypass_regNext_16_3_df_is_ws_11;
  reg                 io_in_r_bypass_regNext_16_3_stall_11;
  reg        [15:0]   io_in_r_bypass_regNext_17_0_data_11;
  reg                 io_in_r_bypass_regNext_17_0_load_store_11;
  reg                 io_in_r_bypass_regNext_17_0_df_is_ws_11;
  reg                 io_in_r_bypass_regNext_17_0_stall_11;
  reg        [15:0]   io_in_r_bypass_regNext_17_1_data_11;
  reg                 io_in_r_bypass_regNext_17_1_load_store_11;
  reg                 io_in_r_bypass_regNext_17_1_df_is_ws_11;
  reg                 io_in_r_bypass_regNext_17_1_stall_11;
  reg        [15:0]   io_in_r_bypass_regNext_17_2_data_11;
  reg                 io_in_r_bypass_regNext_17_2_load_store_11;
  reg                 io_in_r_bypass_regNext_17_2_df_is_ws_11;
  reg                 io_in_r_bypass_regNext_17_2_stall_11;
  reg        [15:0]   io_in_r_bypass_regNext_17_3_data_11;
  reg                 io_in_r_bypass_regNext_17_3_load_store_11;
  reg                 io_in_r_bypass_regNext_17_3_df_is_ws_11;
  reg                 io_in_r_bypass_regNext_17_3_stall_11;
  reg        [15:0]   io_in_r_bypass_regNext_18_0_data_11;
  reg                 io_in_r_bypass_regNext_18_0_load_store_11;
  reg                 io_in_r_bypass_regNext_18_0_df_is_ws_11;
  reg                 io_in_r_bypass_regNext_18_0_stall_11;
  reg        [15:0]   io_in_r_bypass_regNext_18_1_data_11;
  reg                 io_in_r_bypass_regNext_18_1_load_store_11;
  reg                 io_in_r_bypass_regNext_18_1_df_is_ws_11;
  reg                 io_in_r_bypass_regNext_18_1_stall_11;
  reg        [15:0]   io_in_r_bypass_regNext_18_2_data_11;
  reg                 io_in_r_bypass_regNext_18_2_load_store_11;
  reg                 io_in_r_bypass_regNext_18_2_df_is_ws_11;
  reg                 io_in_r_bypass_regNext_18_2_stall_11;
  reg        [15:0]   io_in_r_bypass_regNext_18_3_data_11;
  reg                 io_in_r_bypass_regNext_18_3_load_store_11;
  reg                 io_in_r_bypass_regNext_18_3_df_is_ws_11;
  reg                 io_in_r_bypass_regNext_18_3_stall_11;
  reg        [15:0]   io_in_r_bypass_regNext_19_0_data_11;
  reg                 io_in_r_bypass_regNext_19_0_load_store_11;
  reg                 io_in_r_bypass_regNext_19_0_df_is_ws_11;
  reg                 io_in_r_bypass_regNext_19_0_stall_11;
  reg        [15:0]   io_in_r_bypass_regNext_19_1_data_11;
  reg                 io_in_r_bypass_regNext_19_1_load_store_11;
  reg                 io_in_r_bypass_regNext_19_1_df_is_ws_11;
  reg                 io_in_r_bypass_regNext_19_1_stall_11;
  reg        [15:0]   io_in_r_bypass_regNext_19_2_data_11;
  reg                 io_in_r_bypass_regNext_19_2_load_store_11;
  reg                 io_in_r_bypass_regNext_19_2_df_is_ws_11;
  reg                 io_in_r_bypass_regNext_19_2_stall_11;
  reg        [15:0]   io_in_r_bypass_regNext_19_3_data_11;
  reg                 io_in_r_bypass_regNext_19_3_load_store_11;
  reg                 io_in_r_bypass_regNext_19_3_df_is_ws_11;
  reg                 io_in_r_bypass_regNext_19_3_stall_11;
  reg        [15:0]   io_in_r_bypass_regNext_20_0_data_11;
  reg                 io_in_r_bypass_regNext_20_0_load_store_11;
  reg                 io_in_r_bypass_regNext_20_0_df_is_ws_11;
  reg                 io_in_r_bypass_regNext_20_0_stall_11;
  reg        [15:0]   io_in_r_bypass_regNext_20_1_data_11;
  reg                 io_in_r_bypass_regNext_20_1_load_store_11;
  reg                 io_in_r_bypass_regNext_20_1_df_is_ws_11;
  reg                 io_in_r_bypass_regNext_20_1_stall_11;
  reg        [15:0]   io_in_r_bypass_regNext_20_2_data_11;
  reg                 io_in_r_bypass_regNext_20_2_load_store_11;
  reg                 io_in_r_bypass_regNext_20_2_df_is_ws_11;
  reg                 io_in_r_bypass_regNext_20_2_stall_11;
  reg        [15:0]   io_in_r_bypass_regNext_20_3_data_11;
  reg                 io_in_r_bypass_regNext_20_3_load_store_11;
  reg                 io_in_r_bypass_regNext_20_3_df_is_ws_11;
  reg                 io_in_r_bypass_regNext_20_3_stall_11;
  reg        [15:0]   io_in_r_bypass_regNext_21_0_data_11;
  reg                 io_in_r_bypass_regNext_21_0_load_store_11;
  reg                 io_in_r_bypass_regNext_21_0_df_is_ws_11;
  reg                 io_in_r_bypass_regNext_21_0_stall_11;
  reg        [15:0]   io_in_r_bypass_regNext_21_1_data_11;
  reg                 io_in_r_bypass_regNext_21_1_load_store_11;
  reg                 io_in_r_bypass_regNext_21_1_df_is_ws_11;
  reg                 io_in_r_bypass_regNext_21_1_stall_11;
  reg        [15:0]   io_in_r_bypass_regNext_21_2_data_11;
  reg                 io_in_r_bypass_regNext_21_2_load_store_11;
  reg                 io_in_r_bypass_regNext_21_2_df_is_ws_11;
  reg                 io_in_r_bypass_regNext_21_2_stall_11;
  reg        [15:0]   io_in_r_bypass_regNext_21_3_data_11;
  reg                 io_in_r_bypass_regNext_21_3_load_store_11;
  reg                 io_in_r_bypass_regNext_21_3_df_is_ws_11;
  reg                 io_in_r_bypass_regNext_21_3_stall_11;
  reg        [15:0]   io_in_r_bypass_regNext_22_0_data_11;
  reg                 io_in_r_bypass_regNext_22_0_load_store_11;
  reg                 io_in_r_bypass_regNext_22_0_df_is_ws_11;
  reg                 io_in_r_bypass_regNext_22_0_stall_11;
  reg        [15:0]   io_in_r_bypass_regNext_22_1_data_11;
  reg                 io_in_r_bypass_regNext_22_1_load_store_11;
  reg                 io_in_r_bypass_regNext_22_1_df_is_ws_11;
  reg                 io_in_r_bypass_regNext_22_1_stall_11;
  reg        [15:0]   io_in_r_bypass_regNext_22_2_data_11;
  reg                 io_in_r_bypass_regNext_22_2_load_store_11;
  reg                 io_in_r_bypass_regNext_22_2_df_is_ws_11;
  reg                 io_in_r_bypass_regNext_22_2_stall_11;
  reg        [15:0]   io_in_r_bypass_regNext_22_3_data_11;
  reg                 io_in_r_bypass_regNext_22_3_load_store_11;
  reg                 io_in_r_bypass_regNext_22_3_df_is_ws_11;
  reg                 io_in_r_bypass_regNext_22_3_stall_11;
  reg        [15:0]   io_in_r_bypass_regNext_23_0_data_11;
  reg                 io_in_r_bypass_regNext_23_0_load_store_11;
  reg                 io_in_r_bypass_regNext_23_0_df_is_ws_11;
  reg                 io_in_r_bypass_regNext_23_0_stall_11;
  reg        [15:0]   io_in_r_bypass_regNext_23_1_data_11;
  reg                 io_in_r_bypass_regNext_23_1_load_store_11;
  reg                 io_in_r_bypass_regNext_23_1_df_is_ws_11;
  reg                 io_in_r_bypass_regNext_23_1_stall_11;
  reg        [15:0]   io_in_r_bypass_regNext_23_2_data_11;
  reg                 io_in_r_bypass_regNext_23_2_load_store_11;
  reg                 io_in_r_bypass_regNext_23_2_df_is_ws_11;
  reg                 io_in_r_bypass_regNext_23_2_stall_11;
  reg        [15:0]   io_in_r_bypass_regNext_23_3_data_11;
  reg                 io_in_r_bypass_regNext_23_3_load_store_11;
  reg                 io_in_r_bypass_regNext_23_3_df_is_ws_11;
  reg                 io_in_r_bypass_regNext_23_3_stall_11;
  reg        [15:0]   io_in_r_bypass_regNext_24_0_data_11;
  reg                 io_in_r_bypass_regNext_24_0_load_store_11;
  reg                 io_in_r_bypass_regNext_24_0_df_is_ws_11;
  reg                 io_in_r_bypass_regNext_24_0_stall_11;
  reg        [15:0]   io_in_r_bypass_regNext_24_1_data_11;
  reg                 io_in_r_bypass_regNext_24_1_load_store_11;
  reg                 io_in_r_bypass_regNext_24_1_df_is_ws_11;
  reg                 io_in_r_bypass_regNext_24_1_stall_11;
  reg        [15:0]   io_in_r_bypass_regNext_24_2_data_11;
  reg                 io_in_r_bypass_regNext_24_2_load_store_11;
  reg                 io_in_r_bypass_regNext_24_2_df_is_ws_11;
  reg                 io_in_r_bypass_regNext_24_2_stall_11;
  reg        [15:0]   io_in_r_bypass_regNext_24_3_data_11;
  reg                 io_in_r_bypass_regNext_24_3_load_store_11;
  reg                 io_in_r_bypass_regNext_24_3_df_is_ws_11;
  reg                 io_in_r_bypass_regNext_24_3_stall_11;
  reg        [15:0]   io_in_r_bypass_regNext_25_0_data_11;
  reg                 io_in_r_bypass_regNext_25_0_load_store_11;
  reg                 io_in_r_bypass_regNext_25_0_df_is_ws_11;
  reg                 io_in_r_bypass_regNext_25_0_stall_11;
  reg        [15:0]   io_in_r_bypass_regNext_25_1_data_11;
  reg                 io_in_r_bypass_regNext_25_1_load_store_11;
  reg                 io_in_r_bypass_regNext_25_1_df_is_ws_11;
  reg                 io_in_r_bypass_regNext_25_1_stall_11;
  reg        [15:0]   io_in_r_bypass_regNext_25_2_data_11;
  reg                 io_in_r_bypass_regNext_25_2_load_store_11;
  reg                 io_in_r_bypass_regNext_25_2_df_is_ws_11;
  reg                 io_in_r_bypass_regNext_25_2_stall_11;
  reg        [15:0]   io_in_r_bypass_regNext_25_3_data_11;
  reg                 io_in_r_bypass_regNext_25_3_load_store_11;
  reg                 io_in_r_bypass_regNext_25_3_df_is_ws_11;
  reg                 io_in_r_bypass_regNext_25_3_stall_11;
  reg        [15:0]   io_in_r_bypass_regNext_26_0_data_11;
  reg                 io_in_r_bypass_regNext_26_0_load_store_11;
  reg                 io_in_r_bypass_regNext_26_0_df_is_ws_11;
  reg                 io_in_r_bypass_regNext_26_0_stall_11;
  reg        [15:0]   io_in_r_bypass_regNext_26_1_data_11;
  reg                 io_in_r_bypass_regNext_26_1_load_store_11;
  reg                 io_in_r_bypass_regNext_26_1_df_is_ws_11;
  reg                 io_in_r_bypass_regNext_26_1_stall_11;
  reg        [15:0]   io_in_r_bypass_regNext_26_2_data_11;
  reg                 io_in_r_bypass_regNext_26_2_load_store_11;
  reg                 io_in_r_bypass_regNext_26_2_df_is_ws_11;
  reg                 io_in_r_bypass_regNext_26_2_stall_11;
  reg        [15:0]   io_in_r_bypass_regNext_26_3_data_11;
  reg                 io_in_r_bypass_regNext_26_3_load_store_11;
  reg                 io_in_r_bypass_regNext_26_3_df_is_ws_11;
  reg                 io_in_r_bypass_regNext_26_3_stall_11;
  reg        [15:0]   io_in_r_bypass_regNext_27_0_data_11;
  reg                 io_in_r_bypass_regNext_27_0_load_store_11;
  reg                 io_in_r_bypass_regNext_27_0_df_is_ws_11;
  reg                 io_in_r_bypass_regNext_27_0_stall_11;
  reg        [15:0]   io_in_r_bypass_regNext_27_1_data_11;
  reg                 io_in_r_bypass_regNext_27_1_load_store_11;
  reg                 io_in_r_bypass_regNext_27_1_df_is_ws_11;
  reg                 io_in_r_bypass_regNext_27_1_stall_11;
  reg        [15:0]   io_in_r_bypass_regNext_27_2_data_11;
  reg                 io_in_r_bypass_regNext_27_2_load_store_11;
  reg                 io_in_r_bypass_regNext_27_2_df_is_ws_11;
  reg                 io_in_r_bypass_regNext_27_2_stall_11;
  reg        [15:0]   io_in_r_bypass_regNext_27_3_data_11;
  reg                 io_in_r_bypass_regNext_27_3_load_store_11;
  reg                 io_in_r_bypass_regNext_27_3_df_is_ws_11;
  reg                 io_in_r_bypass_regNext_27_3_stall_11;
  reg        [15:0]   io_in_r_bypass_regNext_28_0_data_11;
  reg                 io_in_r_bypass_regNext_28_0_load_store_11;
  reg                 io_in_r_bypass_regNext_28_0_df_is_ws_11;
  reg                 io_in_r_bypass_regNext_28_0_stall_11;
  reg        [15:0]   io_in_r_bypass_regNext_28_1_data_11;
  reg                 io_in_r_bypass_regNext_28_1_load_store_11;
  reg                 io_in_r_bypass_regNext_28_1_df_is_ws_11;
  reg                 io_in_r_bypass_regNext_28_1_stall_11;
  reg        [15:0]   io_in_r_bypass_regNext_28_2_data_11;
  reg                 io_in_r_bypass_regNext_28_2_load_store_11;
  reg                 io_in_r_bypass_regNext_28_2_df_is_ws_11;
  reg                 io_in_r_bypass_regNext_28_2_stall_11;
  reg        [15:0]   io_in_r_bypass_regNext_28_3_data_11;
  reg                 io_in_r_bypass_regNext_28_3_load_store_11;
  reg                 io_in_r_bypass_regNext_28_3_df_is_ws_11;
  reg                 io_in_r_bypass_regNext_28_3_stall_11;
  reg        [15:0]   io_in_r_bypass_regNext_29_0_data_11;
  reg                 io_in_r_bypass_regNext_29_0_load_store_11;
  reg                 io_in_r_bypass_regNext_29_0_df_is_ws_11;
  reg                 io_in_r_bypass_regNext_29_0_stall_11;
  reg        [15:0]   io_in_r_bypass_regNext_29_1_data_11;
  reg                 io_in_r_bypass_regNext_29_1_load_store_11;
  reg                 io_in_r_bypass_regNext_29_1_df_is_ws_11;
  reg                 io_in_r_bypass_regNext_29_1_stall_11;
  reg        [15:0]   io_in_r_bypass_regNext_29_2_data_11;
  reg                 io_in_r_bypass_regNext_29_2_load_store_11;
  reg                 io_in_r_bypass_regNext_29_2_df_is_ws_11;
  reg                 io_in_r_bypass_regNext_29_2_stall_11;
  reg        [15:0]   io_in_r_bypass_regNext_29_3_data_11;
  reg                 io_in_r_bypass_regNext_29_3_load_store_11;
  reg                 io_in_r_bypass_regNext_29_3_df_is_ws_11;
  reg                 io_in_r_bypass_regNext_29_3_stall_11;
  reg        [15:0]   io_in_r_bypass_regNext_30_0_data_11;
  reg                 io_in_r_bypass_regNext_30_0_load_store_11;
  reg                 io_in_r_bypass_regNext_30_0_df_is_ws_11;
  reg                 io_in_r_bypass_regNext_30_0_stall_11;
  reg        [15:0]   io_in_r_bypass_regNext_30_1_data_11;
  reg                 io_in_r_bypass_regNext_30_1_load_store_11;
  reg                 io_in_r_bypass_regNext_30_1_df_is_ws_11;
  reg                 io_in_r_bypass_regNext_30_1_stall_11;
  reg        [15:0]   io_in_r_bypass_regNext_30_2_data_11;
  reg                 io_in_r_bypass_regNext_30_2_load_store_11;
  reg                 io_in_r_bypass_regNext_30_2_df_is_ws_11;
  reg                 io_in_r_bypass_regNext_30_2_stall_11;
  reg        [15:0]   io_in_r_bypass_regNext_30_3_data_11;
  reg                 io_in_r_bypass_regNext_30_3_load_store_11;
  reg                 io_in_r_bypass_regNext_30_3_df_is_ws_11;
  reg                 io_in_r_bypass_regNext_30_3_stall_11;
  reg        [15:0]   io_in_r_bypass_regNext_31_0_data_11;
  reg                 io_in_r_bypass_regNext_31_0_load_store_11;
  reg                 io_in_r_bypass_regNext_31_0_df_is_ws_11;
  reg                 io_in_r_bypass_regNext_31_0_stall_11;
  reg        [15:0]   io_in_r_bypass_regNext_31_1_data_11;
  reg                 io_in_r_bypass_regNext_31_1_load_store_11;
  reg                 io_in_r_bypass_regNext_31_1_df_is_ws_11;
  reg                 io_in_r_bypass_regNext_31_1_stall_11;
  reg        [15:0]   io_in_r_bypass_regNext_31_2_data_11;
  reg                 io_in_r_bypass_regNext_31_2_load_store_11;
  reg                 io_in_r_bypass_regNext_31_2_df_is_ws_11;
  reg                 io_in_r_bypass_regNext_31_2_stall_11;
  reg        [15:0]   io_in_r_bypass_regNext_31_3_data_11;
  reg                 io_in_r_bypass_regNext_31_3_load_store_11;
  reg                 io_in_r_bypass_regNext_31_3_df_is_ws_11;
  reg                 io_in_r_bypass_regNext_31_3_stall_11;
  reg        [15:0]   io_in_r_bypass_regNext_0_0_data_12;
  reg                 io_in_r_bypass_regNext_0_0_load_store_12;
  reg                 io_in_r_bypass_regNext_0_0_df_is_ws_12;
  reg                 io_in_r_bypass_regNext_0_0_stall_12;
  reg        [15:0]   io_in_r_bypass_regNext_0_1_data_12;
  reg                 io_in_r_bypass_regNext_0_1_load_store_12;
  reg                 io_in_r_bypass_regNext_0_1_df_is_ws_12;
  reg                 io_in_r_bypass_regNext_0_1_stall_12;
  reg        [15:0]   io_in_r_bypass_regNext_0_2_data_12;
  reg                 io_in_r_bypass_regNext_0_2_load_store_12;
  reg                 io_in_r_bypass_regNext_0_2_df_is_ws_12;
  reg                 io_in_r_bypass_regNext_0_2_stall_12;
  reg        [15:0]   io_in_r_bypass_regNext_0_3_data_12;
  reg                 io_in_r_bypass_regNext_0_3_load_store_12;
  reg                 io_in_r_bypass_regNext_0_3_df_is_ws_12;
  reg                 io_in_r_bypass_regNext_0_3_stall_12;
  reg        [15:0]   io_in_r_bypass_regNext_1_0_data_12;
  reg                 io_in_r_bypass_regNext_1_0_load_store_12;
  reg                 io_in_r_bypass_regNext_1_0_df_is_ws_12;
  reg                 io_in_r_bypass_regNext_1_0_stall_12;
  reg        [15:0]   io_in_r_bypass_regNext_1_1_data_12;
  reg                 io_in_r_bypass_regNext_1_1_load_store_12;
  reg                 io_in_r_bypass_regNext_1_1_df_is_ws_12;
  reg                 io_in_r_bypass_regNext_1_1_stall_12;
  reg        [15:0]   io_in_r_bypass_regNext_1_2_data_12;
  reg                 io_in_r_bypass_regNext_1_2_load_store_12;
  reg                 io_in_r_bypass_regNext_1_2_df_is_ws_12;
  reg                 io_in_r_bypass_regNext_1_2_stall_12;
  reg        [15:0]   io_in_r_bypass_regNext_1_3_data_12;
  reg                 io_in_r_bypass_regNext_1_3_load_store_12;
  reg                 io_in_r_bypass_regNext_1_3_df_is_ws_12;
  reg                 io_in_r_bypass_regNext_1_3_stall_12;
  reg        [15:0]   io_in_r_bypass_regNext_2_0_data_12;
  reg                 io_in_r_bypass_regNext_2_0_load_store_12;
  reg                 io_in_r_bypass_regNext_2_0_df_is_ws_12;
  reg                 io_in_r_bypass_regNext_2_0_stall_12;
  reg        [15:0]   io_in_r_bypass_regNext_2_1_data_12;
  reg                 io_in_r_bypass_regNext_2_1_load_store_12;
  reg                 io_in_r_bypass_regNext_2_1_df_is_ws_12;
  reg                 io_in_r_bypass_regNext_2_1_stall_12;
  reg        [15:0]   io_in_r_bypass_regNext_2_2_data_12;
  reg                 io_in_r_bypass_regNext_2_2_load_store_12;
  reg                 io_in_r_bypass_regNext_2_2_df_is_ws_12;
  reg                 io_in_r_bypass_regNext_2_2_stall_12;
  reg        [15:0]   io_in_r_bypass_regNext_2_3_data_12;
  reg                 io_in_r_bypass_regNext_2_3_load_store_12;
  reg                 io_in_r_bypass_regNext_2_3_df_is_ws_12;
  reg                 io_in_r_bypass_regNext_2_3_stall_12;
  reg        [15:0]   io_in_r_bypass_regNext_3_0_data_12;
  reg                 io_in_r_bypass_regNext_3_0_load_store_12;
  reg                 io_in_r_bypass_regNext_3_0_df_is_ws_12;
  reg                 io_in_r_bypass_regNext_3_0_stall_12;
  reg        [15:0]   io_in_r_bypass_regNext_3_1_data_12;
  reg                 io_in_r_bypass_regNext_3_1_load_store_12;
  reg                 io_in_r_bypass_regNext_3_1_df_is_ws_12;
  reg                 io_in_r_bypass_regNext_3_1_stall_12;
  reg        [15:0]   io_in_r_bypass_regNext_3_2_data_12;
  reg                 io_in_r_bypass_regNext_3_2_load_store_12;
  reg                 io_in_r_bypass_regNext_3_2_df_is_ws_12;
  reg                 io_in_r_bypass_regNext_3_2_stall_12;
  reg        [15:0]   io_in_r_bypass_regNext_3_3_data_12;
  reg                 io_in_r_bypass_regNext_3_3_load_store_12;
  reg                 io_in_r_bypass_regNext_3_3_df_is_ws_12;
  reg                 io_in_r_bypass_regNext_3_3_stall_12;
  reg        [15:0]   io_in_r_bypass_regNext_4_0_data_12;
  reg                 io_in_r_bypass_regNext_4_0_load_store_12;
  reg                 io_in_r_bypass_regNext_4_0_df_is_ws_12;
  reg                 io_in_r_bypass_regNext_4_0_stall_12;
  reg        [15:0]   io_in_r_bypass_regNext_4_1_data_12;
  reg                 io_in_r_bypass_regNext_4_1_load_store_12;
  reg                 io_in_r_bypass_regNext_4_1_df_is_ws_12;
  reg                 io_in_r_bypass_regNext_4_1_stall_12;
  reg        [15:0]   io_in_r_bypass_regNext_4_2_data_12;
  reg                 io_in_r_bypass_regNext_4_2_load_store_12;
  reg                 io_in_r_bypass_regNext_4_2_df_is_ws_12;
  reg                 io_in_r_bypass_regNext_4_2_stall_12;
  reg        [15:0]   io_in_r_bypass_regNext_4_3_data_12;
  reg                 io_in_r_bypass_regNext_4_3_load_store_12;
  reg                 io_in_r_bypass_regNext_4_3_df_is_ws_12;
  reg                 io_in_r_bypass_regNext_4_3_stall_12;
  reg        [15:0]   io_in_r_bypass_regNext_5_0_data_12;
  reg                 io_in_r_bypass_regNext_5_0_load_store_12;
  reg                 io_in_r_bypass_regNext_5_0_df_is_ws_12;
  reg                 io_in_r_bypass_regNext_5_0_stall_12;
  reg        [15:0]   io_in_r_bypass_regNext_5_1_data_12;
  reg                 io_in_r_bypass_regNext_5_1_load_store_12;
  reg                 io_in_r_bypass_regNext_5_1_df_is_ws_12;
  reg                 io_in_r_bypass_regNext_5_1_stall_12;
  reg        [15:0]   io_in_r_bypass_regNext_5_2_data_12;
  reg                 io_in_r_bypass_regNext_5_2_load_store_12;
  reg                 io_in_r_bypass_regNext_5_2_df_is_ws_12;
  reg                 io_in_r_bypass_regNext_5_2_stall_12;
  reg        [15:0]   io_in_r_bypass_regNext_5_3_data_12;
  reg                 io_in_r_bypass_regNext_5_3_load_store_12;
  reg                 io_in_r_bypass_regNext_5_3_df_is_ws_12;
  reg                 io_in_r_bypass_regNext_5_3_stall_12;
  reg        [15:0]   io_in_r_bypass_regNext_6_0_data_12;
  reg                 io_in_r_bypass_regNext_6_0_load_store_12;
  reg                 io_in_r_bypass_regNext_6_0_df_is_ws_12;
  reg                 io_in_r_bypass_regNext_6_0_stall_12;
  reg        [15:0]   io_in_r_bypass_regNext_6_1_data_12;
  reg                 io_in_r_bypass_regNext_6_1_load_store_12;
  reg                 io_in_r_bypass_regNext_6_1_df_is_ws_12;
  reg                 io_in_r_bypass_regNext_6_1_stall_12;
  reg        [15:0]   io_in_r_bypass_regNext_6_2_data_12;
  reg                 io_in_r_bypass_regNext_6_2_load_store_12;
  reg                 io_in_r_bypass_regNext_6_2_df_is_ws_12;
  reg                 io_in_r_bypass_regNext_6_2_stall_12;
  reg        [15:0]   io_in_r_bypass_regNext_6_3_data_12;
  reg                 io_in_r_bypass_regNext_6_3_load_store_12;
  reg                 io_in_r_bypass_regNext_6_3_df_is_ws_12;
  reg                 io_in_r_bypass_regNext_6_3_stall_12;
  reg        [15:0]   io_in_r_bypass_regNext_7_0_data_12;
  reg                 io_in_r_bypass_regNext_7_0_load_store_12;
  reg                 io_in_r_bypass_regNext_7_0_df_is_ws_12;
  reg                 io_in_r_bypass_regNext_7_0_stall_12;
  reg        [15:0]   io_in_r_bypass_regNext_7_1_data_12;
  reg                 io_in_r_bypass_regNext_7_1_load_store_12;
  reg                 io_in_r_bypass_regNext_7_1_df_is_ws_12;
  reg                 io_in_r_bypass_regNext_7_1_stall_12;
  reg        [15:0]   io_in_r_bypass_regNext_7_2_data_12;
  reg                 io_in_r_bypass_regNext_7_2_load_store_12;
  reg                 io_in_r_bypass_regNext_7_2_df_is_ws_12;
  reg                 io_in_r_bypass_regNext_7_2_stall_12;
  reg        [15:0]   io_in_r_bypass_regNext_7_3_data_12;
  reg                 io_in_r_bypass_regNext_7_3_load_store_12;
  reg                 io_in_r_bypass_regNext_7_3_df_is_ws_12;
  reg                 io_in_r_bypass_regNext_7_3_stall_12;
  reg        [15:0]   io_in_r_bypass_regNext_8_0_data_12;
  reg                 io_in_r_bypass_regNext_8_0_load_store_12;
  reg                 io_in_r_bypass_regNext_8_0_df_is_ws_12;
  reg                 io_in_r_bypass_regNext_8_0_stall_12;
  reg        [15:0]   io_in_r_bypass_regNext_8_1_data_12;
  reg                 io_in_r_bypass_regNext_8_1_load_store_12;
  reg                 io_in_r_bypass_regNext_8_1_df_is_ws_12;
  reg                 io_in_r_bypass_regNext_8_1_stall_12;
  reg        [15:0]   io_in_r_bypass_regNext_8_2_data_12;
  reg                 io_in_r_bypass_regNext_8_2_load_store_12;
  reg                 io_in_r_bypass_regNext_8_2_df_is_ws_12;
  reg                 io_in_r_bypass_regNext_8_2_stall_12;
  reg        [15:0]   io_in_r_bypass_regNext_8_3_data_12;
  reg                 io_in_r_bypass_regNext_8_3_load_store_12;
  reg                 io_in_r_bypass_regNext_8_3_df_is_ws_12;
  reg                 io_in_r_bypass_regNext_8_3_stall_12;
  reg        [15:0]   io_in_r_bypass_regNext_9_0_data_12;
  reg                 io_in_r_bypass_regNext_9_0_load_store_12;
  reg                 io_in_r_bypass_regNext_9_0_df_is_ws_12;
  reg                 io_in_r_bypass_regNext_9_0_stall_12;
  reg        [15:0]   io_in_r_bypass_regNext_9_1_data_12;
  reg                 io_in_r_bypass_regNext_9_1_load_store_12;
  reg                 io_in_r_bypass_regNext_9_1_df_is_ws_12;
  reg                 io_in_r_bypass_regNext_9_1_stall_12;
  reg        [15:0]   io_in_r_bypass_regNext_9_2_data_12;
  reg                 io_in_r_bypass_regNext_9_2_load_store_12;
  reg                 io_in_r_bypass_regNext_9_2_df_is_ws_12;
  reg                 io_in_r_bypass_regNext_9_2_stall_12;
  reg        [15:0]   io_in_r_bypass_regNext_9_3_data_12;
  reg                 io_in_r_bypass_regNext_9_3_load_store_12;
  reg                 io_in_r_bypass_regNext_9_3_df_is_ws_12;
  reg                 io_in_r_bypass_regNext_9_3_stall_12;
  reg        [15:0]   io_in_r_bypass_regNext_10_0_data_12;
  reg                 io_in_r_bypass_regNext_10_0_load_store_12;
  reg                 io_in_r_bypass_regNext_10_0_df_is_ws_12;
  reg                 io_in_r_bypass_regNext_10_0_stall_12;
  reg        [15:0]   io_in_r_bypass_regNext_10_1_data_12;
  reg                 io_in_r_bypass_regNext_10_1_load_store_12;
  reg                 io_in_r_bypass_regNext_10_1_df_is_ws_12;
  reg                 io_in_r_bypass_regNext_10_1_stall_12;
  reg        [15:0]   io_in_r_bypass_regNext_10_2_data_12;
  reg                 io_in_r_bypass_regNext_10_2_load_store_12;
  reg                 io_in_r_bypass_regNext_10_2_df_is_ws_12;
  reg                 io_in_r_bypass_regNext_10_2_stall_12;
  reg        [15:0]   io_in_r_bypass_regNext_10_3_data_12;
  reg                 io_in_r_bypass_regNext_10_3_load_store_12;
  reg                 io_in_r_bypass_regNext_10_3_df_is_ws_12;
  reg                 io_in_r_bypass_regNext_10_3_stall_12;
  reg        [15:0]   io_in_r_bypass_regNext_11_0_data_12;
  reg                 io_in_r_bypass_regNext_11_0_load_store_12;
  reg                 io_in_r_bypass_regNext_11_0_df_is_ws_12;
  reg                 io_in_r_bypass_regNext_11_0_stall_12;
  reg        [15:0]   io_in_r_bypass_regNext_11_1_data_12;
  reg                 io_in_r_bypass_regNext_11_1_load_store_12;
  reg                 io_in_r_bypass_regNext_11_1_df_is_ws_12;
  reg                 io_in_r_bypass_regNext_11_1_stall_12;
  reg        [15:0]   io_in_r_bypass_regNext_11_2_data_12;
  reg                 io_in_r_bypass_regNext_11_2_load_store_12;
  reg                 io_in_r_bypass_regNext_11_2_df_is_ws_12;
  reg                 io_in_r_bypass_regNext_11_2_stall_12;
  reg        [15:0]   io_in_r_bypass_regNext_11_3_data_12;
  reg                 io_in_r_bypass_regNext_11_3_load_store_12;
  reg                 io_in_r_bypass_regNext_11_3_df_is_ws_12;
  reg                 io_in_r_bypass_regNext_11_3_stall_12;
  reg        [15:0]   io_in_r_bypass_regNext_12_0_data_12;
  reg                 io_in_r_bypass_regNext_12_0_load_store_12;
  reg                 io_in_r_bypass_regNext_12_0_df_is_ws_12;
  reg                 io_in_r_bypass_regNext_12_0_stall_12;
  reg        [15:0]   io_in_r_bypass_regNext_12_1_data_12;
  reg                 io_in_r_bypass_regNext_12_1_load_store_12;
  reg                 io_in_r_bypass_regNext_12_1_df_is_ws_12;
  reg                 io_in_r_bypass_regNext_12_1_stall_12;
  reg        [15:0]   io_in_r_bypass_regNext_12_2_data_12;
  reg                 io_in_r_bypass_regNext_12_2_load_store_12;
  reg                 io_in_r_bypass_regNext_12_2_df_is_ws_12;
  reg                 io_in_r_bypass_regNext_12_2_stall_12;
  reg        [15:0]   io_in_r_bypass_regNext_12_3_data_12;
  reg                 io_in_r_bypass_regNext_12_3_load_store_12;
  reg                 io_in_r_bypass_regNext_12_3_df_is_ws_12;
  reg                 io_in_r_bypass_regNext_12_3_stall_12;
  reg        [15:0]   io_in_r_bypass_regNext_13_0_data_12;
  reg                 io_in_r_bypass_regNext_13_0_load_store_12;
  reg                 io_in_r_bypass_regNext_13_0_df_is_ws_12;
  reg                 io_in_r_bypass_regNext_13_0_stall_12;
  reg        [15:0]   io_in_r_bypass_regNext_13_1_data_12;
  reg                 io_in_r_bypass_regNext_13_1_load_store_12;
  reg                 io_in_r_bypass_regNext_13_1_df_is_ws_12;
  reg                 io_in_r_bypass_regNext_13_1_stall_12;
  reg        [15:0]   io_in_r_bypass_regNext_13_2_data_12;
  reg                 io_in_r_bypass_regNext_13_2_load_store_12;
  reg                 io_in_r_bypass_regNext_13_2_df_is_ws_12;
  reg                 io_in_r_bypass_regNext_13_2_stall_12;
  reg        [15:0]   io_in_r_bypass_regNext_13_3_data_12;
  reg                 io_in_r_bypass_regNext_13_3_load_store_12;
  reg                 io_in_r_bypass_regNext_13_3_df_is_ws_12;
  reg                 io_in_r_bypass_regNext_13_3_stall_12;
  reg        [15:0]   io_in_r_bypass_regNext_14_0_data_12;
  reg                 io_in_r_bypass_regNext_14_0_load_store_12;
  reg                 io_in_r_bypass_regNext_14_0_df_is_ws_12;
  reg                 io_in_r_bypass_regNext_14_0_stall_12;
  reg        [15:0]   io_in_r_bypass_regNext_14_1_data_12;
  reg                 io_in_r_bypass_regNext_14_1_load_store_12;
  reg                 io_in_r_bypass_regNext_14_1_df_is_ws_12;
  reg                 io_in_r_bypass_regNext_14_1_stall_12;
  reg        [15:0]   io_in_r_bypass_regNext_14_2_data_12;
  reg                 io_in_r_bypass_regNext_14_2_load_store_12;
  reg                 io_in_r_bypass_regNext_14_2_df_is_ws_12;
  reg                 io_in_r_bypass_regNext_14_2_stall_12;
  reg        [15:0]   io_in_r_bypass_regNext_14_3_data_12;
  reg                 io_in_r_bypass_regNext_14_3_load_store_12;
  reg                 io_in_r_bypass_regNext_14_3_df_is_ws_12;
  reg                 io_in_r_bypass_regNext_14_3_stall_12;
  reg        [15:0]   io_in_r_bypass_regNext_15_0_data_12;
  reg                 io_in_r_bypass_regNext_15_0_load_store_12;
  reg                 io_in_r_bypass_regNext_15_0_df_is_ws_12;
  reg                 io_in_r_bypass_regNext_15_0_stall_12;
  reg        [15:0]   io_in_r_bypass_regNext_15_1_data_12;
  reg                 io_in_r_bypass_regNext_15_1_load_store_12;
  reg                 io_in_r_bypass_regNext_15_1_df_is_ws_12;
  reg                 io_in_r_bypass_regNext_15_1_stall_12;
  reg        [15:0]   io_in_r_bypass_regNext_15_2_data_12;
  reg                 io_in_r_bypass_regNext_15_2_load_store_12;
  reg                 io_in_r_bypass_regNext_15_2_df_is_ws_12;
  reg                 io_in_r_bypass_regNext_15_2_stall_12;
  reg        [15:0]   io_in_r_bypass_regNext_15_3_data_12;
  reg                 io_in_r_bypass_regNext_15_3_load_store_12;
  reg                 io_in_r_bypass_regNext_15_3_df_is_ws_12;
  reg                 io_in_r_bypass_regNext_15_3_stall_12;
  reg        [15:0]   io_in_r_bypass_regNext_16_0_data_12;
  reg                 io_in_r_bypass_regNext_16_0_load_store_12;
  reg                 io_in_r_bypass_regNext_16_0_df_is_ws_12;
  reg                 io_in_r_bypass_regNext_16_0_stall_12;
  reg        [15:0]   io_in_r_bypass_regNext_16_1_data_12;
  reg                 io_in_r_bypass_regNext_16_1_load_store_12;
  reg                 io_in_r_bypass_regNext_16_1_df_is_ws_12;
  reg                 io_in_r_bypass_regNext_16_1_stall_12;
  reg        [15:0]   io_in_r_bypass_regNext_16_2_data_12;
  reg                 io_in_r_bypass_regNext_16_2_load_store_12;
  reg                 io_in_r_bypass_regNext_16_2_df_is_ws_12;
  reg                 io_in_r_bypass_regNext_16_2_stall_12;
  reg        [15:0]   io_in_r_bypass_regNext_16_3_data_12;
  reg                 io_in_r_bypass_regNext_16_3_load_store_12;
  reg                 io_in_r_bypass_regNext_16_3_df_is_ws_12;
  reg                 io_in_r_bypass_regNext_16_3_stall_12;
  reg        [15:0]   io_in_r_bypass_regNext_17_0_data_12;
  reg                 io_in_r_bypass_regNext_17_0_load_store_12;
  reg                 io_in_r_bypass_regNext_17_0_df_is_ws_12;
  reg                 io_in_r_bypass_regNext_17_0_stall_12;
  reg        [15:0]   io_in_r_bypass_regNext_17_1_data_12;
  reg                 io_in_r_bypass_regNext_17_1_load_store_12;
  reg                 io_in_r_bypass_regNext_17_1_df_is_ws_12;
  reg                 io_in_r_bypass_regNext_17_1_stall_12;
  reg        [15:0]   io_in_r_bypass_regNext_17_2_data_12;
  reg                 io_in_r_bypass_regNext_17_2_load_store_12;
  reg                 io_in_r_bypass_regNext_17_2_df_is_ws_12;
  reg                 io_in_r_bypass_regNext_17_2_stall_12;
  reg        [15:0]   io_in_r_bypass_regNext_17_3_data_12;
  reg                 io_in_r_bypass_regNext_17_3_load_store_12;
  reg                 io_in_r_bypass_regNext_17_3_df_is_ws_12;
  reg                 io_in_r_bypass_regNext_17_3_stall_12;
  reg        [15:0]   io_in_r_bypass_regNext_18_0_data_12;
  reg                 io_in_r_bypass_regNext_18_0_load_store_12;
  reg                 io_in_r_bypass_regNext_18_0_df_is_ws_12;
  reg                 io_in_r_bypass_regNext_18_0_stall_12;
  reg        [15:0]   io_in_r_bypass_regNext_18_1_data_12;
  reg                 io_in_r_bypass_regNext_18_1_load_store_12;
  reg                 io_in_r_bypass_regNext_18_1_df_is_ws_12;
  reg                 io_in_r_bypass_regNext_18_1_stall_12;
  reg        [15:0]   io_in_r_bypass_regNext_18_2_data_12;
  reg                 io_in_r_bypass_regNext_18_2_load_store_12;
  reg                 io_in_r_bypass_regNext_18_2_df_is_ws_12;
  reg                 io_in_r_bypass_regNext_18_2_stall_12;
  reg        [15:0]   io_in_r_bypass_regNext_18_3_data_12;
  reg                 io_in_r_bypass_regNext_18_3_load_store_12;
  reg                 io_in_r_bypass_regNext_18_3_df_is_ws_12;
  reg                 io_in_r_bypass_regNext_18_3_stall_12;
  reg        [15:0]   io_in_r_bypass_regNext_19_0_data_12;
  reg                 io_in_r_bypass_regNext_19_0_load_store_12;
  reg                 io_in_r_bypass_regNext_19_0_df_is_ws_12;
  reg                 io_in_r_bypass_regNext_19_0_stall_12;
  reg        [15:0]   io_in_r_bypass_regNext_19_1_data_12;
  reg                 io_in_r_bypass_regNext_19_1_load_store_12;
  reg                 io_in_r_bypass_regNext_19_1_df_is_ws_12;
  reg                 io_in_r_bypass_regNext_19_1_stall_12;
  reg        [15:0]   io_in_r_bypass_regNext_19_2_data_12;
  reg                 io_in_r_bypass_regNext_19_2_load_store_12;
  reg                 io_in_r_bypass_regNext_19_2_df_is_ws_12;
  reg                 io_in_r_bypass_regNext_19_2_stall_12;
  reg        [15:0]   io_in_r_bypass_regNext_19_3_data_12;
  reg                 io_in_r_bypass_regNext_19_3_load_store_12;
  reg                 io_in_r_bypass_regNext_19_3_df_is_ws_12;
  reg                 io_in_r_bypass_regNext_19_3_stall_12;
  reg        [15:0]   io_in_r_bypass_regNext_20_0_data_12;
  reg                 io_in_r_bypass_regNext_20_0_load_store_12;
  reg                 io_in_r_bypass_regNext_20_0_df_is_ws_12;
  reg                 io_in_r_bypass_regNext_20_0_stall_12;
  reg        [15:0]   io_in_r_bypass_regNext_20_1_data_12;
  reg                 io_in_r_bypass_regNext_20_1_load_store_12;
  reg                 io_in_r_bypass_regNext_20_1_df_is_ws_12;
  reg                 io_in_r_bypass_regNext_20_1_stall_12;
  reg        [15:0]   io_in_r_bypass_regNext_20_2_data_12;
  reg                 io_in_r_bypass_regNext_20_2_load_store_12;
  reg                 io_in_r_bypass_regNext_20_2_df_is_ws_12;
  reg                 io_in_r_bypass_regNext_20_2_stall_12;
  reg        [15:0]   io_in_r_bypass_regNext_20_3_data_12;
  reg                 io_in_r_bypass_regNext_20_3_load_store_12;
  reg                 io_in_r_bypass_regNext_20_3_df_is_ws_12;
  reg                 io_in_r_bypass_regNext_20_3_stall_12;
  reg        [15:0]   io_in_r_bypass_regNext_21_0_data_12;
  reg                 io_in_r_bypass_regNext_21_0_load_store_12;
  reg                 io_in_r_bypass_regNext_21_0_df_is_ws_12;
  reg                 io_in_r_bypass_regNext_21_0_stall_12;
  reg        [15:0]   io_in_r_bypass_regNext_21_1_data_12;
  reg                 io_in_r_bypass_regNext_21_1_load_store_12;
  reg                 io_in_r_bypass_regNext_21_1_df_is_ws_12;
  reg                 io_in_r_bypass_regNext_21_1_stall_12;
  reg        [15:0]   io_in_r_bypass_regNext_21_2_data_12;
  reg                 io_in_r_bypass_regNext_21_2_load_store_12;
  reg                 io_in_r_bypass_regNext_21_2_df_is_ws_12;
  reg                 io_in_r_bypass_regNext_21_2_stall_12;
  reg        [15:0]   io_in_r_bypass_regNext_21_3_data_12;
  reg                 io_in_r_bypass_regNext_21_3_load_store_12;
  reg                 io_in_r_bypass_regNext_21_3_df_is_ws_12;
  reg                 io_in_r_bypass_regNext_21_3_stall_12;
  reg        [15:0]   io_in_r_bypass_regNext_22_0_data_12;
  reg                 io_in_r_bypass_regNext_22_0_load_store_12;
  reg                 io_in_r_bypass_regNext_22_0_df_is_ws_12;
  reg                 io_in_r_bypass_regNext_22_0_stall_12;
  reg        [15:0]   io_in_r_bypass_regNext_22_1_data_12;
  reg                 io_in_r_bypass_regNext_22_1_load_store_12;
  reg                 io_in_r_bypass_regNext_22_1_df_is_ws_12;
  reg                 io_in_r_bypass_regNext_22_1_stall_12;
  reg        [15:0]   io_in_r_bypass_regNext_22_2_data_12;
  reg                 io_in_r_bypass_regNext_22_2_load_store_12;
  reg                 io_in_r_bypass_regNext_22_2_df_is_ws_12;
  reg                 io_in_r_bypass_regNext_22_2_stall_12;
  reg        [15:0]   io_in_r_bypass_regNext_22_3_data_12;
  reg                 io_in_r_bypass_regNext_22_3_load_store_12;
  reg                 io_in_r_bypass_regNext_22_3_df_is_ws_12;
  reg                 io_in_r_bypass_regNext_22_3_stall_12;
  reg        [15:0]   io_in_r_bypass_regNext_23_0_data_12;
  reg                 io_in_r_bypass_regNext_23_0_load_store_12;
  reg                 io_in_r_bypass_regNext_23_0_df_is_ws_12;
  reg                 io_in_r_bypass_regNext_23_0_stall_12;
  reg        [15:0]   io_in_r_bypass_regNext_23_1_data_12;
  reg                 io_in_r_bypass_regNext_23_1_load_store_12;
  reg                 io_in_r_bypass_regNext_23_1_df_is_ws_12;
  reg                 io_in_r_bypass_regNext_23_1_stall_12;
  reg        [15:0]   io_in_r_bypass_regNext_23_2_data_12;
  reg                 io_in_r_bypass_regNext_23_2_load_store_12;
  reg                 io_in_r_bypass_regNext_23_2_df_is_ws_12;
  reg                 io_in_r_bypass_regNext_23_2_stall_12;
  reg        [15:0]   io_in_r_bypass_regNext_23_3_data_12;
  reg                 io_in_r_bypass_regNext_23_3_load_store_12;
  reg                 io_in_r_bypass_regNext_23_3_df_is_ws_12;
  reg                 io_in_r_bypass_regNext_23_3_stall_12;
  reg        [15:0]   io_in_r_bypass_regNext_24_0_data_12;
  reg                 io_in_r_bypass_regNext_24_0_load_store_12;
  reg                 io_in_r_bypass_regNext_24_0_df_is_ws_12;
  reg                 io_in_r_bypass_regNext_24_0_stall_12;
  reg        [15:0]   io_in_r_bypass_regNext_24_1_data_12;
  reg                 io_in_r_bypass_regNext_24_1_load_store_12;
  reg                 io_in_r_bypass_regNext_24_1_df_is_ws_12;
  reg                 io_in_r_bypass_regNext_24_1_stall_12;
  reg        [15:0]   io_in_r_bypass_regNext_24_2_data_12;
  reg                 io_in_r_bypass_regNext_24_2_load_store_12;
  reg                 io_in_r_bypass_regNext_24_2_df_is_ws_12;
  reg                 io_in_r_bypass_regNext_24_2_stall_12;
  reg        [15:0]   io_in_r_bypass_regNext_24_3_data_12;
  reg                 io_in_r_bypass_regNext_24_3_load_store_12;
  reg                 io_in_r_bypass_regNext_24_3_df_is_ws_12;
  reg                 io_in_r_bypass_regNext_24_3_stall_12;
  reg        [15:0]   io_in_r_bypass_regNext_25_0_data_12;
  reg                 io_in_r_bypass_regNext_25_0_load_store_12;
  reg                 io_in_r_bypass_regNext_25_0_df_is_ws_12;
  reg                 io_in_r_bypass_regNext_25_0_stall_12;
  reg        [15:0]   io_in_r_bypass_regNext_25_1_data_12;
  reg                 io_in_r_bypass_regNext_25_1_load_store_12;
  reg                 io_in_r_bypass_regNext_25_1_df_is_ws_12;
  reg                 io_in_r_bypass_regNext_25_1_stall_12;
  reg        [15:0]   io_in_r_bypass_regNext_25_2_data_12;
  reg                 io_in_r_bypass_regNext_25_2_load_store_12;
  reg                 io_in_r_bypass_regNext_25_2_df_is_ws_12;
  reg                 io_in_r_bypass_regNext_25_2_stall_12;
  reg        [15:0]   io_in_r_bypass_regNext_25_3_data_12;
  reg                 io_in_r_bypass_regNext_25_3_load_store_12;
  reg                 io_in_r_bypass_regNext_25_3_df_is_ws_12;
  reg                 io_in_r_bypass_regNext_25_3_stall_12;
  reg        [15:0]   io_in_r_bypass_regNext_26_0_data_12;
  reg                 io_in_r_bypass_regNext_26_0_load_store_12;
  reg                 io_in_r_bypass_regNext_26_0_df_is_ws_12;
  reg                 io_in_r_bypass_regNext_26_0_stall_12;
  reg        [15:0]   io_in_r_bypass_regNext_26_1_data_12;
  reg                 io_in_r_bypass_regNext_26_1_load_store_12;
  reg                 io_in_r_bypass_regNext_26_1_df_is_ws_12;
  reg                 io_in_r_bypass_regNext_26_1_stall_12;
  reg        [15:0]   io_in_r_bypass_regNext_26_2_data_12;
  reg                 io_in_r_bypass_regNext_26_2_load_store_12;
  reg                 io_in_r_bypass_regNext_26_2_df_is_ws_12;
  reg                 io_in_r_bypass_regNext_26_2_stall_12;
  reg        [15:0]   io_in_r_bypass_regNext_26_3_data_12;
  reg                 io_in_r_bypass_regNext_26_3_load_store_12;
  reg                 io_in_r_bypass_regNext_26_3_df_is_ws_12;
  reg                 io_in_r_bypass_regNext_26_3_stall_12;
  reg        [15:0]   io_in_r_bypass_regNext_27_0_data_12;
  reg                 io_in_r_bypass_regNext_27_0_load_store_12;
  reg                 io_in_r_bypass_regNext_27_0_df_is_ws_12;
  reg                 io_in_r_bypass_regNext_27_0_stall_12;
  reg        [15:0]   io_in_r_bypass_regNext_27_1_data_12;
  reg                 io_in_r_bypass_regNext_27_1_load_store_12;
  reg                 io_in_r_bypass_regNext_27_1_df_is_ws_12;
  reg                 io_in_r_bypass_regNext_27_1_stall_12;
  reg        [15:0]   io_in_r_bypass_regNext_27_2_data_12;
  reg                 io_in_r_bypass_regNext_27_2_load_store_12;
  reg                 io_in_r_bypass_regNext_27_2_df_is_ws_12;
  reg                 io_in_r_bypass_regNext_27_2_stall_12;
  reg        [15:0]   io_in_r_bypass_regNext_27_3_data_12;
  reg                 io_in_r_bypass_regNext_27_3_load_store_12;
  reg                 io_in_r_bypass_regNext_27_3_df_is_ws_12;
  reg                 io_in_r_bypass_regNext_27_3_stall_12;
  reg        [15:0]   io_in_r_bypass_regNext_28_0_data_12;
  reg                 io_in_r_bypass_regNext_28_0_load_store_12;
  reg                 io_in_r_bypass_regNext_28_0_df_is_ws_12;
  reg                 io_in_r_bypass_regNext_28_0_stall_12;
  reg        [15:0]   io_in_r_bypass_regNext_28_1_data_12;
  reg                 io_in_r_bypass_regNext_28_1_load_store_12;
  reg                 io_in_r_bypass_regNext_28_1_df_is_ws_12;
  reg                 io_in_r_bypass_regNext_28_1_stall_12;
  reg        [15:0]   io_in_r_bypass_regNext_28_2_data_12;
  reg                 io_in_r_bypass_regNext_28_2_load_store_12;
  reg                 io_in_r_bypass_regNext_28_2_df_is_ws_12;
  reg                 io_in_r_bypass_regNext_28_2_stall_12;
  reg        [15:0]   io_in_r_bypass_regNext_28_3_data_12;
  reg                 io_in_r_bypass_regNext_28_3_load_store_12;
  reg                 io_in_r_bypass_regNext_28_3_df_is_ws_12;
  reg                 io_in_r_bypass_regNext_28_3_stall_12;
  reg        [15:0]   io_in_r_bypass_regNext_29_0_data_12;
  reg                 io_in_r_bypass_regNext_29_0_load_store_12;
  reg                 io_in_r_bypass_regNext_29_0_df_is_ws_12;
  reg                 io_in_r_bypass_regNext_29_0_stall_12;
  reg        [15:0]   io_in_r_bypass_regNext_29_1_data_12;
  reg                 io_in_r_bypass_regNext_29_1_load_store_12;
  reg                 io_in_r_bypass_regNext_29_1_df_is_ws_12;
  reg                 io_in_r_bypass_regNext_29_1_stall_12;
  reg        [15:0]   io_in_r_bypass_regNext_29_2_data_12;
  reg                 io_in_r_bypass_regNext_29_2_load_store_12;
  reg                 io_in_r_bypass_regNext_29_2_df_is_ws_12;
  reg                 io_in_r_bypass_regNext_29_2_stall_12;
  reg        [15:0]   io_in_r_bypass_regNext_29_3_data_12;
  reg                 io_in_r_bypass_regNext_29_3_load_store_12;
  reg                 io_in_r_bypass_regNext_29_3_df_is_ws_12;
  reg                 io_in_r_bypass_regNext_29_3_stall_12;
  reg        [15:0]   io_in_r_bypass_regNext_30_0_data_12;
  reg                 io_in_r_bypass_regNext_30_0_load_store_12;
  reg                 io_in_r_bypass_regNext_30_0_df_is_ws_12;
  reg                 io_in_r_bypass_regNext_30_0_stall_12;
  reg        [15:0]   io_in_r_bypass_regNext_30_1_data_12;
  reg                 io_in_r_bypass_regNext_30_1_load_store_12;
  reg                 io_in_r_bypass_regNext_30_1_df_is_ws_12;
  reg                 io_in_r_bypass_regNext_30_1_stall_12;
  reg        [15:0]   io_in_r_bypass_regNext_30_2_data_12;
  reg                 io_in_r_bypass_regNext_30_2_load_store_12;
  reg                 io_in_r_bypass_regNext_30_2_df_is_ws_12;
  reg                 io_in_r_bypass_regNext_30_2_stall_12;
  reg        [15:0]   io_in_r_bypass_regNext_30_3_data_12;
  reg                 io_in_r_bypass_regNext_30_3_load_store_12;
  reg                 io_in_r_bypass_regNext_30_3_df_is_ws_12;
  reg                 io_in_r_bypass_regNext_30_3_stall_12;
  reg        [15:0]   io_in_r_bypass_regNext_31_0_data_12;
  reg                 io_in_r_bypass_regNext_31_0_load_store_12;
  reg                 io_in_r_bypass_regNext_31_0_df_is_ws_12;
  reg                 io_in_r_bypass_regNext_31_0_stall_12;
  reg        [15:0]   io_in_r_bypass_regNext_31_1_data_12;
  reg                 io_in_r_bypass_regNext_31_1_load_store_12;
  reg                 io_in_r_bypass_regNext_31_1_df_is_ws_12;
  reg                 io_in_r_bypass_regNext_31_1_stall_12;
  reg        [15:0]   io_in_r_bypass_regNext_31_2_data_12;
  reg                 io_in_r_bypass_regNext_31_2_load_store_12;
  reg                 io_in_r_bypass_regNext_31_2_df_is_ws_12;
  reg                 io_in_r_bypass_regNext_31_2_stall_12;
  reg        [15:0]   io_in_r_bypass_regNext_31_3_data_12;
  reg                 io_in_r_bypass_regNext_31_3_load_store_12;
  reg                 io_in_r_bypass_regNext_31_3_df_is_ws_12;
  reg                 io_in_r_bypass_regNext_31_3_stall_12;
  reg        [15:0]   io_in_r_bypass_regNext_0_0_data_13;
  reg                 io_in_r_bypass_regNext_0_0_load_store_13;
  reg                 io_in_r_bypass_regNext_0_0_df_is_ws_13;
  reg                 io_in_r_bypass_regNext_0_0_stall_13;
  reg        [15:0]   io_in_r_bypass_regNext_0_1_data_13;
  reg                 io_in_r_bypass_regNext_0_1_load_store_13;
  reg                 io_in_r_bypass_regNext_0_1_df_is_ws_13;
  reg                 io_in_r_bypass_regNext_0_1_stall_13;
  reg        [15:0]   io_in_r_bypass_regNext_0_2_data_13;
  reg                 io_in_r_bypass_regNext_0_2_load_store_13;
  reg                 io_in_r_bypass_regNext_0_2_df_is_ws_13;
  reg                 io_in_r_bypass_regNext_0_2_stall_13;
  reg        [15:0]   io_in_r_bypass_regNext_0_3_data_13;
  reg                 io_in_r_bypass_regNext_0_3_load_store_13;
  reg                 io_in_r_bypass_regNext_0_3_df_is_ws_13;
  reg                 io_in_r_bypass_regNext_0_3_stall_13;
  reg        [15:0]   io_in_r_bypass_regNext_1_0_data_13;
  reg                 io_in_r_bypass_regNext_1_0_load_store_13;
  reg                 io_in_r_bypass_regNext_1_0_df_is_ws_13;
  reg                 io_in_r_bypass_regNext_1_0_stall_13;
  reg        [15:0]   io_in_r_bypass_regNext_1_1_data_13;
  reg                 io_in_r_bypass_regNext_1_1_load_store_13;
  reg                 io_in_r_bypass_regNext_1_1_df_is_ws_13;
  reg                 io_in_r_bypass_regNext_1_1_stall_13;
  reg        [15:0]   io_in_r_bypass_regNext_1_2_data_13;
  reg                 io_in_r_bypass_regNext_1_2_load_store_13;
  reg                 io_in_r_bypass_regNext_1_2_df_is_ws_13;
  reg                 io_in_r_bypass_regNext_1_2_stall_13;
  reg        [15:0]   io_in_r_bypass_regNext_1_3_data_13;
  reg                 io_in_r_bypass_regNext_1_3_load_store_13;
  reg                 io_in_r_bypass_regNext_1_3_df_is_ws_13;
  reg                 io_in_r_bypass_regNext_1_3_stall_13;
  reg        [15:0]   io_in_r_bypass_regNext_2_0_data_13;
  reg                 io_in_r_bypass_regNext_2_0_load_store_13;
  reg                 io_in_r_bypass_regNext_2_0_df_is_ws_13;
  reg                 io_in_r_bypass_regNext_2_0_stall_13;
  reg        [15:0]   io_in_r_bypass_regNext_2_1_data_13;
  reg                 io_in_r_bypass_regNext_2_1_load_store_13;
  reg                 io_in_r_bypass_regNext_2_1_df_is_ws_13;
  reg                 io_in_r_bypass_regNext_2_1_stall_13;
  reg        [15:0]   io_in_r_bypass_regNext_2_2_data_13;
  reg                 io_in_r_bypass_regNext_2_2_load_store_13;
  reg                 io_in_r_bypass_regNext_2_2_df_is_ws_13;
  reg                 io_in_r_bypass_regNext_2_2_stall_13;
  reg        [15:0]   io_in_r_bypass_regNext_2_3_data_13;
  reg                 io_in_r_bypass_regNext_2_3_load_store_13;
  reg                 io_in_r_bypass_regNext_2_3_df_is_ws_13;
  reg                 io_in_r_bypass_regNext_2_3_stall_13;
  reg        [15:0]   io_in_r_bypass_regNext_3_0_data_13;
  reg                 io_in_r_bypass_regNext_3_0_load_store_13;
  reg                 io_in_r_bypass_regNext_3_0_df_is_ws_13;
  reg                 io_in_r_bypass_regNext_3_0_stall_13;
  reg        [15:0]   io_in_r_bypass_regNext_3_1_data_13;
  reg                 io_in_r_bypass_regNext_3_1_load_store_13;
  reg                 io_in_r_bypass_regNext_3_1_df_is_ws_13;
  reg                 io_in_r_bypass_regNext_3_1_stall_13;
  reg        [15:0]   io_in_r_bypass_regNext_3_2_data_13;
  reg                 io_in_r_bypass_regNext_3_2_load_store_13;
  reg                 io_in_r_bypass_regNext_3_2_df_is_ws_13;
  reg                 io_in_r_bypass_regNext_3_2_stall_13;
  reg        [15:0]   io_in_r_bypass_regNext_3_3_data_13;
  reg                 io_in_r_bypass_regNext_3_3_load_store_13;
  reg                 io_in_r_bypass_regNext_3_3_df_is_ws_13;
  reg                 io_in_r_bypass_regNext_3_3_stall_13;
  reg        [15:0]   io_in_r_bypass_regNext_4_0_data_13;
  reg                 io_in_r_bypass_regNext_4_0_load_store_13;
  reg                 io_in_r_bypass_regNext_4_0_df_is_ws_13;
  reg                 io_in_r_bypass_regNext_4_0_stall_13;
  reg        [15:0]   io_in_r_bypass_regNext_4_1_data_13;
  reg                 io_in_r_bypass_regNext_4_1_load_store_13;
  reg                 io_in_r_bypass_regNext_4_1_df_is_ws_13;
  reg                 io_in_r_bypass_regNext_4_1_stall_13;
  reg        [15:0]   io_in_r_bypass_regNext_4_2_data_13;
  reg                 io_in_r_bypass_regNext_4_2_load_store_13;
  reg                 io_in_r_bypass_regNext_4_2_df_is_ws_13;
  reg                 io_in_r_bypass_regNext_4_2_stall_13;
  reg        [15:0]   io_in_r_bypass_regNext_4_3_data_13;
  reg                 io_in_r_bypass_regNext_4_3_load_store_13;
  reg                 io_in_r_bypass_regNext_4_3_df_is_ws_13;
  reg                 io_in_r_bypass_regNext_4_3_stall_13;
  reg        [15:0]   io_in_r_bypass_regNext_5_0_data_13;
  reg                 io_in_r_bypass_regNext_5_0_load_store_13;
  reg                 io_in_r_bypass_regNext_5_0_df_is_ws_13;
  reg                 io_in_r_bypass_regNext_5_0_stall_13;
  reg        [15:0]   io_in_r_bypass_regNext_5_1_data_13;
  reg                 io_in_r_bypass_regNext_5_1_load_store_13;
  reg                 io_in_r_bypass_regNext_5_1_df_is_ws_13;
  reg                 io_in_r_bypass_regNext_5_1_stall_13;
  reg        [15:0]   io_in_r_bypass_regNext_5_2_data_13;
  reg                 io_in_r_bypass_regNext_5_2_load_store_13;
  reg                 io_in_r_bypass_regNext_5_2_df_is_ws_13;
  reg                 io_in_r_bypass_regNext_5_2_stall_13;
  reg        [15:0]   io_in_r_bypass_regNext_5_3_data_13;
  reg                 io_in_r_bypass_regNext_5_3_load_store_13;
  reg                 io_in_r_bypass_regNext_5_3_df_is_ws_13;
  reg                 io_in_r_bypass_regNext_5_3_stall_13;
  reg        [15:0]   io_in_r_bypass_regNext_6_0_data_13;
  reg                 io_in_r_bypass_regNext_6_0_load_store_13;
  reg                 io_in_r_bypass_regNext_6_0_df_is_ws_13;
  reg                 io_in_r_bypass_regNext_6_0_stall_13;
  reg        [15:0]   io_in_r_bypass_regNext_6_1_data_13;
  reg                 io_in_r_bypass_regNext_6_1_load_store_13;
  reg                 io_in_r_bypass_regNext_6_1_df_is_ws_13;
  reg                 io_in_r_bypass_regNext_6_1_stall_13;
  reg        [15:0]   io_in_r_bypass_regNext_6_2_data_13;
  reg                 io_in_r_bypass_regNext_6_2_load_store_13;
  reg                 io_in_r_bypass_regNext_6_2_df_is_ws_13;
  reg                 io_in_r_bypass_regNext_6_2_stall_13;
  reg        [15:0]   io_in_r_bypass_regNext_6_3_data_13;
  reg                 io_in_r_bypass_regNext_6_3_load_store_13;
  reg                 io_in_r_bypass_regNext_6_3_df_is_ws_13;
  reg                 io_in_r_bypass_regNext_6_3_stall_13;
  reg        [15:0]   io_in_r_bypass_regNext_7_0_data_13;
  reg                 io_in_r_bypass_regNext_7_0_load_store_13;
  reg                 io_in_r_bypass_regNext_7_0_df_is_ws_13;
  reg                 io_in_r_bypass_regNext_7_0_stall_13;
  reg        [15:0]   io_in_r_bypass_regNext_7_1_data_13;
  reg                 io_in_r_bypass_regNext_7_1_load_store_13;
  reg                 io_in_r_bypass_regNext_7_1_df_is_ws_13;
  reg                 io_in_r_bypass_regNext_7_1_stall_13;
  reg        [15:0]   io_in_r_bypass_regNext_7_2_data_13;
  reg                 io_in_r_bypass_regNext_7_2_load_store_13;
  reg                 io_in_r_bypass_regNext_7_2_df_is_ws_13;
  reg                 io_in_r_bypass_regNext_7_2_stall_13;
  reg        [15:0]   io_in_r_bypass_regNext_7_3_data_13;
  reg                 io_in_r_bypass_regNext_7_3_load_store_13;
  reg                 io_in_r_bypass_regNext_7_3_df_is_ws_13;
  reg                 io_in_r_bypass_regNext_7_3_stall_13;
  reg        [15:0]   io_in_r_bypass_regNext_8_0_data_13;
  reg                 io_in_r_bypass_regNext_8_0_load_store_13;
  reg                 io_in_r_bypass_regNext_8_0_df_is_ws_13;
  reg                 io_in_r_bypass_regNext_8_0_stall_13;
  reg        [15:0]   io_in_r_bypass_regNext_8_1_data_13;
  reg                 io_in_r_bypass_regNext_8_1_load_store_13;
  reg                 io_in_r_bypass_regNext_8_1_df_is_ws_13;
  reg                 io_in_r_bypass_regNext_8_1_stall_13;
  reg        [15:0]   io_in_r_bypass_regNext_8_2_data_13;
  reg                 io_in_r_bypass_regNext_8_2_load_store_13;
  reg                 io_in_r_bypass_regNext_8_2_df_is_ws_13;
  reg                 io_in_r_bypass_regNext_8_2_stall_13;
  reg        [15:0]   io_in_r_bypass_regNext_8_3_data_13;
  reg                 io_in_r_bypass_regNext_8_3_load_store_13;
  reg                 io_in_r_bypass_regNext_8_3_df_is_ws_13;
  reg                 io_in_r_bypass_regNext_8_3_stall_13;
  reg        [15:0]   io_in_r_bypass_regNext_9_0_data_13;
  reg                 io_in_r_bypass_regNext_9_0_load_store_13;
  reg                 io_in_r_bypass_regNext_9_0_df_is_ws_13;
  reg                 io_in_r_bypass_regNext_9_0_stall_13;
  reg        [15:0]   io_in_r_bypass_regNext_9_1_data_13;
  reg                 io_in_r_bypass_regNext_9_1_load_store_13;
  reg                 io_in_r_bypass_regNext_9_1_df_is_ws_13;
  reg                 io_in_r_bypass_regNext_9_1_stall_13;
  reg        [15:0]   io_in_r_bypass_regNext_9_2_data_13;
  reg                 io_in_r_bypass_regNext_9_2_load_store_13;
  reg                 io_in_r_bypass_regNext_9_2_df_is_ws_13;
  reg                 io_in_r_bypass_regNext_9_2_stall_13;
  reg        [15:0]   io_in_r_bypass_regNext_9_3_data_13;
  reg                 io_in_r_bypass_regNext_9_3_load_store_13;
  reg                 io_in_r_bypass_regNext_9_3_df_is_ws_13;
  reg                 io_in_r_bypass_regNext_9_3_stall_13;
  reg        [15:0]   io_in_r_bypass_regNext_10_0_data_13;
  reg                 io_in_r_bypass_regNext_10_0_load_store_13;
  reg                 io_in_r_bypass_regNext_10_0_df_is_ws_13;
  reg                 io_in_r_bypass_regNext_10_0_stall_13;
  reg        [15:0]   io_in_r_bypass_regNext_10_1_data_13;
  reg                 io_in_r_bypass_regNext_10_1_load_store_13;
  reg                 io_in_r_bypass_regNext_10_1_df_is_ws_13;
  reg                 io_in_r_bypass_regNext_10_1_stall_13;
  reg        [15:0]   io_in_r_bypass_regNext_10_2_data_13;
  reg                 io_in_r_bypass_regNext_10_2_load_store_13;
  reg                 io_in_r_bypass_regNext_10_2_df_is_ws_13;
  reg                 io_in_r_bypass_regNext_10_2_stall_13;
  reg        [15:0]   io_in_r_bypass_regNext_10_3_data_13;
  reg                 io_in_r_bypass_regNext_10_3_load_store_13;
  reg                 io_in_r_bypass_regNext_10_3_df_is_ws_13;
  reg                 io_in_r_bypass_regNext_10_3_stall_13;
  reg        [15:0]   io_in_r_bypass_regNext_11_0_data_13;
  reg                 io_in_r_bypass_regNext_11_0_load_store_13;
  reg                 io_in_r_bypass_regNext_11_0_df_is_ws_13;
  reg                 io_in_r_bypass_regNext_11_0_stall_13;
  reg        [15:0]   io_in_r_bypass_regNext_11_1_data_13;
  reg                 io_in_r_bypass_regNext_11_1_load_store_13;
  reg                 io_in_r_bypass_regNext_11_1_df_is_ws_13;
  reg                 io_in_r_bypass_regNext_11_1_stall_13;
  reg        [15:0]   io_in_r_bypass_regNext_11_2_data_13;
  reg                 io_in_r_bypass_regNext_11_2_load_store_13;
  reg                 io_in_r_bypass_regNext_11_2_df_is_ws_13;
  reg                 io_in_r_bypass_regNext_11_2_stall_13;
  reg        [15:0]   io_in_r_bypass_regNext_11_3_data_13;
  reg                 io_in_r_bypass_regNext_11_3_load_store_13;
  reg                 io_in_r_bypass_regNext_11_3_df_is_ws_13;
  reg                 io_in_r_bypass_regNext_11_3_stall_13;
  reg        [15:0]   io_in_r_bypass_regNext_12_0_data_13;
  reg                 io_in_r_bypass_regNext_12_0_load_store_13;
  reg                 io_in_r_bypass_regNext_12_0_df_is_ws_13;
  reg                 io_in_r_bypass_regNext_12_0_stall_13;
  reg        [15:0]   io_in_r_bypass_regNext_12_1_data_13;
  reg                 io_in_r_bypass_regNext_12_1_load_store_13;
  reg                 io_in_r_bypass_regNext_12_1_df_is_ws_13;
  reg                 io_in_r_bypass_regNext_12_1_stall_13;
  reg        [15:0]   io_in_r_bypass_regNext_12_2_data_13;
  reg                 io_in_r_bypass_regNext_12_2_load_store_13;
  reg                 io_in_r_bypass_regNext_12_2_df_is_ws_13;
  reg                 io_in_r_bypass_regNext_12_2_stall_13;
  reg        [15:0]   io_in_r_bypass_regNext_12_3_data_13;
  reg                 io_in_r_bypass_regNext_12_3_load_store_13;
  reg                 io_in_r_bypass_regNext_12_3_df_is_ws_13;
  reg                 io_in_r_bypass_regNext_12_3_stall_13;
  reg        [15:0]   io_in_r_bypass_regNext_13_0_data_13;
  reg                 io_in_r_bypass_regNext_13_0_load_store_13;
  reg                 io_in_r_bypass_regNext_13_0_df_is_ws_13;
  reg                 io_in_r_bypass_regNext_13_0_stall_13;
  reg        [15:0]   io_in_r_bypass_regNext_13_1_data_13;
  reg                 io_in_r_bypass_regNext_13_1_load_store_13;
  reg                 io_in_r_bypass_regNext_13_1_df_is_ws_13;
  reg                 io_in_r_bypass_regNext_13_1_stall_13;
  reg        [15:0]   io_in_r_bypass_regNext_13_2_data_13;
  reg                 io_in_r_bypass_regNext_13_2_load_store_13;
  reg                 io_in_r_bypass_regNext_13_2_df_is_ws_13;
  reg                 io_in_r_bypass_regNext_13_2_stall_13;
  reg        [15:0]   io_in_r_bypass_regNext_13_3_data_13;
  reg                 io_in_r_bypass_regNext_13_3_load_store_13;
  reg                 io_in_r_bypass_regNext_13_3_df_is_ws_13;
  reg                 io_in_r_bypass_regNext_13_3_stall_13;
  reg        [15:0]   io_in_r_bypass_regNext_14_0_data_13;
  reg                 io_in_r_bypass_regNext_14_0_load_store_13;
  reg                 io_in_r_bypass_regNext_14_0_df_is_ws_13;
  reg                 io_in_r_bypass_regNext_14_0_stall_13;
  reg        [15:0]   io_in_r_bypass_regNext_14_1_data_13;
  reg                 io_in_r_bypass_regNext_14_1_load_store_13;
  reg                 io_in_r_bypass_regNext_14_1_df_is_ws_13;
  reg                 io_in_r_bypass_regNext_14_1_stall_13;
  reg        [15:0]   io_in_r_bypass_regNext_14_2_data_13;
  reg                 io_in_r_bypass_regNext_14_2_load_store_13;
  reg                 io_in_r_bypass_regNext_14_2_df_is_ws_13;
  reg                 io_in_r_bypass_regNext_14_2_stall_13;
  reg        [15:0]   io_in_r_bypass_regNext_14_3_data_13;
  reg                 io_in_r_bypass_regNext_14_3_load_store_13;
  reg                 io_in_r_bypass_regNext_14_3_df_is_ws_13;
  reg                 io_in_r_bypass_regNext_14_3_stall_13;
  reg        [15:0]   io_in_r_bypass_regNext_15_0_data_13;
  reg                 io_in_r_bypass_regNext_15_0_load_store_13;
  reg                 io_in_r_bypass_regNext_15_0_df_is_ws_13;
  reg                 io_in_r_bypass_regNext_15_0_stall_13;
  reg        [15:0]   io_in_r_bypass_regNext_15_1_data_13;
  reg                 io_in_r_bypass_regNext_15_1_load_store_13;
  reg                 io_in_r_bypass_regNext_15_1_df_is_ws_13;
  reg                 io_in_r_bypass_regNext_15_1_stall_13;
  reg        [15:0]   io_in_r_bypass_regNext_15_2_data_13;
  reg                 io_in_r_bypass_regNext_15_2_load_store_13;
  reg                 io_in_r_bypass_regNext_15_2_df_is_ws_13;
  reg                 io_in_r_bypass_regNext_15_2_stall_13;
  reg        [15:0]   io_in_r_bypass_regNext_15_3_data_13;
  reg                 io_in_r_bypass_regNext_15_3_load_store_13;
  reg                 io_in_r_bypass_regNext_15_3_df_is_ws_13;
  reg                 io_in_r_bypass_regNext_15_3_stall_13;
  reg        [15:0]   io_in_r_bypass_regNext_16_0_data_13;
  reg                 io_in_r_bypass_regNext_16_0_load_store_13;
  reg                 io_in_r_bypass_regNext_16_0_df_is_ws_13;
  reg                 io_in_r_bypass_regNext_16_0_stall_13;
  reg        [15:0]   io_in_r_bypass_regNext_16_1_data_13;
  reg                 io_in_r_bypass_regNext_16_1_load_store_13;
  reg                 io_in_r_bypass_regNext_16_1_df_is_ws_13;
  reg                 io_in_r_bypass_regNext_16_1_stall_13;
  reg        [15:0]   io_in_r_bypass_regNext_16_2_data_13;
  reg                 io_in_r_bypass_regNext_16_2_load_store_13;
  reg                 io_in_r_bypass_regNext_16_2_df_is_ws_13;
  reg                 io_in_r_bypass_regNext_16_2_stall_13;
  reg        [15:0]   io_in_r_bypass_regNext_16_3_data_13;
  reg                 io_in_r_bypass_regNext_16_3_load_store_13;
  reg                 io_in_r_bypass_regNext_16_3_df_is_ws_13;
  reg                 io_in_r_bypass_regNext_16_3_stall_13;
  reg        [15:0]   io_in_r_bypass_regNext_17_0_data_13;
  reg                 io_in_r_bypass_regNext_17_0_load_store_13;
  reg                 io_in_r_bypass_regNext_17_0_df_is_ws_13;
  reg                 io_in_r_bypass_regNext_17_0_stall_13;
  reg        [15:0]   io_in_r_bypass_regNext_17_1_data_13;
  reg                 io_in_r_bypass_regNext_17_1_load_store_13;
  reg                 io_in_r_bypass_regNext_17_1_df_is_ws_13;
  reg                 io_in_r_bypass_regNext_17_1_stall_13;
  reg        [15:0]   io_in_r_bypass_regNext_17_2_data_13;
  reg                 io_in_r_bypass_regNext_17_2_load_store_13;
  reg                 io_in_r_bypass_regNext_17_2_df_is_ws_13;
  reg                 io_in_r_bypass_regNext_17_2_stall_13;
  reg        [15:0]   io_in_r_bypass_regNext_17_3_data_13;
  reg                 io_in_r_bypass_regNext_17_3_load_store_13;
  reg                 io_in_r_bypass_regNext_17_3_df_is_ws_13;
  reg                 io_in_r_bypass_regNext_17_3_stall_13;
  reg        [15:0]   io_in_r_bypass_regNext_18_0_data_13;
  reg                 io_in_r_bypass_regNext_18_0_load_store_13;
  reg                 io_in_r_bypass_regNext_18_0_df_is_ws_13;
  reg                 io_in_r_bypass_regNext_18_0_stall_13;
  reg        [15:0]   io_in_r_bypass_regNext_18_1_data_13;
  reg                 io_in_r_bypass_regNext_18_1_load_store_13;
  reg                 io_in_r_bypass_regNext_18_1_df_is_ws_13;
  reg                 io_in_r_bypass_regNext_18_1_stall_13;
  reg        [15:0]   io_in_r_bypass_regNext_18_2_data_13;
  reg                 io_in_r_bypass_regNext_18_2_load_store_13;
  reg                 io_in_r_bypass_regNext_18_2_df_is_ws_13;
  reg                 io_in_r_bypass_regNext_18_2_stall_13;
  reg        [15:0]   io_in_r_bypass_regNext_18_3_data_13;
  reg                 io_in_r_bypass_regNext_18_3_load_store_13;
  reg                 io_in_r_bypass_regNext_18_3_df_is_ws_13;
  reg                 io_in_r_bypass_regNext_18_3_stall_13;
  reg        [15:0]   io_in_r_bypass_regNext_19_0_data_13;
  reg                 io_in_r_bypass_regNext_19_0_load_store_13;
  reg                 io_in_r_bypass_regNext_19_0_df_is_ws_13;
  reg                 io_in_r_bypass_regNext_19_0_stall_13;
  reg        [15:0]   io_in_r_bypass_regNext_19_1_data_13;
  reg                 io_in_r_bypass_regNext_19_1_load_store_13;
  reg                 io_in_r_bypass_regNext_19_1_df_is_ws_13;
  reg                 io_in_r_bypass_regNext_19_1_stall_13;
  reg        [15:0]   io_in_r_bypass_regNext_19_2_data_13;
  reg                 io_in_r_bypass_regNext_19_2_load_store_13;
  reg                 io_in_r_bypass_regNext_19_2_df_is_ws_13;
  reg                 io_in_r_bypass_regNext_19_2_stall_13;
  reg        [15:0]   io_in_r_bypass_regNext_19_3_data_13;
  reg                 io_in_r_bypass_regNext_19_3_load_store_13;
  reg                 io_in_r_bypass_regNext_19_3_df_is_ws_13;
  reg                 io_in_r_bypass_regNext_19_3_stall_13;
  reg        [15:0]   io_in_r_bypass_regNext_20_0_data_13;
  reg                 io_in_r_bypass_regNext_20_0_load_store_13;
  reg                 io_in_r_bypass_regNext_20_0_df_is_ws_13;
  reg                 io_in_r_bypass_regNext_20_0_stall_13;
  reg        [15:0]   io_in_r_bypass_regNext_20_1_data_13;
  reg                 io_in_r_bypass_regNext_20_1_load_store_13;
  reg                 io_in_r_bypass_regNext_20_1_df_is_ws_13;
  reg                 io_in_r_bypass_regNext_20_1_stall_13;
  reg        [15:0]   io_in_r_bypass_regNext_20_2_data_13;
  reg                 io_in_r_bypass_regNext_20_2_load_store_13;
  reg                 io_in_r_bypass_regNext_20_2_df_is_ws_13;
  reg                 io_in_r_bypass_regNext_20_2_stall_13;
  reg        [15:0]   io_in_r_bypass_regNext_20_3_data_13;
  reg                 io_in_r_bypass_regNext_20_3_load_store_13;
  reg                 io_in_r_bypass_regNext_20_3_df_is_ws_13;
  reg                 io_in_r_bypass_regNext_20_3_stall_13;
  reg        [15:0]   io_in_r_bypass_regNext_21_0_data_13;
  reg                 io_in_r_bypass_regNext_21_0_load_store_13;
  reg                 io_in_r_bypass_regNext_21_0_df_is_ws_13;
  reg                 io_in_r_bypass_regNext_21_0_stall_13;
  reg        [15:0]   io_in_r_bypass_regNext_21_1_data_13;
  reg                 io_in_r_bypass_regNext_21_1_load_store_13;
  reg                 io_in_r_bypass_regNext_21_1_df_is_ws_13;
  reg                 io_in_r_bypass_regNext_21_1_stall_13;
  reg        [15:0]   io_in_r_bypass_regNext_21_2_data_13;
  reg                 io_in_r_bypass_regNext_21_2_load_store_13;
  reg                 io_in_r_bypass_regNext_21_2_df_is_ws_13;
  reg                 io_in_r_bypass_regNext_21_2_stall_13;
  reg        [15:0]   io_in_r_bypass_regNext_21_3_data_13;
  reg                 io_in_r_bypass_regNext_21_3_load_store_13;
  reg                 io_in_r_bypass_regNext_21_3_df_is_ws_13;
  reg                 io_in_r_bypass_regNext_21_3_stall_13;
  reg        [15:0]   io_in_r_bypass_regNext_22_0_data_13;
  reg                 io_in_r_bypass_regNext_22_0_load_store_13;
  reg                 io_in_r_bypass_regNext_22_0_df_is_ws_13;
  reg                 io_in_r_bypass_regNext_22_0_stall_13;
  reg        [15:0]   io_in_r_bypass_regNext_22_1_data_13;
  reg                 io_in_r_bypass_regNext_22_1_load_store_13;
  reg                 io_in_r_bypass_regNext_22_1_df_is_ws_13;
  reg                 io_in_r_bypass_regNext_22_1_stall_13;
  reg        [15:0]   io_in_r_bypass_regNext_22_2_data_13;
  reg                 io_in_r_bypass_regNext_22_2_load_store_13;
  reg                 io_in_r_bypass_regNext_22_2_df_is_ws_13;
  reg                 io_in_r_bypass_regNext_22_2_stall_13;
  reg        [15:0]   io_in_r_bypass_regNext_22_3_data_13;
  reg                 io_in_r_bypass_regNext_22_3_load_store_13;
  reg                 io_in_r_bypass_regNext_22_3_df_is_ws_13;
  reg                 io_in_r_bypass_regNext_22_3_stall_13;
  reg        [15:0]   io_in_r_bypass_regNext_23_0_data_13;
  reg                 io_in_r_bypass_regNext_23_0_load_store_13;
  reg                 io_in_r_bypass_regNext_23_0_df_is_ws_13;
  reg                 io_in_r_bypass_regNext_23_0_stall_13;
  reg        [15:0]   io_in_r_bypass_regNext_23_1_data_13;
  reg                 io_in_r_bypass_regNext_23_1_load_store_13;
  reg                 io_in_r_bypass_regNext_23_1_df_is_ws_13;
  reg                 io_in_r_bypass_regNext_23_1_stall_13;
  reg        [15:0]   io_in_r_bypass_regNext_23_2_data_13;
  reg                 io_in_r_bypass_regNext_23_2_load_store_13;
  reg                 io_in_r_bypass_regNext_23_2_df_is_ws_13;
  reg                 io_in_r_bypass_regNext_23_2_stall_13;
  reg        [15:0]   io_in_r_bypass_regNext_23_3_data_13;
  reg                 io_in_r_bypass_regNext_23_3_load_store_13;
  reg                 io_in_r_bypass_regNext_23_3_df_is_ws_13;
  reg                 io_in_r_bypass_regNext_23_3_stall_13;
  reg        [15:0]   io_in_r_bypass_regNext_24_0_data_13;
  reg                 io_in_r_bypass_regNext_24_0_load_store_13;
  reg                 io_in_r_bypass_regNext_24_0_df_is_ws_13;
  reg                 io_in_r_bypass_regNext_24_0_stall_13;
  reg        [15:0]   io_in_r_bypass_regNext_24_1_data_13;
  reg                 io_in_r_bypass_regNext_24_1_load_store_13;
  reg                 io_in_r_bypass_regNext_24_1_df_is_ws_13;
  reg                 io_in_r_bypass_regNext_24_1_stall_13;
  reg        [15:0]   io_in_r_bypass_regNext_24_2_data_13;
  reg                 io_in_r_bypass_regNext_24_2_load_store_13;
  reg                 io_in_r_bypass_regNext_24_2_df_is_ws_13;
  reg                 io_in_r_bypass_regNext_24_2_stall_13;
  reg        [15:0]   io_in_r_bypass_regNext_24_3_data_13;
  reg                 io_in_r_bypass_regNext_24_3_load_store_13;
  reg                 io_in_r_bypass_regNext_24_3_df_is_ws_13;
  reg                 io_in_r_bypass_regNext_24_3_stall_13;
  reg        [15:0]   io_in_r_bypass_regNext_25_0_data_13;
  reg                 io_in_r_bypass_regNext_25_0_load_store_13;
  reg                 io_in_r_bypass_regNext_25_0_df_is_ws_13;
  reg                 io_in_r_bypass_regNext_25_0_stall_13;
  reg        [15:0]   io_in_r_bypass_regNext_25_1_data_13;
  reg                 io_in_r_bypass_regNext_25_1_load_store_13;
  reg                 io_in_r_bypass_regNext_25_1_df_is_ws_13;
  reg                 io_in_r_bypass_regNext_25_1_stall_13;
  reg        [15:0]   io_in_r_bypass_regNext_25_2_data_13;
  reg                 io_in_r_bypass_regNext_25_2_load_store_13;
  reg                 io_in_r_bypass_regNext_25_2_df_is_ws_13;
  reg                 io_in_r_bypass_regNext_25_2_stall_13;
  reg        [15:0]   io_in_r_bypass_regNext_25_3_data_13;
  reg                 io_in_r_bypass_regNext_25_3_load_store_13;
  reg                 io_in_r_bypass_regNext_25_3_df_is_ws_13;
  reg                 io_in_r_bypass_regNext_25_3_stall_13;
  reg        [15:0]   io_in_r_bypass_regNext_26_0_data_13;
  reg                 io_in_r_bypass_regNext_26_0_load_store_13;
  reg                 io_in_r_bypass_regNext_26_0_df_is_ws_13;
  reg                 io_in_r_bypass_regNext_26_0_stall_13;
  reg        [15:0]   io_in_r_bypass_regNext_26_1_data_13;
  reg                 io_in_r_bypass_regNext_26_1_load_store_13;
  reg                 io_in_r_bypass_regNext_26_1_df_is_ws_13;
  reg                 io_in_r_bypass_regNext_26_1_stall_13;
  reg        [15:0]   io_in_r_bypass_regNext_26_2_data_13;
  reg                 io_in_r_bypass_regNext_26_2_load_store_13;
  reg                 io_in_r_bypass_regNext_26_2_df_is_ws_13;
  reg                 io_in_r_bypass_regNext_26_2_stall_13;
  reg        [15:0]   io_in_r_bypass_regNext_26_3_data_13;
  reg                 io_in_r_bypass_regNext_26_3_load_store_13;
  reg                 io_in_r_bypass_regNext_26_3_df_is_ws_13;
  reg                 io_in_r_bypass_regNext_26_3_stall_13;
  reg        [15:0]   io_in_r_bypass_regNext_27_0_data_13;
  reg                 io_in_r_bypass_regNext_27_0_load_store_13;
  reg                 io_in_r_bypass_regNext_27_0_df_is_ws_13;
  reg                 io_in_r_bypass_regNext_27_0_stall_13;
  reg        [15:0]   io_in_r_bypass_regNext_27_1_data_13;
  reg                 io_in_r_bypass_regNext_27_1_load_store_13;
  reg                 io_in_r_bypass_regNext_27_1_df_is_ws_13;
  reg                 io_in_r_bypass_regNext_27_1_stall_13;
  reg        [15:0]   io_in_r_bypass_regNext_27_2_data_13;
  reg                 io_in_r_bypass_regNext_27_2_load_store_13;
  reg                 io_in_r_bypass_regNext_27_2_df_is_ws_13;
  reg                 io_in_r_bypass_regNext_27_2_stall_13;
  reg        [15:0]   io_in_r_bypass_regNext_27_3_data_13;
  reg                 io_in_r_bypass_regNext_27_3_load_store_13;
  reg                 io_in_r_bypass_regNext_27_3_df_is_ws_13;
  reg                 io_in_r_bypass_regNext_27_3_stall_13;
  reg        [15:0]   io_in_r_bypass_regNext_28_0_data_13;
  reg                 io_in_r_bypass_regNext_28_0_load_store_13;
  reg                 io_in_r_bypass_regNext_28_0_df_is_ws_13;
  reg                 io_in_r_bypass_regNext_28_0_stall_13;
  reg        [15:0]   io_in_r_bypass_regNext_28_1_data_13;
  reg                 io_in_r_bypass_regNext_28_1_load_store_13;
  reg                 io_in_r_bypass_regNext_28_1_df_is_ws_13;
  reg                 io_in_r_bypass_regNext_28_1_stall_13;
  reg        [15:0]   io_in_r_bypass_regNext_28_2_data_13;
  reg                 io_in_r_bypass_regNext_28_2_load_store_13;
  reg                 io_in_r_bypass_regNext_28_2_df_is_ws_13;
  reg                 io_in_r_bypass_regNext_28_2_stall_13;
  reg        [15:0]   io_in_r_bypass_regNext_28_3_data_13;
  reg                 io_in_r_bypass_regNext_28_3_load_store_13;
  reg                 io_in_r_bypass_regNext_28_3_df_is_ws_13;
  reg                 io_in_r_bypass_regNext_28_3_stall_13;
  reg        [15:0]   io_in_r_bypass_regNext_29_0_data_13;
  reg                 io_in_r_bypass_regNext_29_0_load_store_13;
  reg                 io_in_r_bypass_regNext_29_0_df_is_ws_13;
  reg                 io_in_r_bypass_regNext_29_0_stall_13;
  reg        [15:0]   io_in_r_bypass_regNext_29_1_data_13;
  reg                 io_in_r_bypass_regNext_29_1_load_store_13;
  reg                 io_in_r_bypass_regNext_29_1_df_is_ws_13;
  reg                 io_in_r_bypass_regNext_29_1_stall_13;
  reg        [15:0]   io_in_r_bypass_regNext_29_2_data_13;
  reg                 io_in_r_bypass_regNext_29_2_load_store_13;
  reg                 io_in_r_bypass_regNext_29_2_df_is_ws_13;
  reg                 io_in_r_bypass_regNext_29_2_stall_13;
  reg        [15:0]   io_in_r_bypass_regNext_29_3_data_13;
  reg                 io_in_r_bypass_regNext_29_3_load_store_13;
  reg                 io_in_r_bypass_regNext_29_3_df_is_ws_13;
  reg                 io_in_r_bypass_regNext_29_3_stall_13;
  reg        [15:0]   io_in_r_bypass_regNext_30_0_data_13;
  reg                 io_in_r_bypass_regNext_30_0_load_store_13;
  reg                 io_in_r_bypass_regNext_30_0_df_is_ws_13;
  reg                 io_in_r_bypass_regNext_30_0_stall_13;
  reg        [15:0]   io_in_r_bypass_regNext_30_1_data_13;
  reg                 io_in_r_bypass_regNext_30_1_load_store_13;
  reg                 io_in_r_bypass_regNext_30_1_df_is_ws_13;
  reg                 io_in_r_bypass_regNext_30_1_stall_13;
  reg        [15:0]   io_in_r_bypass_regNext_30_2_data_13;
  reg                 io_in_r_bypass_regNext_30_2_load_store_13;
  reg                 io_in_r_bypass_regNext_30_2_df_is_ws_13;
  reg                 io_in_r_bypass_regNext_30_2_stall_13;
  reg        [15:0]   io_in_r_bypass_regNext_30_3_data_13;
  reg                 io_in_r_bypass_regNext_30_3_load_store_13;
  reg                 io_in_r_bypass_regNext_30_3_df_is_ws_13;
  reg                 io_in_r_bypass_regNext_30_3_stall_13;
  reg        [15:0]   io_in_r_bypass_regNext_31_0_data_13;
  reg                 io_in_r_bypass_regNext_31_0_load_store_13;
  reg                 io_in_r_bypass_regNext_31_0_df_is_ws_13;
  reg                 io_in_r_bypass_regNext_31_0_stall_13;
  reg        [15:0]   io_in_r_bypass_regNext_31_1_data_13;
  reg                 io_in_r_bypass_regNext_31_1_load_store_13;
  reg                 io_in_r_bypass_regNext_31_1_df_is_ws_13;
  reg                 io_in_r_bypass_regNext_31_1_stall_13;
  reg        [15:0]   io_in_r_bypass_regNext_31_2_data_13;
  reg                 io_in_r_bypass_regNext_31_2_load_store_13;
  reg                 io_in_r_bypass_regNext_31_2_df_is_ws_13;
  reg                 io_in_r_bypass_regNext_31_2_stall_13;
  reg        [15:0]   io_in_r_bypass_regNext_31_3_data_13;
  reg                 io_in_r_bypass_regNext_31_3_load_store_13;
  reg                 io_in_r_bypass_regNext_31_3_df_is_ws_13;
  reg                 io_in_r_bypass_regNext_31_3_stall_13;
  reg        [15:0]   io_in_r_bypass_regNext_0_0_data_14;
  reg                 io_in_r_bypass_regNext_0_0_load_store_14;
  reg                 io_in_r_bypass_regNext_0_0_df_is_ws_14;
  reg                 io_in_r_bypass_regNext_0_0_stall_14;
  reg        [15:0]   io_in_r_bypass_regNext_0_1_data_14;
  reg                 io_in_r_bypass_regNext_0_1_load_store_14;
  reg                 io_in_r_bypass_regNext_0_1_df_is_ws_14;
  reg                 io_in_r_bypass_regNext_0_1_stall_14;
  reg        [15:0]   io_in_r_bypass_regNext_0_2_data_14;
  reg                 io_in_r_bypass_regNext_0_2_load_store_14;
  reg                 io_in_r_bypass_regNext_0_2_df_is_ws_14;
  reg                 io_in_r_bypass_regNext_0_2_stall_14;
  reg        [15:0]   io_in_r_bypass_regNext_0_3_data_14;
  reg                 io_in_r_bypass_regNext_0_3_load_store_14;
  reg                 io_in_r_bypass_regNext_0_3_df_is_ws_14;
  reg                 io_in_r_bypass_regNext_0_3_stall_14;
  reg        [15:0]   io_in_r_bypass_regNext_1_0_data_14;
  reg                 io_in_r_bypass_regNext_1_0_load_store_14;
  reg                 io_in_r_bypass_regNext_1_0_df_is_ws_14;
  reg                 io_in_r_bypass_regNext_1_0_stall_14;
  reg        [15:0]   io_in_r_bypass_regNext_1_1_data_14;
  reg                 io_in_r_bypass_regNext_1_1_load_store_14;
  reg                 io_in_r_bypass_regNext_1_1_df_is_ws_14;
  reg                 io_in_r_bypass_regNext_1_1_stall_14;
  reg        [15:0]   io_in_r_bypass_regNext_1_2_data_14;
  reg                 io_in_r_bypass_regNext_1_2_load_store_14;
  reg                 io_in_r_bypass_regNext_1_2_df_is_ws_14;
  reg                 io_in_r_bypass_regNext_1_2_stall_14;
  reg        [15:0]   io_in_r_bypass_regNext_1_3_data_14;
  reg                 io_in_r_bypass_regNext_1_3_load_store_14;
  reg                 io_in_r_bypass_regNext_1_3_df_is_ws_14;
  reg                 io_in_r_bypass_regNext_1_3_stall_14;
  reg        [15:0]   io_in_r_bypass_regNext_2_0_data_14;
  reg                 io_in_r_bypass_regNext_2_0_load_store_14;
  reg                 io_in_r_bypass_regNext_2_0_df_is_ws_14;
  reg                 io_in_r_bypass_regNext_2_0_stall_14;
  reg        [15:0]   io_in_r_bypass_regNext_2_1_data_14;
  reg                 io_in_r_bypass_regNext_2_1_load_store_14;
  reg                 io_in_r_bypass_regNext_2_1_df_is_ws_14;
  reg                 io_in_r_bypass_regNext_2_1_stall_14;
  reg        [15:0]   io_in_r_bypass_regNext_2_2_data_14;
  reg                 io_in_r_bypass_regNext_2_2_load_store_14;
  reg                 io_in_r_bypass_regNext_2_2_df_is_ws_14;
  reg                 io_in_r_bypass_regNext_2_2_stall_14;
  reg        [15:0]   io_in_r_bypass_regNext_2_3_data_14;
  reg                 io_in_r_bypass_regNext_2_3_load_store_14;
  reg                 io_in_r_bypass_regNext_2_3_df_is_ws_14;
  reg                 io_in_r_bypass_regNext_2_3_stall_14;
  reg        [15:0]   io_in_r_bypass_regNext_3_0_data_14;
  reg                 io_in_r_bypass_regNext_3_0_load_store_14;
  reg                 io_in_r_bypass_regNext_3_0_df_is_ws_14;
  reg                 io_in_r_bypass_regNext_3_0_stall_14;
  reg        [15:0]   io_in_r_bypass_regNext_3_1_data_14;
  reg                 io_in_r_bypass_regNext_3_1_load_store_14;
  reg                 io_in_r_bypass_regNext_3_1_df_is_ws_14;
  reg                 io_in_r_bypass_regNext_3_1_stall_14;
  reg        [15:0]   io_in_r_bypass_regNext_3_2_data_14;
  reg                 io_in_r_bypass_regNext_3_2_load_store_14;
  reg                 io_in_r_bypass_regNext_3_2_df_is_ws_14;
  reg                 io_in_r_bypass_regNext_3_2_stall_14;
  reg        [15:0]   io_in_r_bypass_regNext_3_3_data_14;
  reg                 io_in_r_bypass_regNext_3_3_load_store_14;
  reg                 io_in_r_bypass_regNext_3_3_df_is_ws_14;
  reg                 io_in_r_bypass_regNext_3_3_stall_14;
  reg        [15:0]   io_in_r_bypass_regNext_4_0_data_14;
  reg                 io_in_r_bypass_regNext_4_0_load_store_14;
  reg                 io_in_r_bypass_regNext_4_0_df_is_ws_14;
  reg                 io_in_r_bypass_regNext_4_0_stall_14;
  reg        [15:0]   io_in_r_bypass_regNext_4_1_data_14;
  reg                 io_in_r_bypass_regNext_4_1_load_store_14;
  reg                 io_in_r_bypass_regNext_4_1_df_is_ws_14;
  reg                 io_in_r_bypass_regNext_4_1_stall_14;
  reg        [15:0]   io_in_r_bypass_regNext_4_2_data_14;
  reg                 io_in_r_bypass_regNext_4_2_load_store_14;
  reg                 io_in_r_bypass_regNext_4_2_df_is_ws_14;
  reg                 io_in_r_bypass_regNext_4_2_stall_14;
  reg        [15:0]   io_in_r_bypass_regNext_4_3_data_14;
  reg                 io_in_r_bypass_regNext_4_3_load_store_14;
  reg                 io_in_r_bypass_regNext_4_3_df_is_ws_14;
  reg                 io_in_r_bypass_regNext_4_3_stall_14;
  reg        [15:0]   io_in_r_bypass_regNext_5_0_data_14;
  reg                 io_in_r_bypass_regNext_5_0_load_store_14;
  reg                 io_in_r_bypass_regNext_5_0_df_is_ws_14;
  reg                 io_in_r_bypass_regNext_5_0_stall_14;
  reg        [15:0]   io_in_r_bypass_regNext_5_1_data_14;
  reg                 io_in_r_bypass_regNext_5_1_load_store_14;
  reg                 io_in_r_bypass_regNext_5_1_df_is_ws_14;
  reg                 io_in_r_bypass_regNext_5_1_stall_14;
  reg        [15:0]   io_in_r_bypass_regNext_5_2_data_14;
  reg                 io_in_r_bypass_regNext_5_2_load_store_14;
  reg                 io_in_r_bypass_regNext_5_2_df_is_ws_14;
  reg                 io_in_r_bypass_regNext_5_2_stall_14;
  reg        [15:0]   io_in_r_bypass_regNext_5_3_data_14;
  reg                 io_in_r_bypass_regNext_5_3_load_store_14;
  reg                 io_in_r_bypass_regNext_5_3_df_is_ws_14;
  reg                 io_in_r_bypass_regNext_5_3_stall_14;
  reg        [15:0]   io_in_r_bypass_regNext_6_0_data_14;
  reg                 io_in_r_bypass_regNext_6_0_load_store_14;
  reg                 io_in_r_bypass_regNext_6_0_df_is_ws_14;
  reg                 io_in_r_bypass_regNext_6_0_stall_14;
  reg        [15:0]   io_in_r_bypass_regNext_6_1_data_14;
  reg                 io_in_r_bypass_regNext_6_1_load_store_14;
  reg                 io_in_r_bypass_regNext_6_1_df_is_ws_14;
  reg                 io_in_r_bypass_regNext_6_1_stall_14;
  reg        [15:0]   io_in_r_bypass_regNext_6_2_data_14;
  reg                 io_in_r_bypass_regNext_6_2_load_store_14;
  reg                 io_in_r_bypass_regNext_6_2_df_is_ws_14;
  reg                 io_in_r_bypass_regNext_6_2_stall_14;
  reg        [15:0]   io_in_r_bypass_regNext_6_3_data_14;
  reg                 io_in_r_bypass_regNext_6_3_load_store_14;
  reg                 io_in_r_bypass_regNext_6_3_df_is_ws_14;
  reg                 io_in_r_bypass_regNext_6_3_stall_14;
  reg        [15:0]   io_in_r_bypass_regNext_7_0_data_14;
  reg                 io_in_r_bypass_regNext_7_0_load_store_14;
  reg                 io_in_r_bypass_regNext_7_0_df_is_ws_14;
  reg                 io_in_r_bypass_regNext_7_0_stall_14;
  reg        [15:0]   io_in_r_bypass_regNext_7_1_data_14;
  reg                 io_in_r_bypass_regNext_7_1_load_store_14;
  reg                 io_in_r_bypass_regNext_7_1_df_is_ws_14;
  reg                 io_in_r_bypass_regNext_7_1_stall_14;
  reg        [15:0]   io_in_r_bypass_regNext_7_2_data_14;
  reg                 io_in_r_bypass_regNext_7_2_load_store_14;
  reg                 io_in_r_bypass_regNext_7_2_df_is_ws_14;
  reg                 io_in_r_bypass_regNext_7_2_stall_14;
  reg        [15:0]   io_in_r_bypass_regNext_7_3_data_14;
  reg                 io_in_r_bypass_regNext_7_3_load_store_14;
  reg                 io_in_r_bypass_regNext_7_3_df_is_ws_14;
  reg                 io_in_r_bypass_regNext_7_3_stall_14;
  reg        [15:0]   io_in_r_bypass_regNext_8_0_data_14;
  reg                 io_in_r_bypass_regNext_8_0_load_store_14;
  reg                 io_in_r_bypass_regNext_8_0_df_is_ws_14;
  reg                 io_in_r_bypass_regNext_8_0_stall_14;
  reg        [15:0]   io_in_r_bypass_regNext_8_1_data_14;
  reg                 io_in_r_bypass_regNext_8_1_load_store_14;
  reg                 io_in_r_bypass_regNext_8_1_df_is_ws_14;
  reg                 io_in_r_bypass_regNext_8_1_stall_14;
  reg        [15:0]   io_in_r_bypass_regNext_8_2_data_14;
  reg                 io_in_r_bypass_regNext_8_2_load_store_14;
  reg                 io_in_r_bypass_regNext_8_2_df_is_ws_14;
  reg                 io_in_r_bypass_regNext_8_2_stall_14;
  reg        [15:0]   io_in_r_bypass_regNext_8_3_data_14;
  reg                 io_in_r_bypass_regNext_8_3_load_store_14;
  reg                 io_in_r_bypass_regNext_8_3_df_is_ws_14;
  reg                 io_in_r_bypass_regNext_8_3_stall_14;
  reg        [15:0]   io_in_r_bypass_regNext_9_0_data_14;
  reg                 io_in_r_bypass_regNext_9_0_load_store_14;
  reg                 io_in_r_bypass_regNext_9_0_df_is_ws_14;
  reg                 io_in_r_bypass_regNext_9_0_stall_14;
  reg        [15:0]   io_in_r_bypass_regNext_9_1_data_14;
  reg                 io_in_r_bypass_regNext_9_1_load_store_14;
  reg                 io_in_r_bypass_regNext_9_1_df_is_ws_14;
  reg                 io_in_r_bypass_regNext_9_1_stall_14;
  reg        [15:0]   io_in_r_bypass_regNext_9_2_data_14;
  reg                 io_in_r_bypass_regNext_9_2_load_store_14;
  reg                 io_in_r_bypass_regNext_9_2_df_is_ws_14;
  reg                 io_in_r_bypass_regNext_9_2_stall_14;
  reg        [15:0]   io_in_r_bypass_regNext_9_3_data_14;
  reg                 io_in_r_bypass_regNext_9_3_load_store_14;
  reg                 io_in_r_bypass_regNext_9_3_df_is_ws_14;
  reg                 io_in_r_bypass_regNext_9_3_stall_14;
  reg        [15:0]   io_in_r_bypass_regNext_10_0_data_14;
  reg                 io_in_r_bypass_regNext_10_0_load_store_14;
  reg                 io_in_r_bypass_regNext_10_0_df_is_ws_14;
  reg                 io_in_r_bypass_regNext_10_0_stall_14;
  reg        [15:0]   io_in_r_bypass_regNext_10_1_data_14;
  reg                 io_in_r_bypass_regNext_10_1_load_store_14;
  reg                 io_in_r_bypass_regNext_10_1_df_is_ws_14;
  reg                 io_in_r_bypass_regNext_10_1_stall_14;
  reg        [15:0]   io_in_r_bypass_regNext_10_2_data_14;
  reg                 io_in_r_bypass_regNext_10_2_load_store_14;
  reg                 io_in_r_bypass_regNext_10_2_df_is_ws_14;
  reg                 io_in_r_bypass_regNext_10_2_stall_14;
  reg        [15:0]   io_in_r_bypass_regNext_10_3_data_14;
  reg                 io_in_r_bypass_regNext_10_3_load_store_14;
  reg                 io_in_r_bypass_regNext_10_3_df_is_ws_14;
  reg                 io_in_r_bypass_regNext_10_3_stall_14;
  reg        [15:0]   io_in_r_bypass_regNext_11_0_data_14;
  reg                 io_in_r_bypass_regNext_11_0_load_store_14;
  reg                 io_in_r_bypass_regNext_11_0_df_is_ws_14;
  reg                 io_in_r_bypass_regNext_11_0_stall_14;
  reg        [15:0]   io_in_r_bypass_regNext_11_1_data_14;
  reg                 io_in_r_bypass_regNext_11_1_load_store_14;
  reg                 io_in_r_bypass_regNext_11_1_df_is_ws_14;
  reg                 io_in_r_bypass_regNext_11_1_stall_14;
  reg        [15:0]   io_in_r_bypass_regNext_11_2_data_14;
  reg                 io_in_r_bypass_regNext_11_2_load_store_14;
  reg                 io_in_r_bypass_regNext_11_2_df_is_ws_14;
  reg                 io_in_r_bypass_regNext_11_2_stall_14;
  reg        [15:0]   io_in_r_bypass_regNext_11_3_data_14;
  reg                 io_in_r_bypass_regNext_11_3_load_store_14;
  reg                 io_in_r_bypass_regNext_11_3_df_is_ws_14;
  reg                 io_in_r_bypass_regNext_11_3_stall_14;
  reg        [15:0]   io_in_r_bypass_regNext_12_0_data_14;
  reg                 io_in_r_bypass_regNext_12_0_load_store_14;
  reg                 io_in_r_bypass_regNext_12_0_df_is_ws_14;
  reg                 io_in_r_bypass_regNext_12_0_stall_14;
  reg        [15:0]   io_in_r_bypass_regNext_12_1_data_14;
  reg                 io_in_r_bypass_regNext_12_1_load_store_14;
  reg                 io_in_r_bypass_regNext_12_1_df_is_ws_14;
  reg                 io_in_r_bypass_regNext_12_1_stall_14;
  reg        [15:0]   io_in_r_bypass_regNext_12_2_data_14;
  reg                 io_in_r_bypass_regNext_12_2_load_store_14;
  reg                 io_in_r_bypass_regNext_12_2_df_is_ws_14;
  reg                 io_in_r_bypass_regNext_12_2_stall_14;
  reg        [15:0]   io_in_r_bypass_regNext_12_3_data_14;
  reg                 io_in_r_bypass_regNext_12_3_load_store_14;
  reg                 io_in_r_bypass_regNext_12_3_df_is_ws_14;
  reg                 io_in_r_bypass_regNext_12_3_stall_14;
  reg        [15:0]   io_in_r_bypass_regNext_13_0_data_14;
  reg                 io_in_r_bypass_regNext_13_0_load_store_14;
  reg                 io_in_r_bypass_regNext_13_0_df_is_ws_14;
  reg                 io_in_r_bypass_regNext_13_0_stall_14;
  reg        [15:0]   io_in_r_bypass_regNext_13_1_data_14;
  reg                 io_in_r_bypass_regNext_13_1_load_store_14;
  reg                 io_in_r_bypass_regNext_13_1_df_is_ws_14;
  reg                 io_in_r_bypass_regNext_13_1_stall_14;
  reg        [15:0]   io_in_r_bypass_regNext_13_2_data_14;
  reg                 io_in_r_bypass_regNext_13_2_load_store_14;
  reg                 io_in_r_bypass_regNext_13_2_df_is_ws_14;
  reg                 io_in_r_bypass_regNext_13_2_stall_14;
  reg        [15:0]   io_in_r_bypass_regNext_13_3_data_14;
  reg                 io_in_r_bypass_regNext_13_3_load_store_14;
  reg                 io_in_r_bypass_regNext_13_3_df_is_ws_14;
  reg                 io_in_r_bypass_regNext_13_3_stall_14;
  reg        [15:0]   io_in_r_bypass_regNext_14_0_data_14;
  reg                 io_in_r_bypass_regNext_14_0_load_store_14;
  reg                 io_in_r_bypass_regNext_14_0_df_is_ws_14;
  reg                 io_in_r_bypass_regNext_14_0_stall_14;
  reg        [15:0]   io_in_r_bypass_regNext_14_1_data_14;
  reg                 io_in_r_bypass_regNext_14_1_load_store_14;
  reg                 io_in_r_bypass_regNext_14_1_df_is_ws_14;
  reg                 io_in_r_bypass_regNext_14_1_stall_14;
  reg        [15:0]   io_in_r_bypass_regNext_14_2_data_14;
  reg                 io_in_r_bypass_regNext_14_2_load_store_14;
  reg                 io_in_r_bypass_regNext_14_2_df_is_ws_14;
  reg                 io_in_r_bypass_regNext_14_2_stall_14;
  reg        [15:0]   io_in_r_bypass_regNext_14_3_data_14;
  reg                 io_in_r_bypass_regNext_14_3_load_store_14;
  reg                 io_in_r_bypass_regNext_14_3_df_is_ws_14;
  reg                 io_in_r_bypass_regNext_14_3_stall_14;
  reg        [15:0]   io_in_r_bypass_regNext_15_0_data_14;
  reg                 io_in_r_bypass_regNext_15_0_load_store_14;
  reg                 io_in_r_bypass_regNext_15_0_df_is_ws_14;
  reg                 io_in_r_bypass_regNext_15_0_stall_14;
  reg        [15:0]   io_in_r_bypass_regNext_15_1_data_14;
  reg                 io_in_r_bypass_regNext_15_1_load_store_14;
  reg                 io_in_r_bypass_regNext_15_1_df_is_ws_14;
  reg                 io_in_r_bypass_regNext_15_1_stall_14;
  reg        [15:0]   io_in_r_bypass_regNext_15_2_data_14;
  reg                 io_in_r_bypass_regNext_15_2_load_store_14;
  reg                 io_in_r_bypass_regNext_15_2_df_is_ws_14;
  reg                 io_in_r_bypass_regNext_15_2_stall_14;
  reg        [15:0]   io_in_r_bypass_regNext_15_3_data_14;
  reg                 io_in_r_bypass_regNext_15_3_load_store_14;
  reg                 io_in_r_bypass_regNext_15_3_df_is_ws_14;
  reg                 io_in_r_bypass_regNext_15_3_stall_14;
  reg        [15:0]   io_in_r_bypass_regNext_16_0_data_14;
  reg                 io_in_r_bypass_regNext_16_0_load_store_14;
  reg                 io_in_r_bypass_regNext_16_0_df_is_ws_14;
  reg                 io_in_r_bypass_regNext_16_0_stall_14;
  reg        [15:0]   io_in_r_bypass_regNext_16_1_data_14;
  reg                 io_in_r_bypass_regNext_16_1_load_store_14;
  reg                 io_in_r_bypass_regNext_16_1_df_is_ws_14;
  reg                 io_in_r_bypass_regNext_16_1_stall_14;
  reg        [15:0]   io_in_r_bypass_regNext_16_2_data_14;
  reg                 io_in_r_bypass_regNext_16_2_load_store_14;
  reg                 io_in_r_bypass_regNext_16_2_df_is_ws_14;
  reg                 io_in_r_bypass_regNext_16_2_stall_14;
  reg        [15:0]   io_in_r_bypass_regNext_16_3_data_14;
  reg                 io_in_r_bypass_regNext_16_3_load_store_14;
  reg                 io_in_r_bypass_regNext_16_3_df_is_ws_14;
  reg                 io_in_r_bypass_regNext_16_3_stall_14;
  reg        [15:0]   io_in_r_bypass_regNext_17_0_data_14;
  reg                 io_in_r_bypass_regNext_17_0_load_store_14;
  reg                 io_in_r_bypass_regNext_17_0_df_is_ws_14;
  reg                 io_in_r_bypass_regNext_17_0_stall_14;
  reg        [15:0]   io_in_r_bypass_regNext_17_1_data_14;
  reg                 io_in_r_bypass_regNext_17_1_load_store_14;
  reg                 io_in_r_bypass_regNext_17_1_df_is_ws_14;
  reg                 io_in_r_bypass_regNext_17_1_stall_14;
  reg        [15:0]   io_in_r_bypass_regNext_17_2_data_14;
  reg                 io_in_r_bypass_regNext_17_2_load_store_14;
  reg                 io_in_r_bypass_regNext_17_2_df_is_ws_14;
  reg                 io_in_r_bypass_regNext_17_2_stall_14;
  reg        [15:0]   io_in_r_bypass_regNext_17_3_data_14;
  reg                 io_in_r_bypass_regNext_17_3_load_store_14;
  reg                 io_in_r_bypass_regNext_17_3_df_is_ws_14;
  reg                 io_in_r_bypass_regNext_17_3_stall_14;
  reg        [15:0]   io_in_r_bypass_regNext_18_0_data_14;
  reg                 io_in_r_bypass_regNext_18_0_load_store_14;
  reg                 io_in_r_bypass_regNext_18_0_df_is_ws_14;
  reg                 io_in_r_bypass_regNext_18_0_stall_14;
  reg        [15:0]   io_in_r_bypass_regNext_18_1_data_14;
  reg                 io_in_r_bypass_regNext_18_1_load_store_14;
  reg                 io_in_r_bypass_regNext_18_1_df_is_ws_14;
  reg                 io_in_r_bypass_regNext_18_1_stall_14;
  reg        [15:0]   io_in_r_bypass_regNext_18_2_data_14;
  reg                 io_in_r_bypass_regNext_18_2_load_store_14;
  reg                 io_in_r_bypass_regNext_18_2_df_is_ws_14;
  reg                 io_in_r_bypass_regNext_18_2_stall_14;
  reg        [15:0]   io_in_r_bypass_regNext_18_3_data_14;
  reg                 io_in_r_bypass_regNext_18_3_load_store_14;
  reg                 io_in_r_bypass_regNext_18_3_df_is_ws_14;
  reg                 io_in_r_bypass_regNext_18_3_stall_14;
  reg        [15:0]   io_in_r_bypass_regNext_19_0_data_14;
  reg                 io_in_r_bypass_regNext_19_0_load_store_14;
  reg                 io_in_r_bypass_regNext_19_0_df_is_ws_14;
  reg                 io_in_r_bypass_regNext_19_0_stall_14;
  reg        [15:0]   io_in_r_bypass_regNext_19_1_data_14;
  reg                 io_in_r_bypass_regNext_19_1_load_store_14;
  reg                 io_in_r_bypass_regNext_19_1_df_is_ws_14;
  reg                 io_in_r_bypass_regNext_19_1_stall_14;
  reg        [15:0]   io_in_r_bypass_regNext_19_2_data_14;
  reg                 io_in_r_bypass_regNext_19_2_load_store_14;
  reg                 io_in_r_bypass_regNext_19_2_df_is_ws_14;
  reg                 io_in_r_bypass_regNext_19_2_stall_14;
  reg        [15:0]   io_in_r_bypass_regNext_19_3_data_14;
  reg                 io_in_r_bypass_regNext_19_3_load_store_14;
  reg                 io_in_r_bypass_regNext_19_3_df_is_ws_14;
  reg                 io_in_r_bypass_regNext_19_3_stall_14;
  reg        [15:0]   io_in_r_bypass_regNext_20_0_data_14;
  reg                 io_in_r_bypass_regNext_20_0_load_store_14;
  reg                 io_in_r_bypass_regNext_20_0_df_is_ws_14;
  reg                 io_in_r_bypass_regNext_20_0_stall_14;
  reg        [15:0]   io_in_r_bypass_regNext_20_1_data_14;
  reg                 io_in_r_bypass_regNext_20_1_load_store_14;
  reg                 io_in_r_bypass_regNext_20_1_df_is_ws_14;
  reg                 io_in_r_bypass_regNext_20_1_stall_14;
  reg        [15:0]   io_in_r_bypass_regNext_20_2_data_14;
  reg                 io_in_r_bypass_regNext_20_2_load_store_14;
  reg                 io_in_r_bypass_regNext_20_2_df_is_ws_14;
  reg                 io_in_r_bypass_regNext_20_2_stall_14;
  reg        [15:0]   io_in_r_bypass_regNext_20_3_data_14;
  reg                 io_in_r_bypass_regNext_20_3_load_store_14;
  reg                 io_in_r_bypass_regNext_20_3_df_is_ws_14;
  reg                 io_in_r_bypass_regNext_20_3_stall_14;
  reg        [15:0]   io_in_r_bypass_regNext_21_0_data_14;
  reg                 io_in_r_bypass_regNext_21_0_load_store_14;
  reg                 io_in_r_bypass_regNext_21_0_df_is_ws_14;
  reg                 io_in_r_bypass_regNext_21_0_stall_14;
  reg        [15:0]   io_in_r_bypass_regNext_21_1_data_14;
  reg                 io_in_r_bypass_regNext_21_1_load_store_14;
  reg                 io_in_r_bypass_regNext_21_1_df_is_ws_14;
  reg                 io_in_r_bypass_regNext_21_1_stall_14;
  reg        [15:0]   io_in_r_bypass_regNext_21_2_data_14;
  reg                 io_in_r_bypass_regNext_21_2_load_store_14;
  reg                 io_in_r_bypass_regNext_21_2_df_is_ws_14;
  reg                 io_in_r_bypass_regNext_21_2_stall_14;
  reg        [15:0]   io_in_r_bypass_regNext_21_3_data_14;
  reg                 io_in_r_bypass_regNext_21_3_load_store_14;
  reg                 io_in_r_bypass_regNext_21_3_df_is_ws_14;
  reg                 io_in_r_bypass_regNext_21_3_stall_14;
  reg        [15:0]   io_in_r_bypass_regNext_22_0_data_14;
  reg                 io_in_r_bypass_regNext_22_0_load_store_14;
  reg                 io_in_r_bypass_regNext_22_0_df_is_ws_14;
  reg                 io_in_r_bypass_regNext_22_0_stall_14;
  reg        [15:0]   io_in_r_bypass_regNext_22_1_data_14;
  reg                 io_in_r_bypass_regNext_22_1_load_store_14;
  reg                 io_in_r_bypass_regNext_22_1_df_is_ws_14;
  reg                 io_in_r_bypass_regNext_22_1_stall_14;
  reg        [15:0]   io_in_r_bypass_regNext_22_2_data_14;
  reg                 io_in_r_bypass_regNext_22_2_load_store_14;
  reg                 io_in_r_bypass_regNext_22_2_df_is_ws_14;
  reg                 io_in_r_bypass_regNext_22_2_stall_14;
  reg        [15:0]   io_in_r_bypass_regNext_22_3_data_14;
  reg                 io_in_r_bypass_regNext_22_3_load_store_14;
  reg                 io_in_r_bypass_regNext_22_3_df_is_ws_14;
  reg                 io_in_r_bypass_regNext_22_3_stall_14;
  reg        [15:0]   io_in_r_bypass_regNext_23_0_data_14;
  reg                 io_in_r_bypass_regNext_23_0_load_store_14;
  reg                 io_in_r_bypass_regNext_23_0_df_is_ws_14;
  reg                 io_in_r_bypass_regNext_23_0_stall_14;
  reg        [15:0]   io_in_r_bypass_regNext_23_1_data_14;
  reg                 io_in_r_bypass_regNext_23_1_load_store_14;
  reg                 io_in_r_bypass_regNext_23_1_df_is_ws_14;
  reg                 io_in_r_bypass_regNext_23_1_stall_14;
  reg        [15:0]   io_in_r_bypass_regNext_23_2_data_14;
  reg                 io_in_r_bypass_regNext_23_2_load_store_14;
  reg                 io_in_r_bypass_regNext_23_2_df_is_ws_14;
  reg                 io_in_r_bypass_regNext_23_2_stall_14;
  reg        [15:0]   io_in_r_bypass_regNext_23_3_data_14;
  reg                 io_in_r_bypass_regNext_23_3_load_store_14;
  reg                 io_in_r_bypass_regNext_23_3_df_is_ws_14;
  reg                 io_in_r_bypass_regNext_23_3_stall_14;
  reg        [15:0]   io_in_r_bypass_regNext_24_0_data_14;
  reg                 io_in_r_bypass_regNext_24_0_load_store_14;
  reg                 io_in_r_bypass_regNext_24_0_df_is_ws_14;
  reg                 io_in_r_bypass_regNext_24_0_stall_14;
  reg        [15:0]   io_in_r_bypass_regNext_24_1_data_14;
  reg                 io_in_r_bypass_regNext_24_1_load_store_14;
  reg                 io_in_r_bypass_regNext_24_1_df_is_ws_14;
  reg                 io_in_r_bypass_regNext_24_1_stall_14;
  reg        [15:0]   io_in_r_bypass_regNext_24_2_data_14;
  reg                 io_in_r_bypass_regNext_24_2_load_store_14;
  reg                 io_in_r_bypass_regNext_24_2_df_is_ws_14;
  reg                 io_in_r_bypass_regNext_24_2_stall_14;
  reg        [15:0]   io_in_r_bypass_regNext_24_3_data_14;
  reg                 io_in_r_bypass_regNext_24_3_load_store_14;
  reg                 io_in_r_bypass_regNext_24_3_df_is_ws_14;
  reg                 io_in_r_bypass_regNext_24_3_stall_14;
  reg        [15:0]   io_in_r_bypass_regNext_25_0_data_14;
  reg                 io_in_r_bypass_regNext_25_0_load_store_14;
  reg                 io_in_r_bypass_regNext_25_0_df_is_ws_14;
  reg                 io_in_r_bypass_regNext_25_0_stall_14;
  reg        [15:0]   io_in_r_bypass_regNext_25_1_data_14;
  reg                 io_in_r_bypass_regNext_25_1_load_store_14;
  reg                 io_in_r_bypass_regNext_25_1_df_is_ws_14;
  reg                 io_in_r_bypass_regNext_25_1_stall_14;
  reg        [15:0]   io_in_r_bypass_regNext_25_2_data_14;
  reg                 io_in_r_bypass_regNext_25_2_load_store_14;
  reg                 io_in_r_bypass_regNext_25_2_df_is_ws_14;
  reg                 io_in_r_bypass_regNext_25_2_stall_14;
  reg        [15:0]   io_in_r_bypass_regNext_25_3_data_14;
  reg                 io_in_r_bypass_regNext_25_3_load_store_14;
  reg                 io_in_r_bypass_regNext_25_3_df_is_ws_14;
  reg                 io_in_r_bypass_regNext_25_3_stall_14;
  reg        [15:0]   io_in_r_bypass_regNext_26_0_data_14;
  reg                 io_in_r_bypass_regNext_26_0_load_store_14;
  reg                 io_in_r_bypass_regNext_26_0_df_is_ws_14;
  reg                 io_in_r_bypass_regNext_26_0_stall_14;
  reg        [15:0]   io_in_r_bypass_regNext_26_1_data_14;
  reg                 io_in_r_bypass_regNext_26_1_load_store_14;
  reg                 io_in_r_bypass_regNext_26_1_df_is_ws_14;
  reg                 io_in_r_bypass_regNext_26_1_stall_14;
  reg        [15:0]   io_in_r_bypass_regNext_26_2_data_14;
  reg                 io_in_r_bypass_regNext_26_2_load_store_14;
  reg                 io_in_r_bypass_regNext_26_2_df_is_ws_14;
  reg                 io_in_r_bypass_regNext_26_2_stall_14;
  reg        [15:0]   io_in_r_bypass_regNext_26_3_data_14;
  reg                 io_in_r_bypass_regNext_26_3_load_store_14;
  reg                 io_in_r_bypass_regNext_26_3_df_is_ws_14;
  reg                 io_in_r_bypass_regNext_26_3_stall_14;
  reg        [15:0]   io_in_r_bypass_regNext_27_0_data_14;
  reg                 io_in_r_bypass_regNext_27_0_load_store_14;
  reg                 io_in_r_bypass_regNext_27_0_df_is_ws_14;
  reg                 io_in_r_bypass_regNext_27_0_stall_14;
  reg        [15:0]   io_in_r_bypass_regNext_27_1_data_14;
  reg                 io_in_r_bypass_regNext_27_1_load_store_14;
  reg                 io_in_r_bypass_regNext_27_1_df_is_ws_14;
  reg                 io_in_r_bypass_regNext_27_1_stall_14;
  reg        [15:0]   io_in_r_bypass_regNext_27_2_data_14;
  reg                 io_in_r_bypass_regNext_27_2_load_store_14;
  reg                 io_in_r_bypass_regNext_27_2_df_is_ws_14;
  reg                 io_in_r_bypass_regNext_27_2_stall_14;
  reg        [15:0]   io_in_r_bypass_regNext_27_3_data_14;
  reg                 io_in_r_bypass_regNext_27_3_load_store_14;
  reg                 io_in_r_bypass_regNext_27_3_df_is_ws_14;
  reg                 io_in_r_bypass_regNext_27_3_stall_14;
  reg        [15:0]   io_in_r_bypass_regNext_28_0_data_14;
  reg                 io_in_r_bypass_regNext_28_0_load_store_14;
  reg                 io_in_r_bypass_regNext_28_0_df_is_ws_14;
  reg                 io_in_r_bypass_regNext_28_0_stall_14;
  reg        [15:0]   io_in_r_bypass_regNext_28_1_data_14;
  reg                 io_in_r_bypass_regNext_28_1_load_store_14;
  reg                 io_in_r_bypass_regNext_28_1_df_is_ws_14;
  reg                 io_in_r_bypass_regNext_28_1_stall_14;
  reg        [15:0]   io_in_r_bypass_regNext_28_2_data_14;
  reg                 io_in_r_bypass_regNext_28_2_load_store_14;
  reg                 io_in_r_bypass_regNext_28_2_df_is_ws_14;
  reg                 io_in_r_bypass_regNext_28_2_stall_14;
  reg        [15:0]   io_in_r_bypass_regNext_28_3_data_14;
  reg                 io_in_r_bypass_regNext_28_3_load_store_14;
  reg                 io_in_r_bypass_regNext_28_3_df_is_ws_14;
  reg                 io_in_r_bypass_regNext_28_3_stall_14;
  reg        [15:0]   io_in_r_bypass_regNext_29_0_data_14;
  reg                 io_in_r_bypass_regNext_29_0_load_store_14;
  reg                 io_in_r_bypass_regNext_29_0_df_is_ws_14;
  reg                 io_in_r_bypass_regNext_29_0_stall_14;
  reg        [15:0]   io_in_r_bypass_regNext_29_1_data_14;
  reg                 io_in_r_bypass_regNext_29_1_load_store_14;
  reg                 io_in_r_bypass_regNext_29_1_df_is_ws_14;
  reg                 io_in_r_bypass_regNext_29_1_stall_14;
  reg        [15:0]   io_in_r_bypass_regNext_29_2_data_14;
  reg                 io_in_r_bypass_regNext_29_2_load_store_14;
  reg                 io_in_r_bypass_regNext_29_2_df_is_ws_14;
  reg                 io_in_r_bypass_regNext_29_2_stall_14;
  reg        [15:0]   io_in_r_bypass_regNext_29_3_data_14;
  reg                 io_in_r_bypass_regNext_29_3_load_store_14;
  reg                 io_in_r_bypass_regNext_29_3_df_is_ws_14;
  reg                 io_in_r_bypass_regNext_29_3_stall_14;
  reg        [15:0]   io_in_r_bypass_regNext_30_0_data_14;
  reg                 io_in_r_bypass_regNext_30_0_load_store_14;
  reg                 io_in_r_bypass_regNext_30_0_df_is_ws_14;
  reg                 io_in_r_bypass_regNext_30_0_stall_14;
  reg        [15:0]   io_in_r_bypass_regNext_30_1_data_14;
  reg                 io_in_r_bypass_regNext_30_1_load_store_14;
  reg                 io_in_r_bypass_regNext_30_1_df_is_ws_14;
  reg                 io_in_r_bypass_regNext_30_1_stall_14;
  reg        [15:0]   io_in_r_bypass_regNext_30_2_data_14;
  reg                 io_in_r_bypass_regNext_30_2_load_store_14;
  reg                 io_in_r_bypass_regNext_30_2_df_is_ws_14;
  reg                 io_in_r_bypass_regNext_30_2_stall_14;
  reg        [15:0]   io_in_r_bypass_regNext_30_3_data_14;
  reg                 io_in_r_bypass_regNext_30_3_load_store_14;
  reg                 io_in_r_bypass_regNext_30_3_df_is_ws_14;
  reg                 io_in_r_bypass_regNext_30_3_stall_14;
  reg        [15:0]   io_in_r_bypass_regNext_31_0_data_14;
  reg                 io_in_r_bypass_regNext_31_0_load_store_14;
  reg                 io_in_r_bypass_regNext_31_0_df_is_ws_14;
  reg                 io_in_r_bypass_regNext_31_0_stall_14;
  reg        [15:0]   io_in_r_bypass_regNext_31_1_data_14;
  reg                 io_in_r_bypass_regNext_31_1_load_store_14;
  reg                 io_in_r_bypass_regNext_31_1_df_is_ws_14;
  reg                 io_in_r_bypass_regNext_31_1_stall_14;
  reg        [15:0]   io_in_r_bypass_regNext_31_2_data_14;
  reg                 io_in_r_bypass_regNext_31_2_load_store_14;
  reg                 io_in_r_bypass_regNext_31_2_df_is_ws_14;
  reg                 io_in_r_bypass_regNext_31_2_stall_14;
  reg        [15:0]   io_in_r_bypass_regNext_31_3_data_14;
  reg                 io_in_r_bypass_regNext_31_3_load_store_14;
  reg                 io_in_r_bypass_regNext_31_3_df_is_ws_14;
  reg                 io_in_r_bypass_regNext_31_3_stall_14;
  reg        [15:0]   io_in_r_bypass_regNext_0_0_data_15;
  reg                 io_in_r_bypass_regNext_0_0_load_store_15;
  reg                 io_in_r_bypass_regNext_0_0_df_is_ws_15;
  reg                 io_in_r_bypass_regNext_0_0_stall_15;
  reg        [15:0]   io_in_r_bypass_regNext_0_1_data_15;
  reg                 io_in_r_bypass_regNext_0_1_load_store_15;
  reg                 io_in_r_bypass_regNext_0_1_df_is_ws_15;
  reg                 io_in_r_bypass_regNext_0_1_stall_15;
  reg        [15:0]   io_in_r_bypass_regNext_0_2_data_15;
  reg                 io_in_r_bypass_regNext_0_2_load_store_15;
  reg                 io_in_r_bypass_regNext_0_2_df_is_ws_15;
  reg                 io_in_r_bypass_regNext_0_2_stall_15;
  reg        [15:0]   io_in_r_bypass_regNext_0_3_data_15;
  reg                 io_in_r_bypass_regNext_0_3_load_store_15;
  reg                 io_in_r_bypass_regNext_0_3_df_is_ws_15;
  reg                 io_in_r_bypass_regNext_0_3_stall_15;
  reg        [15:0]   io_in_r_bypass_regNext_1_0_data_15;
  reg                 io_in_r_bypass_regNext_1_0_load_store_15;
  reg                 io_in_r_bypass_regNext_1_0_df_is_ws_15;
  reg                 io_in_r_bypass_regNext_1_0_stall_15;
  reg        [15:0]   io_in_r_bypass_regNext_1_1_data_15;
  reg                 io_in_r_bypass_regNext_1_1_load_store_15;
  reg                 io_in_r_bypass_regNext_1_1_df_is_ws_15;
  reg                 io_in_r_bypass_regNext_1_1_stall_15;
  reg        [15:0]   io_in_r_bypass_regNext_1_2_data_15;
  reg                 io_in_r_bypass_regNext_1_2_load_store_15;
  reg                 io_in_r_bypass_regNext_1_2_df_is_ws_15;
  reg                 io_in_r_bypass_regNext_1_2_stall_15;
  reg        [15:0]   io_in_r_bypass_regNext_1_3_data_15;
  reg                 io_in_r_bypass_regNext_1_3_load_store_15;
  reg                 io_in_r_bypass_regNext_1_3_df_is_ws_15;
  reg                 io_in_r_bypass_regNext_1_3_stall_15;
  reg        [15:0]   io_in_r_bypass_regNext_2_0_data_15;
  reg                 io_in_r_bypass_regNext_2_0_load_store_15;
  reg                 io_in_r_bypass_regNext_2_0_df_is_ws_15;
  reg                 io_in_r_bypass_regNext_2_0_stall_15;
  reg        [15:0]   io_in_r_bypass_regNext_2_1_data_15;
  reg                 io_in_r_bypass_regNext_2_1_load_store_15;
  reg                 io_in_r_bypass_regNext_2_1_df_is_ws_15;
  reg                 io_in_r_bypass_regNext_2_1_stall_15;
  reg        [15:0]   io_in_r_bypass_regNext_2_2_data_15;
  reg                 io_in_r_bypass_regNext_2_2_load_store_15;
  reg                 io_in_r_bypass_regNext_2_2_df_is_ws_15;
  reg                 io_in_r_bypass_regNext_2_2_stall_15;
  reg        [15:0]   io_in_r_bypass_regNext_2_3_data_15;
  reg                 io_in_r_bypass_regNext_2_3_load_store_15;
  reg                 io_in_r_bypass_regNext_2_3_df_is_ws_15;
  reg                 io_in_r_bypass_regNext_2_3_stall_15;
  reg        [15:0]   io_in_r_bypass_regNext_3_0_data_15;
  reg                 io_in_r_bypass_regNext_3_0_load_store_15;
  reg                 io_in_r_bypass_regNext_3_0_df_is_ws_15;
  reg                 io_in_r_bypass_regNext_3_0_stall_15;
  reg        [15:0]   io_in_r_bypass_regNext_3_1_data_15;
  reg                 io_in_r_bypass_regNext_3_1_load_store_15;
  reg                 io_in_r_bypass_regNext_3_1_df_is_ws_15;
  reg                 io_in_r_bypass_regNext_3_1_stall_15;
  reg        [15:0]   io_in_r_bypass_regNext_3_2_data_15;
  reg                 io_in_r_bypass_regNext_3_2_load_store_15;
  reg                 io_in_r_bypass_regNext_3_2_df_is_ws_15;
  reg                 io_in_r_bypass_regNext_3_2_stall_15;
  reg        [15:0]   io_in_r_bypass_regNext_3_3_data_15;
  reg                 io_in_r_bypass_regNext_3_3_load_store_15;
  reg                 io_in_r_bypass_regNext_3_3_df_is_ws_15;
  reg                 io_in_r_bypass_regNext_3_3_stall_15;
  reg        [15:0]   io_in_r_bypass_regNext_4_0_data_15;
  reg                 io_in_r_bypass_regNext_4_0_load_store_15;
  reg                 io_in_r_bypass_regNext_4_0_df_is_ws_15;
  reg                 io_in_r_bypass_regNext_4_0_stall_15;
  reg        [15:0]   io_in_r_bypass_regNext_4_1_data_15;
  reg                 io_in_r_bypass_regNext_4_1_load_store_15;
  reg                 io_in_r_bypass_regNext_4_1_df_is_ws_15;
  reg                 io_in_r_bypass_regNext_4_1_stall_15;
  reg        [15:0]   io_in_r_bypass_regNext_4_2_data_15;
  reg                 io_in_r_bypass_regNext_4_2_load_store_15;
  reg                 io_in_r_bypass_regNext_4_2_df_is_ws_15;
  reg                 io_in_r_bypass_regNext_4_2_stall_15;
  reg        [15:0]   io_in_r_bypass_regNext_4_3_data_15;
  reg                 io_in_r_bypass_regNext_4_3_load_store_15;
  reg                 io_in_r_bypass_regNext_4_3_df_is_ws_15;
  reg                 io_in_r_bypass_regNext_4_3_stall_15;
  reg        [15:0]   io_in_r_bypass_regNext_5_0_data_15;
  reg                 io_in_r_bypass_regNext_5_0_load_store_15;
  reg                 io_in_r_bypass_regNext_5_0_df_is_ws_15;
  reg                 io_in_r_bypass_regNext_5_0_stall_15;
  reg        [15:0]   io_in_r_bypass_regNext_5_1_data_15;
  reg                 io_in_r_bypass_regNext_5_1_load_store_15;
  reg                 io_in_r_bypass_regNext_5_1_df_is_ws_15;
  reg                 io_in_r_bypass_regNext_5_1_stall_15;
  reg        [15:0]   io_in_r_bypass_regNext_5_2_data_15;
  reg                 io_in_r_bypass_regNext_5_2_load_store_15;
  reg                 io_in_r_bypass_regNext_5_2_df_is_ws_15;
  reg                 io_in_r_bypass_regNext_5_2_stall_15;
  reg        [15:0]   io_in_r_bypass_regNext_5_3_data_15;
  reg                 io_in_r_bypass_regNext_5_3_load_store_15;
  reg                 io_in_r_bypass_regNext_5_3_df_is_ws_15;
  reg                 io_in_r_bypass_regNext_5_3_stall_15;
  reg        [15:0]   io_in_r_bypass_regNext_6_0_data_15;
  reg                 io_in_r_bypass_regNext_6_0_load_store_15;
  reg                 io_in_r_bypass_regNext_6_0_df_is_ws_15;
  reg                 io_in_r_bypass_regNext_6_0_stall_15;
  reg        [15:0]   io_in_r_bypass_regNext_6_1_data_15;
  reg                 io_in_r_bypass_regNext_6_1_load_store_15;
  reg                 io_in_r_bypass_regNext_6_1_df_is_ws_15;
  reg                 io_in_r_bypass_regNext_6_1_stall_15;
  reg        [15:0]   io_in_r_bypass_regNext_6_2_data_15;
  reg                 io_in_r_bypass_regNext_6_2_load_store_15;
  reg                 io_in_r_bypass_regNext_6_2_df_is_ws_15;
  reg                 io_in_r_bypass_regNext_6_2_stall_15;
  reg        [15:0]   io_in_r_bypass_regNext_6_3_data_15;
  reg                 io_in_r_bypass_regNext_6_3_load_store_15;
  reg                 io_in_r_bypass_regNext_6_3_df_is_ws_15;
  reg                 io_in_r_bypass_regNext_6_3_stall_15;
  reg        [15:0]   io_in_r_bypass_regNext_7_0_data_15;
  reg                 io_in_r_bypass_regNext_7_0_load_store_15;
  reg                 io_in_r_bypass_regNext_7_0_df_is_ws_15;
  reg                 io_in_r_bypass_regNext_7_0_stall_15;
  reg        [15:0]   io_in_r_bypass_regNext_7_1_data_15;
  reg                 io_in_r_bypass_regNext_7_1_load_store_15;
  reg                 io_in_r_bypass_regNext_7_1_df_is_ws_15;
  reg                 io_in_r_bypass_regNext_7_1_stall_15;
  reg        [15:0]   io_in_r_bypass_regNext_7_2_data_15;
  reg                 io_in_r_bypass_regNext_7_2_load_store_15;
  reg                 io_in_r_bypass_regNext_7_2_df_is_ws_15;
  reg                 io_in_r_bypass_regNext_7_2_stall_15;
  reg        [15:0]   io_in_r_bypass_regNext_7_3_data_15;
  reg                 io_in_r_bypass_regNext_7_3_load_store_15;
  reg                 io_in_r_bypass_regNext_7_3_df_is_ws_15;
  reg                 io_in_r_bypass_regNext_7_3_stall_15;
  reg        [15:0]   io_in_r_bypass_regNext_8_0_data_15;
  reg                 io_in_r_bypass_regNext_8_0_load_store_15;
  reg                 io_in_r_bypass_regNext_8_0_df_is_ws_15;
  reg                 io_in_r_bypass_regNext_8_0_stall_15;
  reg        [15:0]   io_in_r_bypass_regNext_8_1_data_15;
  reg                 io_in_r_bypass_regNext_8_1_load_store_15;
  reg                 io_in_r_bypass_regNext_8_1_df_is_ws_15;
  reg                 io_in_r_bypass_regNext_8_1_stall_15;
  reg        [15:0]   io_in_r_bypass_regNext_8_2_data_15;
  reg                 io_in_r_bypass_regNext_8_2_load_store_15;
  reg                 io_in_r_bypass_regNext_8_2_df_is_ws_15;
  reg                 io_in_r_bypass_regNext_8_2_stall_15;
  reg        [15:0]   io_in_r_bypass_regNext_8_3_data_15;
  reg                 io_in_r_bypass_regNext_8_3_load_store_15;
  reg                 io_in_r_bypass_regNext_8_3_df_is_ws_15;
  reg                 io_in_r_bypass_regNext_8_3_stall_15;
  reg        [15:0]   io_in_r_bypass_regNext_9_0_data_15;
  reg                 io_in_r_bypass_regNext_9_0_load_store_15;
  reg                 io_in_r_bypass_regNext_9_0_df_is_ws_15;
  reg                 io_in_r_bypass_regNext_9_0_stall_15;
  reg        [15:0]   io_in_r_bypass_regNext_9_1_data_15;
  reg                 io_in_r_bypass_regNext_9_1_load_store_15;
  reg                 io_in_r_bypass_regNext_9_1_df_is_ws_15;
  reg                 io_in_r_bypass_regNext_9_1_stall_15;
  reg        [15:0]   io_in_r_bypass_regNext_9_2_data_15;
  reg                 io_in_r_bypass_regNext_9_2_load_store_15;
  reg                 io_in_r_bypass_regNext_9_2_df_is_ws_15;
  reg                 io_in_r_bypass_regNext_9_2_stall_15;
  reg        [15:0]   io_in_r_bypass_regNext_9_3_data_15;
  reg                 io_in_r_bypass_regNext_9_3_load_store_15;
  reg                 io_in_r_bypass_regNext_9_3_df_is_ws_15;
  reg                 io_in_r_bypass_regNext_9_3_stall_15;
  reg        [15:0]   io_in_r_bypass_regNext_10_0_data_15;
  reg                 io_in_r_bypass_regNext_10_0_load_store_15;
  reg                 io_in_r_bypass_regNext_10_0_df_is_ws_15;
  reg                 io_in_r_bypass_regNext_10_0_stall_15;
  reg        [15:0]   io_in_r_bypass_regNext_10_1_data_15;
  reg                 io_in_r_bypass_regNext_10_1_load_store_15;
  reg                 io_in_r_bypass_regNext_10_1_df_is_ws_15;
  reg                 io_in_r_bypass_regNext_10_1_stall_15;
  reg        [15:0]   io_in_r_bypass_regNext_10_2_data_15;
  reg                 io_in_r_bypass_regNext_10_2_load_store_15;
  reg                 io_in_r_bypass_regNext_10_2_df_is_ws_15;
  reg                 io_in_r_bypass_regNext_10_2_stall_15;
  reg        [15:0]   io_in_r_bypass_regNext_10_3_data_15;
  reg                 io_in_r_bypass_regNext_10_3_load_store_15;
  reg                 io_in_r_bypass_regNext_10_3_df_is_ws_15;
  reg                 io_in_r_bypass_regNext_10_3_stall_15;
  reg        [15:0]   io_in_r_bypass_regNext_11_0_data_15;
  reg                 io_in_r_bypass_regNext_11_0_load_store_15;
  reg                 io_in_r_bypass_regNext_11_0_df_is_ws_15;
  reg                 io_in_r_bypass_regNext_11_0_stall_15;
  reg        [15:0]   io_in_r_bypass_regNext_11_1_data_15;
  reg                 io_in_r_bypass_regNext_11_1_load_store_15;
  reg                 io_in_r_bypass_regNext_11_1_df_is_ws_15;
  reg                 io_in_r_bypass_regNext_11_1_stall_15;
  reg        [15:0]   io_in_r_bypass_regNext_11_2_data_15;
  reg                 io_in_r_bypass_regNext_11_2_load_store_15;
  reg                 io_in_r_bypass_regNext_11_2_df_is_ws_15;
  reg                 io_in_r_bypass_regNext_11_2_stall_15;
  reg        [15:0]   io_in_r_bypass_regNext_11_3_data_15;
  reg                 io_in_r_bypass_regNext_11_3_load_store_15;
  reg                 io_in_r_bypass_regNext_11_3_df_is_ws_15;
  reg                 io_in_r_bypass_regNext_11_3_stall_15;
  reg        [15:0]   io_in_r_bypass_regNext_12_0_data_15;
  reg                 io_in_r_bypass_regNext_12_0_load_store_15;
  reg                 io_in_r_bypass_regNext_12_0_df_is_ws_15;
  reg                 io_in_r_bypass_regNext_12_0_stall_15;
  reg        [15:0]   io_in_r_bypass_regNext_12_1_data_15;
  reg                 io_in_r_bypass_regNext_12_1_load_store_15;
  reg                 io_in_r_bypass_regNext_12_1_df_is_ws_15;
  reg                 io_in_r_bypass_regNext_12_1_stall_15;
  reg        [15:0]   io_in_r_bypass_regNext_12_2_data_15;
  reg                 io_in_r_bypass_regNext_12_2_load_store_15;
  reg                 io_in_r_bypass_regNext_12_2_df_is_ws_15;
  reg                 io_in_r_bypass_regNext_12_2_stall_15;
  reg        [15:0]   io_in_r_bypass_regNext_12_3_data_15;
  reg                 io_in_r_bypass_regNext_12_3_load_store_15;
  reg                 io_in_r_bypass_regNext_12_3_df_is_ws_15;
  reg                 io_in_r_bypass_regNext_12_3_stall_15;
  reg        [15:0]   io_in_r_bypass_regNext_13_0_data_15;
  reg                 io_in_r_bypass_regNext_13_0_load_store_15;
  reg                 io_in_r_bypass_regNext_13_0_df_is_ws_15;
  reg                 io_in_r_bypass_regNext_13_0_stall_15;
  reg        [15:0]   io_in_r_bypass_regNext_13_1_data_15;
  reg                 io_in_r_bypass_regNext_13_1_load_store_15;
  reg                 io_in_r_bypass_regNext_13_1_df_is_ws_15;
  reg                 io_in_r_bypass_regNext_13_1_stall_15;
  reg        [15:0]   io_in_r_bypass_regNext_13_2_data_15;
  reg                 io_in_r_bypass_regNext_13_2_load_store_15;
  reg                 io_in_r_bypass_regNext_13_2_df_is_ws_15;
  reg                 io_in_r_bypass_regNext_13_2_stall_15;
  reg        [15:0]   io_in_r_bypass_regNext_13_3_data_15;
  reg                 io_in_r_bypass_regNext_13_3_load_store_15;
  reg                 io_in_r_bypass_regNext_13_3_df_is_ws_15;
  reg                 io_in_r_bypass_regNext_13_3_stall_15;
  reg        [15:0]   io_in_r_bypass_regNext_14_0_data_15;
  reg                 io_in_r_bypass_regNext_14_0_load_store_15;
  reg                 io_in_r_bypass_regNext_14_0_df_is_ws_15;
  reg                 io_in_r_bypass_regNext_14_0_stall_15;
  reg        [15:0]   io_in_r_bypass_regNext_14_1_data_15;
  reg                 io_in_r_bypass_regNext_14_1_load_store_15;
  reg                 io_in_r_bypass_regNext_14_1_df_is_ws_15;
  reg                 io_in_r_bypass_regNext_14_1_stall_15;
  reg        [15:0]   io_in_r_bypass_regNext_14_2_data_15;
  reg                 io_in_r_bypass_regNext_14_2_load_store_15;
  reg                 io_in_r_bypass_regNext_14_2_df_is_ws_15;
  reg                 io_in_r_bypass_regNext_14_2_stall_15;
  reg        [15:0]   io_in_r_bypass_regNext_14_3_data_15;
  reg                 io_in_r_bypass_regNext_14_3_load_store_15;
  reg                 io_in_r_bypass_regNext_14_3_df_is_ws_15;
  reg                 io_in_r_bypass_regNext_14_3_stall_15;
  reg        [15:0]   io_in_r_bypass_regNext_15_0_data_15;
  reg                 io_in_r_bypass_regNext_15_0_load_store_15;
  reg                 io_in_r_bypass_regNext_15_0_df_is_ws_15;
  reg                 io_in_r_bypass_regNext_15_0_stall_15;
  reg        [15:0]   io_in_r_bypass_regNext_15_1_data_15;
  reg                 io_in_r_bypass_regNext_15_1_load_store_15;
  reg                 io_in_r_bypass_regNext_15_1_df_is_ws_15;
  reg                 io_in_r_bypass_regNext_15_1_stall_15;
  reg        [15:0]   io_in_r_bypass_regNext_15_2_data_15;
  reg                 io_in_r_bypass_regNext_15_2_load_store_15;
  reg                 io_in_r_bypass_regNext_15_2_df_is_ws_15;
  reg                 io_in_r_bypass_regNext_15_2_stall_15;
  reg        [15:0]   io_in_r_bypass_regNext_15_3_data_15;
  reg                 io_in_r_bypass_regNext_15_3_load_store_15;
  reg                 io_in_r_bypass_regNext_15_3_df_is_ws_15;
  reg                 io_in_r_bypass_regNext_15_3_stall_15;
  reg        [15:0]   io_in_r_bypass_regNext_16_0_data_15;
  reg                 io_in_r_bypass_regNext_16_0_load_store_15;
  reg                 io_in_r_bypass_regNext_16_0_df_is_ws_15;
  reg                 io_in_r_bypass_regNext_16_0_stall_15;
  reg        [15:0]   io_in_r_bypass_regNext_16_1_data_15;
  reg                 io_in_r_bypass_regNext_16_1_load_store_15;
  reg                 io_in_r_bypass_regNext_16_1_df_is_ws_15;
  reg                 io_in_r_bypass_regNext_16_1_stall_15;
  reg        [15:0]   io_in_r_bypass_regNext_16_2_data_15;
  reg                 io_in_r_bypass_regNext_16_2_load_store_15;
  reg                 io_in_r_bypass_regNext_16_2_df_is_ws_15;
  reg                 io_in_r_bypass_regNext_16_2_stall_15;
  reg        [15:0]   io_in_r_bypass_regNext_16_3_data_15;
  reg                 io_in_r_bypass_regNext_16_3_load_store_15;
  reg                 io_in_r_bypass_regNext_16_3_df_is_ws_15;
  reg                 io_in_r_bypass_regNext_16_3_stall_15;
  reg        [15:0]   io_in_r_bypass_regNext_17_0_data_15;
  reg                 io_in_r_bypass_regNext_17_0_load_store_15;
  reg                 io_in_r_bypass_regNext_17_0_df_is_ws_15;
  reg                 io_in_r_bypass_regNext_17_0_stall_15;
  reg        [15:0]   io_in_r_bypass_regNext_17_1_data_15;
  reg                 io_in_r_bypass_regNext_17_1_load_store_15;
  reg                 io_in_r_bypass_regNext_17_1_df_is_ws_15;
  reg                 io_in_r_bypass_regNext_17_1_stall_15;
  reg        [15:0]   io_in_r_bypass_regNext_17_2_data_15;
  reg                 io_in_r_bypass_regNext_17_2_load_store_15;
  reg                 io_in_r_bypass_regNext_17_2_df_is_ws_15;
  reg                 io_in_r_bypass_regNext_17_2_stall_15;
  reg        [15:0]   io_in_r_bypass_regNext_17_3_data_15;
  reg                 io_in_r_bypass_regNext_17_3_load_store_15;
  reg                 io_in_r_bypass_regNext_17_3_df_is_ws_15;
  reg                 io_in_r_bypass_regNext_17_3_stall_15;
  reg        [15:0]   io_in_r_bypass_regNext_18_0_data_15;
  reg                 io_in_r_bypass_regNext_18_0_load_store_15;
  reg                 io_in_r_bypass_regNext_18_0_df_is_ws_15;
  reg                 io_in_r_bypass_regNext_18_0_stall_15;
  reg        [15:0]   io_in_r_bypass_regNext_18_1_data_15;
  reg                 io_in_r_bypass_regNext_18_1_load_store_15;
  reg                 io_in_r_bypass_regNext_18_1_df_is_ws_15;
  reg                 io_in_r_bypass_regNext_18_1_stall_15;
  reg        [15:0]   io_in_r_bypass_regNext_18_2_data_15;
  reg                 io_in_r_bypass_regNext_18_2_load_store_15;
  reg                 io_in_r_bypass_regNext_18_2_df_is_ws_15;
  reg                 io_in_r_bypass_regNext_18_2_stall_15;
  reg        [15:0]   io_in_r_bypass_regNext_18_3_data_15;
  reg                 io_in_r_bypass_regNext_18_3_load_store_15;
  reg                 io_in_r_bypass_regNext_18_3_df_is_ws_15;
  reg                 io_in_r_bypass_regNext_18_3_stall_15;
  reg        [15:0]   io_in_r_bypass_regNext_19_0_data_15;
  reg                 io_in_r_bypass_regNext_19_0_load_store_15;
  reg                 io_in_r_bypass_regNext_19_0_df_is_ws_15;
  reg                 io_in_r_bypass_regNext_19_0_stall_15;
  reg        [15:0]   io_in_r_bypass_regNext_19_1_data_15;
  reg                 io_in_r_bypass_regNext_19_1_load_store_15;
  reg                 io_in_r_bypass_regNext_19_1_df_is_ws_15;
  reg                 io_in_r_bypass_regNext_19_1_stall_15;
  reg        [15:0]   io_in_r_bypass_regNext_19_2_data_15;
  reg                 io_in_r_bypass_regNext_19_2_load_store_15;
  reg                 io_in_r_bypass_regNext_19_2_df_is_ws_15;
  reg                 io_in_r_bypass_regNext_19_2_stall_15;
  reg        [15:0]   io_in_r_bypass_regNext_19_3_data_15;
  reg                 io_in_r_bypass_regNext_19_3_load_store_15;
  reg                 io_in_r_bypass_regNext_19_3_df_is_ws_15;
  reg                 io_in_r_bypass_regNext_19_3_stall_15;
  reg        [15:0]   io_in_r_bypass_regNext_20_0_data_15;
  reg                 io_in_r_bypass_regNext_20_0_load_store_15;
  reg                 io_in_r_bypass_regNext_20_0_df_is_ws_15;
  reg                 io_in_r_bypass_regNext_20_0_stall_15;
  reg        [15:0]   io_in_r_bypass_regNext_20_1_data_15;
  reg                 io_in_r_bypass_regNext_20_1_load_store_15;
  reg                 io_in_r_bypass_regNext_20_1_df_is_ws_15;
  reg                 io_in_r_bypass_regNext_20_1_stall_15;
  reg        [15:0]   io_in_r_bypass_regNext_20_2_data_15;
  reg                 io_in_r_bypass_regNext_20_2_load_store_15;
  reg                 io_in_r_bypass_regNext_20_2_df_is_ws_15;
  reg                 io_in_r_bypass_regNext_20_2_stall_15;
  reg        [15:0]   io_in_r_bypass_regNext_20_3_data_15;
  reg                 io_in_r_bypass_regNext_20_3_load_store_15;
  reg                 io_in_r_bypass_regNext_20_3_df_is_ws_15;
  reg                 io_in_r_bypass_regNext_20_3_stall_15;
  reg        [15:0]   io_in_r_bypass_regNext_21_0_data_15;
  reg                 io_in_r_bypass_regNext_21_0_load_store_15;
  reg                 io_in_r_bypass_regNext_21_0_df_is_ws_15;
  reg                 io_in_r_bypass_regNext_21_0_stall_15;
  reg        [15:0]   io_in_r_bypass_regNext_21_1_data_15;
  reg                 io_in_r_bypass_regNext_21_1_load_store_15;
  reg                 io_in_r_bypass_regNext_21_1_df_is_ws_15;
  reg                 io_in_r_bypass_regNext_21_1_stall_15;
  reg        [15:0]   io_in_r_bypass_regNext_21_2_data_15;
  reg                 io_in_r_bypass_regNext_21_2_load_store_15;
  reg                 io_in_r_bypass_regNext_21_2_df_is_ws_15;
  reg                 io_in_r_bypass_regNext_21_2_stall_15;
  reg        [15:0]   io_in_r_bypass_regNext_21_3_data_15;
  reg                 io_in_r_bypass_regNext_21_3_load_store_15;
  reg                 io_in_r_bypass_regNext_21_3_df_is_ws_15;
  reg                 io_in_r_bypass_regNext_21_3_stall_15;
  reg        [15:0]   io_in_r_bypass_regNext_22_0_data_15;
  reg                 io_in_r_bypass_regNext_22_0_load_store_15;
  reg                 io_in_r_bypass_regNext_22_0_df_is_ws_15;
  reg                 io_in_r_bypass_regNext_22_0_stall_15;
  reg        [15:0]   io_in_r_bypass_regNext_22_1_data_15;
  reg                 io_in_r_bypass_regNext_22_1_load_store_15;
  reg                 io_in_r_bypass_regNext_22_1_df_is_ws_15;
  reg                 io_in_r_bypass_regNext_22_1_stall_15;
  reg        [15:0]   io_in_r_bypass_regNext_22_2_data_15;
  reg                 io_in_r_bypass_regNext_22_2_load_store_15;
  reg                 io_in_r_bypass_regNext_22_2_df_is_ws_15;
  reg                 io_in_r_bypass_regNext_22_2_stall_15;
  reg        [15:0]   io_in_r_bypass_regNext_22_3_data_15;
  reg                 io_in_r_bypass_regNext_22_3_load_store_15;
  reg                 io_in_r_bypass_regNext_22_3_df_is_ws_15;
  reg                 io_in_r_bypass_regNext_22_3_stall_15;
  reg        [15:0]   io_in_r_bypass_regNext_23_0_data_15;
  reg                 io_in_r_bypass_regNext_23_0_load_store_15;
  reg                 io_in_r_bypass_regNext_23_0_df_is_ws_15;
  reg                 io_in_r_bypass_regNext_23_0_stall_15;
  reg        [15:0]   io_in_r_bypass_regNext_23_1_data_15;
  reg                 io_in_r_bypass_regNext_23_1_load_store_15;
  reg                 io_in_r_bypass_regNext_23_1_df_is_ws_15;
  reg                 io_in_r_bypass_regNext_23_1_stall_15;
  reg        [15:0]   io_in_r_bypass_regNext_23_2_data_15;
  reg                 io_in_r_bypass_regNext_23_2_load_store_15;
  reg                 io_in_r_bypass_regNext_23_2_df_is_ws_15;
  reg                 io_in_r_bypass_regNext_23_2_stall_15;
  reg        [15:0]   io_in_r_bypass_regNext_23_3_data_15;
  reg                 io_in_r_bypass_regNext_23_3_load_store_15;
  reg                 io_in_r_bypass_regNext_23_3_df_is_ws_15;
  reg                 io_in_r_bypass_regNext_23_3_stall_15;
  reg        [15:0]   io_in_r_bypass_regNext_24_0_data_15;
  reg                 io_in_r_bypass_regNext_24_0_load_store_15;
  reg                 io_in_r_bypass_regNext_24_0_df_is_ws_15;
  reg                 io_in_r_bypass_regNext_24_0_stall_15;
  reg        [15:0]   io_in_r_bypass_regNext_24_1_data_15;
  reg                 io_in_r_bypass_regNext_24_1_load_store_15;
  reg                 io_in_r_bypass_regNext_24_1_df_is_ws_15;
  reg                 io_in_r_bypass_regNext_24_1_stall_15;
  reg        [15:0]   io_in_r_bypass_regNext_24_2_data_15;
  reg                 io_in_r_bypass_regNext_24_2_load_store_15;
  reg                 io_in_r_bypass_regNext_24_2_df_is_ws_15;
  reg                 io_in_r_bypass_regNext_24_2_stall_15;
  reg        [15:0]   io_in_r_bypass_regNext_24_3_data_15;
  reg                 io_in_r_bypass_regNext_24_3_load_store_15;
  reg                 io_in_r_bypass_regNext_24_3_df_is_ws_15;
  reg                 io_in_r_bypass_regNext_24_3_stall_15;
  reg        [15:0]   io_in_r_bypass_regNext_25_0_data_15;
  reg                 io_in_r_bypass_regNext_25_0_load_store_15;
  reg                 io_in_r_bypass_regNext_25_0_df_is_ws_15;
  reg                 io_in_r_bypass_regNext_25_0_stall_15;
  reg        [15:0]   io_in_r_bypass_regNext_25_1_data_15;
  reg                 io_in_r_bypass_regNext_25_1_load_store_15;
  reg                 io_in_r_bypass_regNext_25_1_df_is_ws_15;
  reg                 io_in_r_bypass_regNext_25_1_stall_15;
  reg        [15:0]   io_in_r_bypass_regNext_25_2_data_15;
  reg                 io_in_r_bypass_regNext_25_2_load_store_15;
  reg                 io_in_r_bypass_regNext_25_2_df_is_ws_15;
  reg                 io_in_r_bypass_regNext_25_2_stall_15;
  reg        [15:0]   io_in_r_bypass_regNext_25_3_data_15;
  reg                 io_in_r_bypass_regNext_25_3_load_store_15;
  reg                 io_in_r_bypass_regNext_25_3_df_is_ws_15;
  reg                 io_in_r_bypass_regNext_25_3_stall_15;
  reg        [15:0]   io_in_r_bypass_regNext_26_0_data_15;
  reg                 io_in_r_bypass_regNext_26_0_load_store_15;
  reg                 io_in_r_bypass_regNext_26_0_df_is_ws_15;
  reg                 io_in_r_bypass_regNext_26_0_stall_15;
  reg        [15:0]   io_in_r_bypass_regNext_26_1_data_15;
  reg                 io_in_r_bypass_regNext_26_1_load_store_15;
  reg                 io_in_r_bypass_regNext_26_1_df_is_ws_15;
  reg                 io_in_r_bypass_regNext_26_1_stall_15;
  reg        [15:0]   io_in_r_bypass_regNext_26_2_data_15;
  reg                 io_in_r_bypass_regNext_26_2_load_store_15;
  reg                 io_in_r_bypass_regNext_26_2_df_is_ws_15;
  reg                 io_in_r_bypass_regNext_26_2_stall_15;
  reg        [15:0]   io_in_r_bypass_regNext_26_3_data_15;
  reg                 io_in_r_bypass_regNext_26_3_load_store_15;
  reg                 io_in_r_bypass_regNext_26_3_df_is_ws_15;
  reg                 io_in_r_bypass_regNext_26_3_stall_15;
  reg        [15:0]   io_in_r_bypass_regNext_27_0_data_15;
  reg                 io_in_r_bypass_regNext_27_0_load_store_15;
  reg                 io_in_r_bypass_regNext_27_0_df_is_ws_15;
  reg                 io_in_r_bypass_regNext_27_0_stall_15;
  reg        [15:0]   io_in_r_bypass_regNext_27_1_data_15;
  reg                 io_in_r_bypass_regNext_27_1_load_store_15;
  reg                 io_in_r_bypass_regNext_27_1_df_is_ws_15;
  reg                 io_in_r_bypass_regNext_27_1_stall_15;
  reg        [15:0]   io_in_r_bypass_regNext_27_2_data_15;
  reg                 io_in_r_bypass_regNext_27_2_load_store_15;
  reg                 io_in_r_bypass_regNext_27_2_df_is_ws_15;
  reg                 io_in_r_bypass_regNext_27_2_stall_15;
  reg        [15:0]   io_in_r_bypass_regNext_27_3_data_15;
  reg                 io_in_r_bypass_regNext_27_3_load_store_15;
  reg                 io_in_r_bypass_regNext_27_3_df_is_ws_15;
  reg                 io_in_r_bypass_regNext_27_3_stall_15;
  reg        [15:0]   io_in_r_bypass_regNext_28_0_data_15;
  reg                 io_in_r_bypass_regNext_28_0_load_store_15;
  reg                 io_in_r_bypass_regNext_28_0_df_is_ws_15;
  reg                 io_in_r_bypass_regNext_28_0_stall_15;
  reg        [15:0]   io_in_r_bypass_regNext_28_1_data_15;
  reg                 io_in_r_bypass_regNext_28_1_load_store_15;
  reg                 io_in_r_bypass_regNext_28_1_df_is_ws_15;
  reg                 io_in_r_bypass_regNext_28_1_stall_15;
  reg        [15:0]   io_in_r_bypass_regNext_28_2_data_15;
  reg                 io_in_r_bypass_regNext_28_2_load_store_15;
  reg                 io_in_r_bypass_regNext_28_2_df_is_ws_15;
  reg                 io_in_r_bypass_regNext_28_2_stall_15;
  reg        [15:0]   io_in_r_bypass_regNext_28_3_data_15;
  reg                 io_in_r_bypass_regNext_28_3_load_store_15;
  reg                 io_in_r_bypass_regNext_28_3_df_is_ws_15;
  reg                 io_in_r_bypass_regNext_28_3_stall_15;
  reg        [15:0]   io_in_r_bypass_regNext_29_0_data_15;
  reg                 io_in_r_bypass_regNext_29_0_load_store_15;
  reg                 io_in_r_bypass_regNext_29_0_df_is_ws_15;
  reg                 io_in_r_bypass_regNext_29_0_stall_15;
  reg        [15:0]   io_in_r_bypass_regNext_29_1_data_15;
  reg                 io_in_r_bypass_regNext_29_1_load_store_15;
  reg                 io_in_r_bypass_regNext_29_1_df_is_ws_15;
  reg                 io_in_r_bypass_regNext_29_1_stall_15;
  reg        [15:0]   io_in_r_bypass_regNext_29_2_data_15;
  reg                 io_in_r_bypass_regNext_29_2_load_store_15;
  reg                 io_in_r_bypass_regNext_29_2_df_is_ws_15;
  reg                 io_in_r_bypass_regNext_29_2_stall_15;
  reg        [15:0]   io_in_r_bypass_regNext_29_3_data_15;
  reg                 io_in_r_bypass_regNext_29_3_load_store_15;
  reg                 io_in_r_bypass_regNext_29_3_df_is_ws_15;
  reg                 io_in_r_bypass_regNext_29_3_stall_15;
  reg        [15:0]   io_in_r_bypass_regNext_30_0_data_15;
  reg                 io_in_r_bypass_regNext_30_0_load_store_15;
  reg                 io_in_r_bypass_regNext_30_0_df_is_ws_15;
  reg                 io_in_r_bypass_regNext_30_0_stall_15;
  reg        [15:0]   io_in_r_bypass_regNext_30_1_data_15;
  reg                 io_in_r_bypass_regNext_30_1_load_store_15;
  reg                 io_in_r_bypass_regNext_30_1_df_is_ws_15;
  reg                 io_in_r_bypass_regNext_30_1_stall_15;
  reg        [15:0]   io_in_r_bypass_regNext_30_2_data_15;
  reg                 io_in_r_bypass_regNext_30_2_load_store_15;
  reg                 io_in_r_bypass_regNext_30_2_df_is_ws_15;
  reg                 io_in_r_bypass_regNext_30_2_stall_15;
  reg        [15:0]   io_in_r_bypass_regNext_30_3_data_15;
  reg                 io_in_r_bypass_regNext_30_3_load_store_15;
  reg                 io_in_r_bypass_regNext_30_3_df_is_ws_15;
  reg                 io_in_r_bypass_regNext_30_3_stall_15;
  reg        [15:0]   io_in_r_bypass_regNext_31_0_data_15;
  reg                 io_in_r_bypass_regNext_31_0_load_store_15;
  reg                 io_in_r_bypass_regNext_31_0_df_is_ws_15;
  reg                 io_in_r_bypass_regNext_31_0_stall_15;
  reg        [15:0]   io_in_r_bypass_regNext_31_1_data_15;
  reg                 io_in_r_bypass_regNext_31_1_load_store_15;
  reg                 io_in_r_bypass_regNext_31_1_df_is_ws_15;
  reg                 io_in_r_bypass_regNext_31_1_stall_15;
  reg        [15:0]   io_in_r_bypass_regNext_31_2_data_15;
  reg                 io_in_r_bypass_regNext_31_2_load_store_15;
  reg                 io_in_r_bypass_regNext_31_2_df_is_ws_15;
  reg                 io_in_r_bypass_regNext_31_2_stall_15;
  reg        [15:0]   io_in_r_bypass_regNext_31_3_data_15;
  reg                 io_in_r_bypass_regNext_31_3_load_store_15;
  reg                 io_in_r_bypass_regNext_31_3_df_is_ws_15;
  reg                 io_in_r_bypass_regNext_31_3_stall_15;
  reg        [15:0]   io_in_r_bypass_regNext_0_0_data_16;
  reg                 io_in_r_bypass_regNext_0_0_load_store_16;
  reg                 io_in_r_bypass_regNext_0_0_df_is_ws_16;
  reg                 io_in_r_bypass_regNext_0_0_stall_16;
  reg        [15:0]   io_in_r_bypass_regNext_0_1_data_16;
  reg                 io_in_r_bypass_regNext_0_1_load_store_16;
  reg                 io_in_r_bypass_regNext_0_1_df_is_ws_16;
  reg                 io_in_r_bypass_regNext_0_1_stall_16;
  reg        [15:0]   io_in_r_bypass_regNext_0_2_data_16;
  reg                 io_in_r_bypass_regNext_0_2_load_store_16;
  reg                 io_in_r_bypass_regNext_0_2_df_is_ws_16;
  reg                 io_in_r_bypass_regNext_0_2_stall_16;
  reg        [15:0]   io_in_r_bypass_regNext_0_3_data_16;
  reg                 io_in_r_bypass_regNext_0_3_load_store_16;
  reg                 io_in_r_bypass_regNext_0_3_df_is_ws_16;
  reg                 io_in_r_bypass_regNext_0_3_stall_16;
  reg        [15:0]   io_in_r_bypass_regNext_1_0_data_16;
  reg                 io_in_r_bypass_regNext_1_0_load_store_16;
  reg                 io_in_r_bypass_regNext_1_0_df_is_ws_16;
  reg                 io_in_r_bypass_regNext_1_0_stall_16;
  reg        [15:0]   io_in_r_bypass_regNext_1_1_data_16;
  reg                 io_in_r_bypass_regNext_1_1_load_store_16;
  reg                 io_in_r_bypass_regNext_1_1_df_is_ws_16;
  reg                 io_in_r_bypass_regNext_1_1_stall_16;
  reg        [15:0]   io_in_r_bypass_regNext_1_2_data_16;
  reg                 io_in_r_bypass_regNext_1_2_load_store_16;
  reg                 io_in_r_bypass_regNext_1_2_df_is_ws_16;
  reg                 io_in_r_bypass_regNext_1_2_stall_16;
  reg        [15:0]   io_in_r_bypass_regNext_1_3_data_16;
  reg                 io_in_r_bypass_regNext_1_3_load_store_16;
  reg                 io_in_r_bypass_regNext_1_3_df_is_ws_16;
  reg                 io_in_r_bypass_regNext_1_3_stall_16;
  reg        [15:0]   io_in_r_bypass_regNext_2_0_data_16;
  reg                 io_in_r_bypass_regNext_2_0_load_store_16;
  reg                 io_in_r_bypass_regNext_2_0_df_is_ws_16;
  reg                 io_in_r_bypass_regNext_2_0_stall_16;
  reg        [15:0]   io_in_r_bypass_regNext_2_1_data_16;
  reg                 io_in_r_bypass_regNext_2_1_load_store_16;
  reg                 io_in_r_bypass_regNext_2_1_df_is_ws_16;
  reg                 io_in_r_bypass_regNext_2_1_stall_16;
  reg        [15:0]   io_in_r_bypass_regNext_2_2_data_16;
  reg                 io_in_r_bypass_regNext_2_2_load_store_16;
  reg                 io_in_r_bypass_regNext_2_2_df_is_ws_16;
  reg                 io_in_r_bypass_regNext_2_2_stall_16;
  reg        [15:0]   io_in_r_bypass_regNext_2_3_data_16;
  reg                 io_in_r_bypass_regNext_2_3_load_store_16;
  reg                 io_in_r_bypass_regNext_2_3_df_is_ws_16;
  reg                 io_in_r_bypass_regNext_2_3_stall_16;
  reg        [15:0]   io_in_r_bypass_regNext_3_0_data_16;
  reg                 io_in_r_bypass_regNext_3_0_load_store_16;
  reg                 io_in_r_bypass_regNext_3_0_df_is_ws_16;
  reg                 io_in_r_bypass_regNext_3_0_stall_16;
  reg        [15:0]   io_in_r_bypass_regNext_3_1_data_16;
  reg                 io_in_r_bypass_regNext_3_1_load_store_16;
  reg                 io_in_r_bypass_regNext_3_1_df_is_ws_16;
  reg                 io_in_r_bypass_regNext_3_1_stall_16;
  reg        [15:0]   io_in_r_bypass_regNext_3_2_data_16;
  reg                 io_in_r_bypass_regNext_3_2_load_store_16;
  reg                 io_in_r_bypass_regNext_3_2_df_is_ws_16;
  reg                 io_in_r_bypass_regNext_3_2_stall_16;
  reg        [15:0]   io_in_r_bypass_regNext_3_3_data_16;
  reg                 io_in_r_bypass_regNext_3_3_load_store_16;
  reg                 io_in_r_bypass_regNext_3_3_df_is_ws_16;
  reg                 io_in_r_bypass_regNext_3_3_stall_16;
  reg        [15:0]   io_in_r_bypass_regNext_4_0_data_16;
  reg                 io_in_r_bypass_regNext_4_0_load_store_16;
  reg                 io_in_r_bypass_regNext_4_0_df_is_ws_16;
  reg                 io_in_r_bypass_regNext_4_0_stall_16;
  reg        [15:0]   io_in_r_bypass_regNext_4_1_data_16;
  reg                 io_in_r_bypass_regNext_4_1_load_store_16;
  reg                 io_in_r_bypass_regNext_4_1_df_is_ws_16;
  reg                 io_in_r_bypass_regNext_4_1_stall_16;
  reg        [15:0]   io_in_r_bypass_regNext_4_2_data_16;
  reg                 io_in_r_bypass_regNext_4_2_load_store_16;
  reg                 io_in_r_bypass_regNext_4_2_df_is_ws_16;
  reg                 io_in_r_bypass_regNext_4_2_stall_16;
  reg        [15:0]   io_in_r_bypass_regNext_4_3_data_16;
  reg                 io_in_r_bypass_regNext_4_3_load_store_16;
  reg                 io_in_r_bypass_regNext_4_3_df_is_ws_16;
  reg                 io_in_r_bypass_regNext_4_3_stall_16;
  reg        [15:0]   io_in_r_bypass_regNext_5_0_data_16;
  reg                 io_in_r_bypass_regNext_5_0_load_store_16;
  reg                 io_in_r_bypass_regNext_5_0_df_is_ws_16;
  reg                 io_in_r_bypass_regNext_5_0_stall_16;
  reg        [15:0]   io_in_r_bypass_regNext_5_1_data_16;
  reg                 io_in_r_bypass_regNext_5_1_load_store_16;
  reg                 io_in_r_bypass_regNext_5_1_df_is_ws_16;
  reg                 io_in_r_bypass_regNext_5_1_stall_16;
  reg        [15:0]   io_in_r_bypass_regNext_5_2_data_16;
  reg                 io_in_r_bypass_regNext_5_2_load_store_16;
  reg                 io_in_r_bypass_regNext_5_2_df_is_ws_16;
  reg                 io_in_r_bypass_regNext_5_2_stall_16;
  reg        [15:0]   io_in_r_bypass_regNext_5_3_data_16;
  reg                 io_in_r_bypass_regNext_5_3_load_store_16;
  reg                 io_in_r_bypass_regNext_5_3_df_is_ws_16;
  reg                 io_in_r_bypass_regNext_5_3_stall_16;
  reg        [15:0]   io_in_r_bypass_regNext_6_0_data_16;
  reg                 io_in_r_bypass_regNext_6_0_load_store_16;
  reg                 io_in_r_bypass_regNext_6_0_df_is_ws_16;
  reg                 io_in_r_bypass_regNext_6_0_stall_16;
  reg        [15:0]   io_in_r_bypass_regNext_6_1_data_16;
  reg                 io_in_r_bypass_regNext_6_1_load_store_16;
  reg                 io_in_r_bypass_regNext_6_1_df_is_ws_16;
  reg                 io_in_r_bypass_regNext_6_1_stall_16;
  reg        [15:0]   io_in_r_bypass_regNext_6_2_data_16;
  reg                 io_in_r_bypass_regNext_6_2_load_store_16;
  reg                 io_in_r_bypass_regNext_6_2_df_is_ws_16;
  reg                 io_in_r_bypass_regNext_6_2_stall_16;
  reg        [15:0]   io_in_r_bypass_regNext_6_3_data_16;
  reg                 io_in_r_bypass_regNext_6_3_load_store_16;
  reg                 io_in_r_bypass_regNext_6_3_df_is_ws_16;
  reg                 io_in_r_bypass_regNext_6_3_stall_16;
  reg        [15:0]   io_in_r_bypass_regNext_7_0_data_16;
  reg                 io_in_r_bypass_regNext_7_0_load_store_16;
  reg                 io_in_r_bypass_regNext_7_0_df_is_ws_16;
  reg                 io_in_r_bypass_regNext_7_0_stall_16;
  reg        [15:0]   io_in_r_bypass_regNext_7_1_data_16;
  reg                 io_in_r_bypass_regNext_7_1_load_store_16;
  reg                 io_in_r_bypass_regNext_7_1_df_is_ws_16;
  reg                 io_in_r_bypass_regNext_7_1_stall_16;
  reg        [15:0]   io_in_r_bypass_regNext_7_2_data_16;
  reg                 io_in_r_bypass_regNext_7_2_load_store_16;
  reg                 io_in_r_bypass_regNext_7_2_df_is_ws_16;
  reg                 io_in_r_bypass_regNext_7_2_stall_16;
  reg        [15:0]   io_in_r_bypass_regNext_7_3_data_16;
  reg                 io_in_r_bypass_regNext_7_3_load_store_16;
  reg                 io_in_r_bypass_regNext_7_3_df_is_ws_16;
  reg                 io_in_r_bypass_regNext_7_3_stall_16;
  reg        [15:0]   io_in_r_bypass_regNext_8_0_data_16;
  reg                 io_in_r_bypass_regNext_8_0_load_store_16;
  reg                 io_in_r_bypass_regNext_8_0_df_is_ws_16;
  reg                 io_in_r_bypass_regNext_8_0_stall_16;
  reg        [15:0]   io_in_r_bypass_regNext_8_1_data_16;
  reg                 io_in_r_bypass_regNext_8_1_load_store_16;
  reg                 io_in_r_bypass_regNext_8_1_df_is_ws_16;
  reg                 io_in_r_bypass_regNext_8_1_stall_16;
  reg        [15:0]   io_in_r_bypass_regNext_8_2_data_16;
  reg                 io_in_r_bypass_regNext_8_2_load_store_16;
  reg                 io_in_r_bypass_regNext_8_2_df_is_ws_16;
  reg                 io_in_r_bypass_regNext_8_2_stall_16;
  reg        [15:0]   io_in_r_bypass_regNext_8_3_data_16;
  reg                 io_in_r_bypass_regNext_8_3_load_store_16;
  reg                 io_in_r_bypass_regNext_8_3_df_is_ws_16;
  reg                 io_in_r_bypass_regNext_8_3_stall_16;
  reg        [15:0]   io_in_r_bypass_regNext_9_0_data_16;
  reg                 io_in_r_bypass_regNext_9_0_load_store_16;
  reg                 io_in_r_bypass_regNext_9_0_df_is_ws_16;
  reg                 io_in_r_bypass_regNext_9_0_stall_16;
  reg        [15:0]   io_in_r_bypass_regNext_9_1_data_16;
  reg                 io_in_r_bypass_regNext_9_1_load_store_16;
  reg                 io_in_r_bypass_regNext_9_1_df_is_ws_16;
  reg                 io_in_r_bypass_regNext_9_1_stall_16;
  reg        [15:0]   io_in_r_bypass_regNext_9_2_data_16;
  reg                 io_in_r_bypass_regNext_9_2_load_store_16;
  reg                 io_in_r_bypass_regNext_9_2_df_is_ws_16;
  reg                 io_in_r_bypass_regNext_9_2_stall_16;
  reg        [15:0]   io_in_r_bypass_regNext_9_3_data_16;
  reg                 io_in_r_bypass_regNext_9_3_load_store_16;
  reg                 io_in_r_bypass_regNext_9_3_df_is_ws_16;
  reg                 io_in_r_bypass_regNext_9_3_stall_16;
  reg        [15:0]   io_in_r_bypass_regNext_10_0_data_16;
  reg                 io_in_r_bypass_regNext_10_0_load_store_16;
  reg                 io_in_r_bypass_regNext_10_0_df_is_ws_16;
  reg                 io_in_r_bypass_regNext_10_0_stall_16;
  reg        [15:0]   io_in_r_bypass_regNext_10_1_data_16;
  reg                 io_in_r_bypass_regNext_10_1_load_store_16;
  reg                 io_in_r_bypass_regNext_10_1_df_is_ws_16;
  reg                 io_in_r_bypass_regNext_10_1_stall_16;
  reg        [15:0]   io_in_r_bypass_regNext_10_2_data_16;
  reg                 io_in_r_bypass_regNext_10_2_load_store_16;
  reg                 io_in_r_bypass_regNext_10_2_df_is_ws_16;
  reg                 io_in_r_bypass_regNext_10_2_stall_16;
  reg        [15:0]   io_in_r_bypass_regNext_10_3_data_16;
  reg                 io_in_r_bypass_regNext_10_3_load_store_16;
  reg                 io_in_r_bypass_regNext_10_3_df_is_ws_16;
  reg                 io_in_r_bypass_regNext_10_3_stall_16;
  reg        [15:0]   io_in_r_bypass_regNext_11_0_data_16;
  reg                 io_in_r_bypass_regNext_11_0_load_store_16;
  reg                 io_in_r_bypass_regNext_11_0_df_is_ws_16;
  reg                 io_in_r_bypass_regNext_11_0_stall_16;
  reg        [15:0]   io_in_r_bypass_regNext_11_1_data_16;
  reg                 io_in_r_bypass_regNext_11_1_load_store_16;
  reg                 io_in_r_bypass_regNext_11_1_df_is_ws_16;
  reg                 io_in_r_bypass_regNext_11_1_stall_16;
  reg        [15:0]   io_in_r_bypass_regNext_11_2_data_16;
  reg                 io_in_r_bypass_regNext_11_2_load_store_16;
  reg                 io_in_r_bypass_regNext_11_2_df_is_ws_16;
  reg                 io_in_r_bypass_regNext_11_2_stall_16;
  reg        [15:0]   io_in_r_bypass_regNext_11_3_data_16;
  reg                 io_in_r_bypass_regNext_11_3_load_store_16;
  reg                 io_in_r_bypass_regNext_11_3_df_is_ws_16;
  reg                 io_in_r_bypass_regNext_11_3_stall_16;
  reg        [15:0]   io_in_r_bypass_regNext_12_0_data_16;
  reg                 io_in_r_bypass_regNext_12_0_load_store_16;
  reg                 io_in_r_bypass_regNext_12_0_df_is_ws_16;
  reg                 io_in_r_bypass_regNext_12_0_stall_16;
  reg        [15:0]   io_in_r_bypass_regNext_12_1_data_16;
  reg                 io_in_r_bypass_regNext_12_1_load_store_16;
  reg                 io_in_r_bypass_regNext_12_1_df_is_ws_16;
  reg                 io_in_r_bypass_regNext_12_1_stall_16;
  reg        [15:0]   io_in_r_bypass_regNext_12_2_data_16;
  reg                 io_in_r_bypass_regNext_12_2_load_store_16;
  reg                 io_in_r_bypass_regNext_12_2_df_is_ws_16;
  reg                 io_in_r_bypass_regNext_12_2_stall_16;
  reg        [15:0]   io_in_r_bypass_regNext_12_3_data_16;
  reg                 io_in_r_bypass_regNext_12_3_load_store_16;
  reg                 io_in_r_bypass_regNext_12_3_df_is_ws_16;
  reg                 io_in_r_bypass_regNext_12_3_stall_16;
  reg        [15:0]   io_in_r_bypass_regNext_13_0_data_16;
  reg                 io_in_r_bypass_regNext_13_0_load_store_16;
  reg                 io_in_r_bypass_regNext_13_0_df_is_ws_16;
  reg                 io_in_r_bypass_regNext_13_0_stall_16;
  reg        [15:0]   io_in_r_bypass_regNext_13_1_data_16;
  reg                 io_in_r_bypass_regNext_13_1_load_store_16;
  reg                 io_in_r_bypass_regNext_13_1_df_is_ws_16;
  reg                 io_in_r_bypass_regNext_13_1_stall_16;
  reg        [15:0]   io_in_r_bypass_regNext_13_2_data_16;
  reg                 io_in_r_bypass_regNext_13_2_load_store_16;
  reg                 io_in_r_bypass_regNext_13_2_df_is_ws_16;
  reg                 io_in_r_bypass_regNext_13_2_stall_16;
  reg        [15:0]   io_in_r_bypass_regNext_13_3_data_16;
  reg                 io_in_r_bypass_regNext_13_3_load_store_16;
  reg                 io_in_r_bypass_regNext_13_3_df_is_ws_16;
  reg                 io_in_r_bypass_regNext_13_3_stall_16;
  reg        [15:0]   io_in_r_bypass_regNext_14_0_data_16;
  reg                 io_in_r_bypass_regNext_14_0_load_store_16;
  reg                 io_in_r_bypass_regNext_14_0_df_is_ws_16;
  reg                 io_in_r_bypass_regNext_14_0_stall_16;
  reg        [15:0]   io_in_r_bypass_regNext_14_1_data_16;
  reg                 io_in_r_bypass_regNext_14_1_load_store_16;
  reg                 io_in_r_bypass_regNext_14_1_df_is_ws_16;
  reg                 io_in_r_bypass_regNext_14_1_stall_16;
  reg        [15:0]   io_in_r_bypass_regNext_14_2_data_16;
  reg                 io_in_r_bypass_regNext_14_2_load_store_16;
  reg                 io_in_r_bypass_regNext_14_2_df_is_ws_16;
  reg                 io_in_r_bypass_regNext_14_2_stall_16;
  reg        [15:0]   io_in_r_bypass_regNext_14_3_data_16;
  reg                 io_in_r_bypass_regNext_14_3_load_store_16;
  reg                 io_in_r_bypass_regNext_14_3_df_is_ws_16;
  reg                 io_in_r_bypass_regNext_14_3_stall_16;
  reg        [15:0]   io_in_r_bypass_regNext_15_0_data_16;
  reg                 io_in_r_bypass_regNext_15_0_load_store_16;
  reg                 io_in_r_bypass_regNext_15_0_df_is_ws_16;
  reg                 io_in_r_bypass_regNext_15_0_stall_16;
  reg        [15:0]   io_in_r_bypass_regNext_15_1_data_16;
  reg                 io_in_r_bypass_regNext_15_1_load_store_16;
  reg                 io_in_r_bypass_regNext_15_1_df_is_ws_16;
  reg                 io_in_r_bypass_regNext_15_1_stall_16;
  reg        [15:0]   io_in_r_bypass_regNext_15_2_data_16;
  reg                 io_in_r_bypass_regNext_15_2_load_store_16;
  reg                 io_in_r_bypass_regNext_15_2_df_is_ws_16;
  reg                 io_in_r_bypass_regNext_15_2_stall_16;
  reg        [15:0]   io_in_r_bypass_regNext_15_3_data_16;
  reg                 io_in_r_bypass_regNext_15_3_load_store_16;
  reg                 io_in_r_bypass_regNext_15_3_df_is_ws_16;
  reg                 io_in_r_bypass_regNext_15_3_stall_16;
  reg        [15:0]   io_in_r_bypass_regNext_16_0_data_16;
  reg                 io_in_r_bypass_regNext_16_0_load_store_16;
  reg                 io_in_r_bypass_regNext_16_0_df_is_ws_16;
  reg                 io_in_r_bypass_regNext_16_0_stall_16;
  reg        [15:0]   io_in_r_bypass_regNext_16_1_data_16;
  reg                 io_in_r_bypass_regNext_16_1_load_store_16;
  reg                 io_in_r_bypass_regNext_16_1_df_is_ws_16;
  reg                 io_in_r_bypass_regNext_16_1_stall_16;
  reg        [15:0]   io_in_r_bypass_regNext_16_2_data_16;
  reg                 io_in_r_bypass_regNext_16_2_load_store_16;
  reg                 io_in_r_bypass_regNext_16_2_df_is_ws_16;
  reg                 io_in_r_bypass_regNext_16_2_stall_16;
  reg        [15:0]   io_in_r_bypass_regNext_16_3_data_16;
  reg                 io_in_r_bypass_regNext_16_3_load_store_16;
  reg                 io_in_r_bypass_regNext_16_3_df_is_ws_16;
  reg                 io_in_r_bypass_regNext_16_3_stall_16;
  reg        [15:0]   io_in_r_bypass_regNext_17_0_data_16;
  reg                 io_in_r_bypass_regNext_17_0_load_store_16;
  reg                 io_in_r_bypass_regNext_17_0_df_is_ws_16;
  reg                 io_in_r_bypass_regNext_17_0_stall_16;
  reg        [15:0]   io_in_r_bypass_regNext_17_1_data_16;
  reg                 io_in_r_bypass_regNext_17_1_load_store_16;
  reg                 io_in_r_bypass_regNext_17_1_df_is_ws_16;
  reg                 io_in_r_bypass_regNext_17_1_stall_16;
  reg        [15:0]   io_in_r_bypass_regNext_17_2_data_16;
  reg                 io_in_r_bypass_regNext_17_2_load_store_16;
  reg                 io_in_r_bypass_regNext_17_2_df_is_ws_16;
  reg                 io_in_r_bypass_regNext_17_2_stall_16;
  reg        [15:0]   io_in_r_bypass_regNext_17_3_data_16;
  reg                 io_in_r_bypass_regNext_17_3_load_store_16;
  reg                 io_in_r_bypass_regNext_17_3_df_is_ws_16;
  reg                 io_in_r_bypass_regNext_17_3_stall_16;
  reg        [15:0]   io_in_r_bypass_regNext_18_0_data_16;
  reg                 io_in_r_bypass_regNext_18_0_load_store_16;
  reg                 io_in_r_bypass_regNext_18_0_df_is_ws_16;
  reg                 io_in_r_bypass_regNext_18_0_stall_16;
  reg        [15:0]   io_in_r_bypass_regNext_18_1_data_16;
  reg                 io_in_r_bypass_regNext_18_1_load_store_16;
  reg                 io_in_r_bypass_regNext_18_1_df_is_ws_16;
  reg                 io_in_r_bypass_regNext_18_1_stall_16;
  reg        [15:0]   io_in_r_bypass_regNext_18_2_data_16;
  reg                 io_in_r_bypass_regNext_18_2_load_store_16;
  reg                 io_in_r_bypass_regNext_18_2_df_is_ws_16;
  reg                 io_in_r_bypass_regNext_18_2_stall_16;
  reg        [15:0]   io_in_r_bypass_regNext_18_3_data_16;
  reg                 io_in_r_bypass_regNext_18_3_load_store_16;
  reg                 io_in_r_bypass_regNext_18_3_df_is_ws_16;
  reg                 io_in_r_bypass_regNext_18_3_stall_16;
  reg        [15:0]   io_in_r_bypass_regNext_19_0_data_16;
  reg                 io_in_r_bypass_regNext_19_0_load_store_16;
  reg                 io_in_r_bypass_regNext_19_0_df_is_ws_16;
  reg                 io_in_r_bypass_regNext_19_0_stall_16;
  reg        [15:0]   io_in_r_bypass_regNext_19_1_data_16;
  reg                 io_in_r_bypass_regNext_19_1_load_store_16;
  reg                 io_in_r_bypass_regNext_19_1_df_is_ws_16;
  reg                 io_in_r_bypass_regNext_19_1_stall_16;
  reg        [15:0]   io_in_r_bypass_regNext_19_2_data_16;
  reg                 io_in_r_bypass_regNext_19_2_load_store_16;
  reg                 io_in_r_bypass_regNext_19_2_df_is_ws_16;
  reg                 io_in_r_bypass_regNext_19_2_stall_16;
  reg        [15:0]   io_in_r_bypass_regNext_19_3_data_16;
  reg                 io_in_r_bypass_regNext_19_3_load_store_16;
  reg                 io_in_r_bypass_regNext_19_3_df_is_ws_16;
  reg                 io_in_r_bypass_regNext_19_3_stall_16;
  reg        [15:0]   io_in_r_bypass_regNext_20_0_data_16;
  reg                 io_in_r_bypass_regNext_20_0_load_store_16;
  reg                 io_in_r_bypass_regNext_20_0_df_is_ws_16;
  reg                 io_in_r_bypass_regNext_20_0_stall_16;
  reg        [15:0]   io_in_r_bypass_regNext_20_1_data_16;
  reg                 io_in_r_bypass_regNext_20_1_load_store_16;
  reg                 io_in_r_bypass_regNext_20_1_df_is_ws_16;
  reg                 io_in_r_bypass_regNext_20_1_stall_16;
  reg        [15:0]   io_in_r_bypass_regNext_20_2_data_16;
  reg                 io_in_r_bypass_regNext_20_2_load_store_16;
  reg                 io_in_r_bypass_regNext_20_2_df_is_ws_16;
  reg                 io_in_r_bypass_regNext_20_2_stall_16;
  reg        [15:0]   io_in_r_bypass_regNext_20_3_data_16;
  reg                 io_in_r_bypass_regNext_20_3_load_store_16;
  reg                 io_in_r_bypass_regNext_20_3_df_is_ws_16;
  reg                 io_in_r_bypass_regNext_20_3_stall_16;
  reg        [15:0]   io_in_r_bypass_regNext_21_0_data_16;
  reg                 io_in_r_bypass_regNext_21_0_load_store_16;
  reg                 io_in_r_bypass_regNext_21_0_df_is_ws_16;
  reg                 io_in_r_bypass_regNext_21_0_stall_16;
  reg        [15:0]   io_in_r_bypass_regNext_21_1_data_16;
  reg                 io_in_r_bypass_regNext_21_1_load_store_16;
  reg                 io_in_r_bypass_regNext_21_1_df_is_ws_16;
  reg                 io_in_r_bypass_regNext_21_1_stall_16;
  reg        [15:0]   io_in_r_bypass_regNext_21_2_data_16;
  reg                 io_in_r_bypass_regNext_21_2_load_store_16;
  reg                 io_in_r_bypass_regNext_21_2_df_is_ws_16;
  reg                 io_in_r_bypass_regNext_21_2_stall_16;
  reg        [15:0]   io_in_r_bypass_regNext_21_3_data_16;
  reg                 io_in_r_bypass_regNext_21_3_load_store_16;
  reg                 io_in_r_bypass_regNext_21_3_df_is_ws_16;
  reg                 io_in_r_bypass_regNext_21_3_stall_16;
  reg        [15:0]   io_in_r_bypass_regNext_22_0_data_16;
  reg                 io_in_r_bypass_regNext_22_0_load_store_16;
  reg                 io_in_r_bypass_regNext_22_0_df_is_ws_16;
  reg                 io_in_r_bypass_regNext_22_0_stall_16;
  reg        [15:0]   io_in_r_bypass_regNext_22_1_data_16;
  reg                 io_in_r_bypass_regNext_22_1_load_store_16;
  reg                 io_in_r_bypass_regNext_22_1_df_is_ws_16;
  reg                 io_in_r_bypass_regNext_22_1_stall_16;
  reg        [15:0]   io_in_r_bypass_regNext_22_2_data_16;
  reg                 io_in_r_bypass_regNext_22_2_load_store_16;
  reg                 io_in_r_bypass_regNext_22_2_df_is_ws_16;
  reg                 io_in_r_bypass_regNext_22_2_stall_16;
  reg        [15:0]   io_in_r_bypass_regNext_22_3_data_16;
  reg                 io_in_r_bypass_regNext_22_3_load_store_16;
  reg                 io_in_r_bypass_regNext_22_3_df_is_ws_16;
  reg                 io_in_r_bypass_regNext_22_3_stall_16;
  reg        [15:0]   io_in_r_bypass_regNext_23_0_data_16;
  reg                 io_in_r_bypass_regNext_23_0_load_store_16;
  reg                 io_in_r_bypass_regNext_23_0_df_is_ws_16;
  reg                 io_in_r_bypass_regNext_23_0_stall_16;
  reg        [15:0]   io_in_r_bypass_regNext_23_1_data_16;
  reg                 io_in_r_bypass_regNext_23_1_load_store_16;
  reg                 io_in_r_bypass_regNext_23_1_df_is_ws_16;
  reg                 io_in_r_bypass_regNext_23_1_stall_16;
  reg        [15:0]   io_in_r_bypass_regNext_23_2_data_16;
  reg                 io_in_r_bypass_regNext_23_2_load_store_16;
  reg                 io_in_r_bypass_regNext_23_2_df_is_ws_16;
  reg                 io_in_r_bypass_regNext_23_2_stall_16;
  reg        [15:0]   io_in_r_bypass_regNext_23_3_data_16;
  reg                 io_in_r_bypass_regNext_23_3_load_store_16;
  reg                 io_in_r_bypass_regNext_23_3_df_is_ws_16;
  reg                 io_in_r_bypass_regNext_23_3_stall_16;
  reg        [15:0]   io_in_r_bypass_regNext_24_0_data_16;
  reg                 io_in_r_bypass_regNext_24_0_load_store_16;
  reg                 io_in_r_bypass_regNext_24_0_df_is_ws_16;
  reg                 io_in_r_bypass_regNext_24_0_stall_16;
  reg        [15:0]   io_in_r_bypass_regNext_24_1_data_16;
  reg                 io_in_r_bypass_regNext_24_1_load_store_16;
  reg                 io_in_r_bypass_regNext_24_1_df_is_ws_16;
  reg                 io_in_r_bypass_regNext_24_1_stall_16;
  reg        [15:0]   io_in_r_bypass_regNext_24_2_data_16;
  reg                 io_in_r_bypass_regNext_24_2_load_store_16;
  reg                 io_in_r_bypass_regNext_24_2_df_is_ws_16;
  reg                 io_in_r_bypass_regNext_24_2_stall_16;
  reg        [15:0]   io_in_r_bypass_regNext_24_3_data_16;
  reg                 io_in_r_bypass_regNext_24_3_load_store_16;
  reg                 io_in_r_bypass_regNext_24_3_df_is_ws_16;
  reg                 io_in_r_bypass_regNext_24_3_stall_16;
  reg        [15:0]   io_in_r_bypass_regNext_25_0_data_16;
  reg                 io_in_r_bypass_regNext_25_0_load_store_16;
  reg                 io_in_r_bypass_regNext_25_0_df_is_ws_16;
  reg                 io_in_r_bypass_regNext_25_0_stall_16;
  reg        [15:0]   io_in_r_bypass_regNext_25_1_data_16;
  reg                 io_in_r_bypass_regNext_25_1_load_store_16;
  reg                 io_in_r_bypass_regNext_25_1_df_is_ws_16;
  reg                 io_in_r_bypass_regNext_25_1_stall_16;
  reg        [15:0]   io_in_r_bypass_regNext_25_2_data_16;
  reg                 io_in_r_bypass_regNext_25_2_load_store_16;
  reg                 io_in_r_bypass_regNext_25_2_df_is_ws_16;
  reg                 io_in_r_bypass_regNext_25_2_stall_16;
  reg        [15:0]   io_in_r_bypass_regNext_25_3_data_16;
  reg                 io_in_r_bypass_regNext_25_3_load_store_16;
  reg                 io_in_r_bypass_regNext_25_3_df_is_ws_16;
  reg                 io_in_r_bypass_regNext_25_3_stall_16;
  reg        [15:0]   io_in_r_bypass_regNext_26_0_data_16;
  reg                 io_in_r_bypass_regNext_26_0_load_store_16;
  reg                 io_in_r_bypass_regNext_26_0_df_is_ws_16;
  reg                 io_in_r_bypass_regNext_26_0_stall_16;
  reg        [15:0]   io_in_r_bypass_regNext_26_1_data_16;
  reg                 io_in_r_bypass_regNext_26_1_load_store_16;
  reg                 io_in_r_bypass_regNext_26_1_df_is_ws_16;
  reg                 io_in_r_bypass_regNext_26_1_stall_16;
  reg        [15:0]   io_in_r_bypass_regNext_26_2_data_16;
  reg                 io_in_r_bypass_regNext_26_2_load_store_16;
  reg                 io_in_r_bypass_regNext_26_2_df_is_ws_16;
  reg                 io_in_r_bypass_regNext_26_2_stall_16;
  reg        [15:0]   io_in_r_bypass_regNext_26_3_data_16;
  reg                 io_in_r_bypass_regNext_26_3_load_store_16;
  reg                 io_in_r_bypass_regNext_26_3_df_is_ws_16;
  reg                 io_in_r_bypass_regNext_26_3_stall_16;
  reg        [15:0]   io_in_r_bypass_regNext_27_0_data_16;
  reg                 io_in_r_bypass_regNext_27_0_load_store_16;
  reg                 io_in_r_bypass_regNext_27_0_df_is_ws_16;
  reg                 io_in_r_bypass_regNext_27_0_stall_16;
  reg        [15:0]   io_in_r_bypass_regNext_27_1_data_16;
  reg                 io_in_r_bypass_regNext_27_1_load_store_16;
  reg                 io_in_r_bypass_regNext_27_1_df_is_ws_16;
  reg                 io_in_r_bypass_regNext_27_1_stall_16;
  reg        [15:0]   io_in_r_bypass_regNext_27_2_data_16;
  reg                 io_in_r_bypass_regNext_27_2_load_store_16;
  reg                 io_in_r_bypass_regNext_27_2_df_is_ws_16;
  reg                 io_in_r_bypass_regNext_27_2_stall_16;
  reg        [15:0]   io_in_r_bypass_regNext_27_3_data_16;
  reg                 io_in_r_bypass_regNext_27_3_load_store_16;
  reg                 io_in_r_bypass_regNext_27_3_df_is_ws_16;
  reg                 io_in_r_bypass_regNext_27_3_stall_16;
  reg        [15:0]   io_in_r_bypass_regNext_28_0_data_16;
  reg                 io_in_r_bypass_regNext_28_0_load_store_16;
  reg                 io_in_r_bypass_regNext_28_0_df_is_ws_16;
  reg                 io_in_r_bypass_regNext_28_0_stall_16;
  reg        [15:0]   io_in_r_bypass_regNext_28_1_data_16;
  reg                 io_in_r_bypass_regNext_28_1_load_store_16;
  reg                 io_in_r_bypass_regNext_28_1_df_is_ws_16;
  reg                 io_in_r_bypass_regNext_28_1_stall_16;
  reg        [15:0]   io_in_r_bypass_regNext_28_2_data_16;
  reg                 io_in_r_bypass_regNext_28_2_load_store_16;
  reg                 io_in_r_bypass_regNext_28_2_df_is_ws_16;
  reg                 io_in_r_bypass_regNext_28_2_stall_16;
  reg        [15:0]   io_in_r_bypass_regNext_28_3_data_16;
  reg                 io_in_r_bypass_regNext_28_3_load_store_16;
  reg                 io_in_r_bypass_regNext_28_3_df_is_ws_16;
  reg                 io_in_r_bypass_regNext_28_3_stall_16;
  reg        [15:0]   io_in_r_bypass_regNext_29_0_data_16;
  reg                 io_in_r_bypass_regNext_29_0_load_store_16;
  reg                 io_in_r_bypass_regNext_29_0_df_is_ws_16;
  reg                 io_in_r_bypass_regNext_29_0_stall_16;
  reg        [15:0]   io_in_r_bypass_regNext_29_1_data_16;
  reg                 io_in_r_bypass_regNext_29_1_load_store_16;
  reg                 io_in_r_bypass_regNext_29_1_df_is_ws_16;
  reg                 io_in_r_bypass_regNext_29_1_stall_16;
  reg        [15:0]   io_in_r_bypass_regNext_29_2_data_16;
  reg                 io_in_r_bypass_regNext_29_2_load_store_16;
  reg                 io_in_r_bypass_regNext_29_2_df_is_ws_16;
  reg                 io_in_r_bypass_regNext_29_2_stall_16;
  reg        [15:0]   io_in_r_bypass_regNext_29_3_data_16;
  reg                 io_in_r_bypass_regNext_29_3_load_store_16;
  reg                 io_in_r_bypass_regNext_29_3_df_is_ws_16;
  reg                 io_in_r_bypass_regNext_29_3_stall_16;
  reg        [15:0]   io_in_r_bypass_regNext_30_0_data_16;
  reg                 io_in_r_bypass_regNext_30_0_load_store_16;
  reg                 io_in_r_bypass_regNext_30_0_df_is_ws_16;
  reg                 io_in_r_bypass_regNext_30_0_stall_16;
  reg        [15:0]   io_in_r_bypass_regNext_30_1_data_16;
  reg                 io_in_r_bypass_regNext_30_1_load_store_16;
  reg                 io_in_r_bypass_regNext_30_1_df_is_ws_16;
  reg                 io_in_r_bypass_regNext_30_1_stall_16;
  reg        [15:0]   io_in_r_bypass_regNext_30_2_data_16;
  reg                 io_in_r_bypass_regNext_30_2_load_store_16;
  reg                 io_in_r_bypass_regNext_30_2_df_is_ws_16;
  reg                 io_in_r_bypass_regNext_30_2_stall_16;
  reg        [15:0]   io_in_r_bypass_regNext_30_3_data_16;
  reg                 io_in_r_bypass_regNext_30_3_load_store_16;
  reg                 io_in_r_bypass_regNext_30_3_df_is_ws_16;
  reg                 io_in_r_bypass_regNext_30_3_stall_16;
  reg        [15:0]   io_in_r_bypass_regNext_31_0_data_16;
  reg                 io_in_r_bypass_regNext_31_0_load_store_16;
  reg                 io_in_r_bypass_regNext_31_0_df_is_ws_16;
  reg                 io_in_r_bypass_regNext_31_0_stall_16;
  reg        [15:0]   io_in_r_bypass_regNext_31_1_data_16;
  reg                 io_in_r_bypass_regNext_31_1_load_store_16;
  reg                 io_in_r_bypass_regNext_31_1_df_is_ws_16;
  reg                 io_in_r_bypass_regNext_31_1_stall_16;
  reg        [15:0]   io_in_r_bypass_regNext_31_2_data_16;
  reg                 io_in_r_bypass_regNext_31_2_load_store_16;
  reg                 io_in_r_bypass_regNext_31_2_df_is_ws_16;
  reg                 io_in_r_bypass_regNext_31_2_stall_16;
  reg        [15:0]   io_in_r_bypass_regNext_31_3_data_16;
  reg                 io_in_r_bypass_regNext_31_3_load_store_16;
  reg                 io_in_r_bypass_regNext_31_3_df_is_ws_16;
  reg                 io_in_r_bypass_regNext_31_3_stall_16;
  reg        [15:0]   io_in_r_bypass_regNext_0_0_data_17;
  reg                 io_in_r_bypass_regNext_0_0_load_store_17;
  reg                 io_in_r_bypass_regNext_0_0_df_is_ws_17;
  reg                 io_in_r_bypass_regNext_0_0_stall_17;
  reg        [15:0]   io_in_r_bypass_regNext_0_1_data_17;
  reg                 io_in_r_bypass_regNext_0_1_load_store_17;
  reg                 io_in_r_bypass_regNext_0_1_df_is_ws_17;
  reg                 io_in_r_bypass_regNext_0_1_stall_17;
  reg        [15:0]   io_in_r_bypass_regNext_0_2_data_17;
  reg                 io_in_r_bypass_regNext_0_2_load_store_17;
  reg                 io_in_r_bypass_regNext_0_2_df_is_ws_17;
  reg                 io_in_r_bypass_regNext_0_2_stall_17;
  reg        [15:0]   io_in_r_bypass_regNext_0_3_data_17;
  reg                 io_in_r_bypass_regNext_0_3_load_store_17;
  reg                 io_in_r_bypass_regNext_0_3_df_is_ws_17;
  reg                 io_in_r_bypass_regNext_0_3_stall_17;
  reg        [15:0]   io_in_r_bypass_regNext_1_0_data_17;
  reg                 io_in_r_bypass_regNext_1_0_load_store_17;
  reg                 io_in_r_bypass_regNext_1_0_df_is_ws_17;
  reg                 io_in_r_bypass_regNext_1_0_stall_17;
  reg        [15:0]   io_in_r_bypass_regNext_1_1_data_17;
  reg                 io_in_r_bypass_regNext_1_1_load_store_17;
  reg                 io_in_r_bypass_regNext_1_1_df_is_ws_17;
  reg                 io_in_r_bypass_regNext_1_1_stall_17;
  reg        [15:0]   io_in_r_bypass_regNext_1_2_data_17;
  reg                 io_in_r_bypass_regNext_1_2_load_store_17;
  reg                 io_in_r_bypass_regNext_1_2_df_is_ws_17;
  reg                 io_in_r_bypass_regNext_1_2_stall_17;
  reg        [15:0]   io_in_r_bypass_regNext_1_3_data_17;
  reg                 io_in_r_bypass_regNext_1_3_load_store_17;
  reg                 io_in_r_bypass_regNext_1_3_df_is_ws_17;
  reg                 io_in_r_bypass_regNext_1_3_stall_17;
  reg        [15:0]   io_in_r_bypass_regNext_2_0_data_17;
  reg                 io_in_r_bypass_regNext_2_0_load_store_17;
  reg                 io_in_r_bypass_regNext_2_0_df_is_ws_17;
  reg                 io_in_r_bypass_regNext_2_0_stall_17;
  reg        [15:0]   io_in_r_bypass_regNext_2_1_data_17;
  reg                 io_in_r_bypass_regNext_2_1_load_store_17;
  reg                 io_in_r_bypass_regNext_2_1_df_is_ws_17;
  reg                 io_in_r_bypass_regNext_2_1_stall_17;
  reg        [15:0]   io_in_r_bypass_regNext_2_2_data_17;
  reg                 io_in_r_bypass_regNext_2_2_load_store_17;
  reg                 io_in_r_bypass_regNext_2_2_df_is_ws_17;
  reg                 io_in_r_bypass_regNext_2_2_stall_17;
  reg        [15:0]   io_in_r_bypass_regNext_2_3_data_17;
  reg                 io_in_r_bypass_regNext_2_3_load_store_17;
  reg                 io_in_r_bypass_regNext_2_3_df_is_ws_17;
  reg                 io_in_r_bypass_regNext_2_3_stall_17;
  reg        [15:0]   io_in_r_bypass_regNext_3_0_data_17;
  reg                 io_in_r_bypass_regNext_3_0_load_store_17;
  reg                 io_in_r_bypass_regNext_3_0_df_is_ws_17;
  reg                 io_in_r_bypass_regNext_3_0_stall_17;
  reg        [15:0]   io_in_r_bypass_regNext_3_1_data_17;
  reg                 io_in_r_bypass_regNext_3_1_load_store_17;
  reg                 io_in_r_bypass_regNext_3_1_df_is_ws_17;
  reg                 io_in_r_bypass_regNext_3_1_stall_17;
  reg        [15:0]   io_in_r_bypass_regNext_3_2_data_17;
  reg                 io_in_r_bypass_regNext_3_2_load_store_17;
  reg                 io_in_r_bypass_regNext_3_2_df_is_ws_17;
  reg                 io_in_r_bypass_regNext_3_2_stall_17;
  reg        [15:0]   io_in_r_bypass_regNext_3_3_data_17;
  reg                 io_in_r_bypass_regNext_3_3_load_store_17;
  reg                 io_in_r_bypass_regNext_3_3_df_is_ws_17;
  reg                 io_in_r_bypass_regNext_3_3_stall_17;
  reg        [15:0]   io_in_r_bypass_regNext_4_0_data_17;
  reg                 io_in_r_bypass_regNext_4_0_load_store_17;
  reg                 io_in_r_bypass_regNext_4_0_df_is_ws_17;
  reg                 io_in_r_bypass_regNext_4_0_stall_17;
  reg        [15:0]   io_in_r_bypass_regNext_4_1_data_17;
  reg                 io_in_r_bypass_regNext_4_1_load_store_17;
  reg                 io_in_r_bypass_regNext_4_1_df_is_ws_17;
  reg                 io_in_r_bypass_regNext_4_1_stall_17;
  reg        [15:0]   io_in_r_bypass_regNext_4_2_data_17;
  reg                 io_in_r_bypass_regNext_4_2_load_store_17;
  reg                 io_in_r_bypass_regNext_4_2_df_is_ws_17;
  reg                 io_in_r_bypass_regNext_4_2_stall_17;
  reg        [15:0]   io_in_r_bypass_regNext_4_3_data_17;
  reg                 io_in_r_bypass_regNext_4_3_load_store_17;
  reg                 io_in_r_bypass_regNext_4_3_df_is_ws_17;
  reg                 io_in_r_bypass_regNext_4_3_stall_17;
  reg        [15:0]   io_in_r_bypass_regNext_5_0_data_17;
  reg                 io_in_r_bypass_regNext_5_0_load_store_17;
  reg                 io_in_r_bypass_regNext_5_0_df_is_ws_17;
  reg                 io_in_r_bypass_regNext_5_0_stall_17;
  reg        [15:0]   io_in_r_bypass_regNext_5_1_data_17;
  reg                 io_in_r_bypass_regNext_5_1_load_store_17;
  reg                 io_in_r_bypass_regNext_5_1_df_is_ws_17;
  reg                 io_in_r_bypass_regNext_5_1_stall_17;
  reg        [15:0]   io_in_r_bypass_regNext_5_2_data_17;
  reg                 io_in_r_bypass_regNext_5_2_load_store_17;
  reg                 io_in_r_bypass_regNext_5_2_df_is_ws_17;
  reg                 io_in_r_bypass_regNext_5_2_stall_17;
  reg        [15:0]   io_in_r_bypass_regNext_5_3_data_17;
  reg                 io_in_r_bypass_regNext_5_3_load_store_17;
  reg                 io_in_r_bypass_regNext_5_3_df_is_ws_17;
  reg                 io_in_r_bypass_regNext_5_3_stall_17;
  reg        [15:0]   io_in_r_bypass_regNext_6_0_data_17;
  reg                 io_in_r_bypass_regNext_6_0_load_store_17;
  reg                 io_in_r_bypass_regNext_6_0_df_is_ws_17;
  reg                 io_in_r_bypass_regNext_6_0_stall_17;
  reg        [15:0]   io_in_r_bypass_regNext_6_1_data_17;
  reg                 io_in_r_bypass_regNext_6_1_load_store_17;
  reg                 io_in_r_bypass_regNext_6_1_df_is_ws_17;
  reg                 io_in_r_bypass_regNext_6_1_stall_17;
  reg        [15:0]   io_in_r_bypass_regNext_6_2_data_17;
  reg                 io_in_r_bypass_regNext_6_2_load_store_17;
  reg                 io_in_r_bypass_regNext_6_2_df_is_ws_17;
  reg                 io_in_r_bypass_regNext_6_2_stall_17;
  reg        [15:0]   io_in_r_bypass_regNext_6_3_data_17;
  reg                 io_in_r_bypass_regNext_6_3_load_store_17;
  reg                 io_in_r_bypass_regNext_6_3_df_is_ws_17;
  reg                 io_in_r_bypass_regNext_6_3_stall_17;
  reg        [15:0]   io_in_r_bypass_regNext_7_0_data_17;
  reg                 io_in_r_bypass_regNext_7_0_load_store_17;
  reg                 io_in_r_bypass_regNext_7_0_df_is_ws_17;
  reg                 io_in_r_bypass_regNext_7_0_stall_17;
  reg        [15:0]   io_in_r_bypass_regNext_7_1_data_17;
  reg                 io_in_r_bypass_regNext_7_1_load_store_17;
  reg                 io_in_r_bypass_regNext_7_1_df_is_ws_17;
  reg                 io_in_r_bypass_regNext_7_1_stall_17;
  reg        [15:0]   io_in_r_bypass_regNext_7_2_data_17;
  reg                 io_in_r_bypass_regNext_7_2_load_store_17;
  reg                 io_in_r_bypass_regNext_7_2_df_is_ws_17;
  reg                 io_in_r_bypass_regNext_7_2_stall_17;
  reg        [15:0]   io_in_r_bypass_regNext_7_3_data_17;
  reg                 io_in_r_bypass_regNext_7_3_load_store_17;
  reg                 io_in_r_bypass_regNext_7_3_df_is_ws_17;
  reg                 io_in_r_bypass_regNext_7_3_stall_17;
  reg        [15:0]   io_in_r_bypass_regNext_8_0_data_17;
  reg                 io_in_r_bypass_regNext_8_0_load_store_17;
  reg                 io_in_r_bypass_regNext_8_0_df_is_ws_17;
  reg                 io_in_r_bypass_regNext_8_0_stall_17;
  reg        [15:0]   io_in_r_bypass_regNext_8_1_data_17;
  reg                 io_in_r_bypass_regNext_8_1_load_store_17;
  reg                 io_in_r_bypass_regNext_8_1_df_is_ws_17;
  reg                 io_in_r_bypass_regNext_8_1_stall_17;
  reg        [15:0]   io_in_r_bypass_regNext_8_2_data_17;
  reg                 io_in_r_bypass_regNext_8_2_load_store_17;
  reg                 io_in_r_bypass_regNext_8_2_df_is_ws_17;
  reg                 io_in_r_bypass_regNext_8_2_stall_17;
  reg        [15:0]   io_in_r_bypass_regNext_8_3_data_17;
  reg                 io_in_r_bypass_regNext_8_3_load_store_17;
  reg                 io_in_r_bypass_regNext_8_3_df_is_ws_17;
  reg                 io_in_r_bypass_regNext_8_3_stall_17;
  reg        [15:0]   io_in_r_bypass_regNext_9_0_data_17;
  reg                 io_in_r_bypass_regNext_9_0_load_store_17;
  reg                 io_in_r_bypass_regNext_9_0_df_is_ws_17;
  reg                 io_in_r_bypass_regNext_9_0_stall_17;
  reg        [15:0]   io_in_r_bypass_regNext_9_1_data_17;
  reg                 io_in_r_bypass_regNext_9_1_load_store_17;
  reg                 io_in_r_bypass_regNext_9_1_df_is_ws_17;
  reg                 io_in_r_bypass_regNext_9_1_stall_17;
  reg        [15:0]   io_in_r_bypass_regNext_9_2_data_17;
  reg                 io_in_r_bypass_regNext_9_2_load_store_17;
  reg                 io_in_r_bypass_regNext_9_2_df_is_ws_17;
  reg                 io_in_r_bypass_regNext_9_2_stall_17;
  reg        [15:0]   io_in_r_bypass_regNext_9_3_data_17;
  reg                 io_in_r_bypass_regNext_9_3_load_store_17;
  reg                 io_in_r_bypass_regNext_9_3_df_is_ws_17;
  reg                 io_in_r_bypass_regNext_9_3_stall_17;
  reg        [15:0]   io_in_r_bypass_regNext_10_0_data_17;
  reg                 io_in_r_bypass_regNext_10_0_load_store_17;
  reg                 io_in_r_bypass_regNext_10_0_df_is_ws_17;
  reg                 io_in_r_bypass_regNext_10_0_stall_17;
  reg        [15:0]   io_in_r_bypass_regNext_10_1_data_17;
  reg                 io_in_r_bypass_regNext_10_1_load_store_17;
  reg                 io_in_r_bypass_regNext_10_1_df_is_ws_17;
  reg                 io_in_r_bypass_regNext_10_1_stall_17;
  reg        [15:0]   io_in_r_bypass_regNext_10_2_data_17;
  reg                 io_in_r_bypass_regNext_10_2_load_store_17;
  reg                 io_in_r_bypass_regNext_10_2_df_is_ws_17;
  reg                 io_in_r_bypass_regNext_10_2_stall_17;
  reg        [15:0]   io_in_r_bypass_regNext_10_3_data_17;
  reg                 io_in_r_bypass_regNext_10_3_load_store_17;
  reg                 io_in_r_bypass_regNext_10_3_df_is_ws_17;
  reg                 io_in_r_bypass_regNext_10_3_stall_17;
  reg        [15:0]   io_in_r_bypass_regNext_11_0_data_17;
  reg                 io_in_r_bypass_regNext_11_0_load_store_17;
  reg                 io_in_r_bypass_regNext_11_0_df_is_ws_17;
  reg                 io_in_r_bypass_regNext_11_0_stall_17;
  reg        [15:0]   io_in_r_bypass_regNext_11_1_data_17;
  reg                 io_in_r_bypass_regNext_11_1_load_store_17;
  reg                 io_in_r_bypass_regNext_11_1_df_is_ws_17;
  reg                 io_in_r_bypass_regNext_11_1_stall_17;
  reg        [15:0]   io_in_r_bypass_regNext_11_2_data_17;
  reg                 io_in_r_bypass_regNext_11_2_load_store_17;
  reg                 io_in_r_bypass_regNext_11_2_df_is_ws_17;
  reg                 io_in_r_bypass_regNext_11_2_stall_17;
  reg        [15:0]   io_in_r_bypass_regNext_11_3_data_17;
  reg                 io_in_r_bypass_regNext_11_3_load_store_17;
  reg                 io_in_r_bypass_regNext_11_3_df_is_ws_17;
  reg                 io_in_r_bypass_regNext_11_3_stall_17;
  reg        [15:0]   io_in_r_bypass_regNext_12_0_data_17;
  reg                 io_in_r_bypass_regNext_12_0_load_store_17;
  reg                 io_in_r_bypass_regNext_12_0_df_is_ws_17;
  reg                 io_in_r_bypass_regNext_12_0_stall_17;
  reg        [15:0]   io_in_r_bypass_regNext_12_1_data_17;
  reg                 io_in_r_bypass_regNext_12_1_load_store_17;
  reg                 io_in_r_bypass_regNext_12_1_df_is_ws_17;
  reg                 io_in_r_bypass_regNext_12_1_stall_17;
  reg        [15:0]   io_in_r_bypass_regNext_12_2_data_17;
  reg                 io_in_r_bypass_regNext_12_2_load_store_17;
  reg                 io_in_r_bypass_regNext_12_2_df_is_ws_17;
  reg                 io_in_r_bypass_regNext_12_2_stall_17;
  reg        [15:0]   io_in_r_bypass_regNext_12_3_data_17;
  reg                 io_in_r_bypass_regNext_12_3_load_store_17;
  reg                 io_in_r_bypass_regNext_12_3_df_is_ws_17;
  reg                 io_in_r_bypass_regNext_12_3_stall_17;
  reg        [15:0]   io_in_r_bypass_regNext_13_0_data_17;
  reg                 io_in_r_bypass_regNext_13_0_load_store_17;
  reg                 io_in_r_bypass_regNext_13_0_df_is_ws_17;
  reg                 io_in_r_bypass_regNext_13_0_stall_17;
  reg        [15:0]   io_in_r_bypass_regNext_13_1_data_17;
  reg                 io_in_r_bypass_regNext_13_1_load_store_17;
  reg                 io_in_r_bypass_regNext_13_1_df_is_ws_17;
  reg                 io_in_r_bypass_regNext_13_1_stall_17;
  reg        [15:0]   io_in_r_bypass_regNext_13_2_data_17;
  reg                 io_in_r_bypass_regNext_13_2_load_store_17;
  reg                 io_in_r_bypass_regNext_13_2_df_is_ws_17;
  reg                 io_in_r_bypass_regNext_13_2_stall_17;
  reg        [15:0]   io_in_r_bypass_regNext_13_3_data_17;
  reg                 io_in_r_bypass_regNext_13_3_load_store_17;
  reg                 io_in_r_bypass_regNext_13_3_df_is_ws_17;
  reg                 io_in_r_bypass_regNext_13_3_stall_17;
  reg        [15:0]   io_in_r_bypass_regNext_14_0_data_17;
  reg                 io_in_r_bypass_regNext_14_0_load_store_17;
  reg                 io_in_r_bypass_regNext_14_0_df_is_ws_17;
  reg                 io_in_r_bypass_regNext_14_0_stall_17;
  reg        [15:0]   io_in_r_bypass_regNext_14_1_data_17;
  reg                 io_in_r_bypass_regNext_14_1_load_store_17;
  reg                 io_in_r_bypass_regNext_14_1_df_is_ws_17;
  reg                 io_in_r_bypass_regNext_14_1_stall_17;
  reg        [15:0]   io_in_r_bypass_regNext_14_2_data_17;
  reg                 io_in_r_bypass_regNext_14_2_load_store_17;
  reg                 io_in_r_bypass_regNext_14_2_df_is_ws_17;
  reg                 io_in_r_bypass_regNext_14_2_stall_17;
  reg        [15:0]   io_in_r_bypass_regNext_14_3_data_17;
  reg                 io_in_r_bypass_regNext_14_3_load_store_17;
  reg                 io_in_r_bypass_regNext_14_3_df_is_ws_17;
  reg                 io_in_r_bypass_regNext_14_3_stall_17;
  reg        [15:0]   io_in_r_bypass_regNext_15_0_data_17;
  reg                 io_in_r_bypass_regNext_15_0_load_store_17;
  reg                 io_in_r_bypass_regNext_15_0_df_is_ws_17;
  reg                 io_in_r_bypass_regNext_15_0_stall_17;
  reg        [15:0]   io_in_r_bypass_regNext_15_1_data_17;
  reg                 io_in_r_bypass_regNext_15_1_load_store_17;
  reg                 io_in_r_bypass_regNext_15_1_df_is_ws_17;
  reg                 io_in_r_bypass_regNext_15_1_stall_17;
  reg        [15:0]   io_in_r_bypass_regNext_15_2_data_17;
  reg                 io_in_r_bypass_regNext_15_2_load_store_17;
  reg                 io_in_r_bypass_regNext_15_2_df_is_ws_17;
  reg                 io_in_r_bypass_regNext_15_2_stall_17;
  reg        [15:0]   io_in_r_bypass_regNext_15_3_data_17;
  reg                 io_in_r_bypass_regNext_15_3_load_store_17;
  reg                 io_in_r_bypass_regNext_15_3_df_is_ws_17;
  reg                 io_in_r_bypass_regNext_15_3_stall_17;
  reg        [15:0]   io_in_r_bypass_regNext_16_0_data_17;
  reg                 io_in_r_bypass_regNext_16_0_load_store_17;
  reg                 io_in_r_bypass_regNext_16_0_df_is_ws_17;
  reg                 io_in_r_bypass_regNext_16_0_stall_17;
  reg        [15:0]   io_in_r_bypass_regNext_16_1_data_17;
  reg                 io_in_r_bypass_regNext_16_1_load_store_17;
  reg                 io_in_r_bypass_regNext_16_1_df_is_ws_17;
  reg                 io_in_r_bypass_regNext_16_1_stall_17;
  reg        [15:0]   io_in_r_bypass_regNext_16_2_data_17;
  reg                 io_in_r_bypass_regNext_16_2_load_store_17;
  reg                 io_in_r_bypass_regNext_16_2_df_is_ws_17;
  reg                 io_in_r_bypass_regNext_16_2_stall_17;
  reg        [15:0]   io_in_r_bypass_regNext_16_3_data_17;
  reg                 io_in_r_bypass_regNext_16_3_load_store_17;
  reg                 io_in_r_bypass_regNext_16_3_df_is_ws_17;
  reg                 io_in_r_bypass_regNext_16_3_stall_17;
  reg        [15:0]   io_in_r_bypass_regNext_17_0_data_17;
  reg                 io_in_r_bypass_regNext_17_0_load_store_17;
  reg                 io_in_r_bypass_regNext_17_0_df_is_ws_17;
  reg                 io_in_r_bypass_regNext_17_0_stall_17;
  reg        [15:0]   io_in_r_bypass_regNext_17_1_data_17;
  reg                 io_in_r_bypass_regNext_17_1_load_store_17;
  reg                 io_in_r_bypass_regNext_17_1_df_is_ws_17;
  reg                 io_in_r_bypass_regNext_17_1_stall_17;
  reg        [15:0]   io_in_r_bypass_regNext_17_2_data_17;
  reg                 io_in_r_bypass_regNext_17_2_load_store_17;
  reg                 io_in_r_bypass_regNext_17_2_df_is_ws_17;
  reg                 io_in_r_bypass_regNext_17_2_stall_17;
  reg        [15:0]   io_in_r_bypass_regNext_17_3_data_17;
  reg                 io_in_r_bypass_regNext_17_3_load_store_17;
  reg                 io_in_r_bypass_regNext_17_3_df_is_ws_17;
  reg                 io_in_r_bypass_regNext_17_3_stall_17;
  reg        [15:0]   io_in_r_bypass_regNext_18_0_data_17;
  reg                 io_in_r_bypass_regNext_18_0_load_store_17;
  reg                 io_in_r_bypass_regNext_18_0_df_is_ws_17;
  reg                 io_in_r_bypass_regNext_18_0_stall_17;
  reg        [15:0]   io_in_r_bypass_regNext_18_1_data_17;
  reg                 io_in_r_bypass_regNext_18_1_load_store_17;
  reg                 io_in_r_bypass_regNext_18_1_df_is_ws_17;
  reg                 io_in_r_bypass_regNext_18_1_stall_17;
  reg        [15:0]   io_in_r_bypass_regNext_18_2_data_17;
  reg                 io_in_r_bypass_regNext_18_2_load_store_17;
  reg                 io_in_r_bypass_regNext_18_2_df_is_ws_17;
  reg                 io_in_r_bypass_regNext_18_2_stall_17;
  reg        [15:0]   io_in_r_bypass_regNext_18_3_data_17;
  reg                 io_in_r_bypass_regNext_18_3_load_store_17;
  reg                 io_in_r_bypass_regNext_18_3_df_is_ws_17;
  reg                 io_in_r_bypass_regNext_18_3_stall_17;
  reg        [15:0]   io_in_r_bypass_regNext_19_0_data_17;
  reg                 io_in_r_bypass_regNext_19_0_load_store_17;
  reg                 io_in_r_bypass_regNext_19_0_df_is_ws_17;
  reg                 io_in_r_bypass_regNext_19_0_stall_17;
  reg        [15:0]   io_in_r_bypass_regNext_19_1_data_17;
  reg                 io_in_r_bypass_regNext_19_1_load_store_17;
  reg                 io_in_r_bypass_regNext_19_1_df_is_ws_17;
  reg                 io_in_r_bypass_regNext_19_1_stall_17;
  reg        [15:0]   io_in_r_bypass_regNext_19_2_data_17;
  reg                 io_in_r_bypass_regNext_19_2_load_store_17;
  reg                 io_in_r_bypass_regNext_19_2_df_is_ws_17;
  reg                 io_in_r_bypass_regNext_19_2_stall_17;
  reg        [15:0]   io_in_r_bypass_regNext_19_3_data_17;
  reg                 io_in_r_bypass_regNext_19_3_load_store_17;
  reg                 io_in_r_bypass_regNext_19_3_df_is_ws_17;
  reg                 io_in_r_bypass_regNext_19_3_stall_17;
  reg        [15:0]   io_in_r_bypass_regNext_20_0_data_17;
  reg                 io_in_r_bypass_regNext_20_0_load_store_17;
  reg                 io_in_r_bypass_regNext_20_0_df_is_ws_17;
  reg                 io_in_r_bypass_regNext_20_0_stall_17;
  reg        [15:0]   io_in_r_bypass_regNext_20_1_data_17;
  reg                 io_in_r_bypass_regNext_20_1_load_store_17;
  reg                 io_in_r_bypass_regNext_20_1_df_is_ws_17;
  reg                 io_in_r_bypass_regNext_20_1_stall_17;
  reg        [15:0]   io_in_r_bypass_regNext_20_2_data_17;
  reg                 io_in_r_bypass_regNext_20_2_load_store_17;
  reg                 io_in_r_bypass_regNext_20_2_df_is_ws_17;
  reg                 io_in_r_bypass_regNext_20_2_stall_17;
  reg        [15:0]   io_in_r_bypass_regNext_20_3_data_17;
  reg                 io_in_r_bypass_regNext_20_3_load_store_17;
  reg                 io_in_r_bypass_regNext_20_3_df_is_ws_17;
  reg                 io_in_r_bypass_regNext_20_3_stall_17;
  reg        [15:0]   io_in_r_bypass_regNext_21_0_data_17;
  reg                 io_in_r_bypass_regNext_21_0_load_store_17;
  reg                 io_in_r_bypass_regNext_21_0_df_is_ws_17;
  reg                 io_in_r_bypass_regNext_21_0_stall_17;
  reg        [15:0]   io_in_r_bypass_regNext_21_1_data_17;
  reg                 io_in_r_bypass_regNext_21_1_load_store_17;
  reg                 io_in_r_bypass_regNext_21_1_df_is_ws_17;
  reg                 io_in_r_bypass_regNext_21_1_stall_17;
  reg        [15:0]   io_in_r_bypass_regNext_21_2_data_17;
  reg                 io_in_r_bypass_regNext_21_2_load_store_17;
  reg                 io_in_r_bypass_regNext_21_2_df_is_ws_17;
  reg                 io_in_r_bypass_regNext_21_2_stall_17;
  reg        [15:0]   io_in_r_bypass_regNext_21_3_data_17;
  reg                 io_in_r_bypass_regNext_21_3_load_store_17;
  reg                 io_in_r_bypass_regNext_21_3_df_is_ws_17;
  reg                 io_in_r_bypass_regNext_21_3_stall_17;
  reg        [15:0]   io_in_r_bypass_regNext_22_0_data_17;
  reg                 io_in_r_bypass_regNext_22_0_load_store_17;
  reg                 io_in_r_bypass_regNext_22_0_df_is_ws_17;
  reg                 io_in_r_bypass_regNext_22_0_stall_17;
  reg        [15:0]   io_in_r_bypass_regNext_22_1_data_17;
  reg                 io_in_r_bypass_regNext_22_1_load_store_17;
  reg                 io_in_r_bypass_regNext_22_1_df_is_ws_17;
  reg                 io_in_r_bypass_regNext_22_1_stall_17;
  reg        [15:0]   io_in_r_bypass_regNext_22_2_data_17;
  reg                 io_in_r_bypass_regNext_22_2_load_store_17;
  reg                 io_in_r_bypass_regNext_22_2_df_is_ws_17;
  reg                 io_in_r_bypass_regNext_22_2_stall_17;
  reg        [15:0]   io_in_r_bypass_regNext_22_3_data_17;
  reg                 io_in_r_bypass_regNext_22_3_load_store_17;
  reg                 io_in_r_bypass_regNext_22_3_df_is_ws_17;
  reg                 io_in_r_bypass_regNext_22_3_stall_17;
  reg        [15:0]   io_in_r_bypass_regNext_23_0_data_17;
  reg                 io_in_r_bypass_regNext_23_0_load_store_17;
  reg                 io_in_r_bypass_regNext_23_0_df_is_ws_17;
  reg                 io_in_r_bypass_regNext_23_0_stall_17;
  reg        [15:0]   io_in_r_bypass_regNext_23_1_data_17;
  reg                 io_in_r_bypass_regNext_23_1_load_store_17;
  reg                 io_in_r_bypass_regNext_23_1_df_is_ws_17;
  reg                 io_in_r_bypass_regNext_23_1_stall_17;
  reg        [15:0]   io_in_r_bypass_regNext_23_2_data_17;
  reg                 io_in_r_bypass_regNext_23_2_load_store_17;
  reg                 io_in_r_bypass_regNext_23_2_df_is_ws_17;
  reg                 io_in_r_bypass_regNext_23_2_stall_17;
  reg        [15:0]   io_in_r_bypass_regNext_23_3_data_17;
  reg                 io_in_r_bypass_regNext_23_3_load_store_17;
  reg                 io_in_r_bypass_regNext_23_3_df_is_ws_17;
  reg                 io_in_r_bypass_regNext_23_3_stall_17;
  reg        [15:0]   io_in_r_bypass_regNext_24_0_data_17;
  reg                 io_in_r_bypass_regNext_24_0_load_store_17;
  reg                 io_in_r_bypass_regNext_24_0_df_is_ws_17;
  reg                 io_in_r_bypass_regNext_24_0_stall_17;
  reg        [15:0]   io_in_r_bypass_regNext_24_1_data_17;
  reg                 io_in_r_bypass_regNext_24_1_load_store_17;
  reg                 io_in_r_bypass_regNext_24_1_df_is_ws_17;
  reg                 io_in_r_bypass_regNext_24_1_stall_17;
  reg        [15:0]   io_in_r_bypass_regNext_24_2_data_17;
  reg                 io_in_r_bypass_regNext_24_2_load_store_17;
  reg                 io_in_r_bypass_regNext_24_2_df_is_ws_17;
  reg                 io_in_r_bypass_regNext_24_2_stall_17;
  reg        [15:0]   io_in_r_bypass_regNext_24_3_data_17;
  reg                 io_in_r_bypass_regNext_24_3_load_store_17;
  reg                 io_in_r_bypass_regNext_24_3_df_is_ws_17;
  reg                 io_in_r_bypass_regNext_24_3_stall_17;
  reg        [15:0]   io_in_r_bypass_regNext_25_0_data_17;
  reg                 io_in_r_bypass_regNext_25_0_load_store_17;
  reg                 io_in_r_bypass_regNext_25_0_df_is_ws_17;
  reg                 io_in_r_bypass_regNext_25_0_stall_17;
  reg        [15:0]   io_in_r_bypass_regNext_25_1_data_17;
  reg                 io_in_r_bypass_regNext_25_1_load_store_17;
  reg                 io_in_r_bypass_regNext_25_1_df_is_ws_17;
  reg                 io_in_r_bypass_regNext_25_1_stall_17;
  reg        [15:0]   io_in_r_bypass_regNext_25_2_data_17;
  reg                 io_in_r_bypass_regNext_25_2_load_store_17;
  reg                 io_in_r_bypass_regNext_25_2_df_is_ws_17;
  reg                 io_in_r_bypass_regNext_25_2_stall_17;
  reg        [15:0]   io_in_r_bypass_regNext_25_3_data_17;
  reg                 io_in_r_bypass_regNext_25_3_load_store_17;
  reg                 io_in_r_bypass_regNext_25_3_df_is_ws_17;
  reg                 io_in_r_bypass_regNext_25_3_stall_17;
  reg        [15:0]   io_in_r_bypass_regNext_26_0_data_17;
  reg                 io_in_r_bypass_regNext_26_0_load_store_17;
  reg                 io_in_r_bypass_regNext_26_0_df_is_ws_17;
  reg                 io_in_r_bypass_regNext_26_0_stall_17;
  reg        [15:0]   io_in_r_bypass_regNext_26_1_data_17;
  reg                 io_in_r_bypass_regNext_26_1_load_store_17;
  reg                 io_in_r_bypass_regNext_26_1_df_is_ws_17;
  reg                 io_in_r_bypass_regNext_26_1_stall_17;
  reg        [15:0]   io_in_r_bypass_regNext_26_2_data_17;
  reg                 io_in_r_bypass_regNext_26_2_load_store_17;
  reg                 io_in_r_bypass_regNext_26_2_df_is_ws_17;
  reg                 io_in_r_bypass_regNext_26_2_stall_17;
  reg        [15:0]   io_in_r_bypass_regNext_26_3_data_17;
  reg                 io_in_r_bypass_regNext_26_3_load_store_17;
  reg                 io_in_r_bypass_regNext_26_3_df_is_ws_17;
  reg                 io_in_r_bypass_regNext_26_3_stall_17;
  reg        [15:0]   io_in_r_bypass_regNext_27_0_data_17;
  reg                 io_in_r_bypass_regNext_27_0_load_store_17;
  reg                 io_in_r_bypass_regNext_27_0_df_is_ws_17;
  reg                 io_in_r_bypass_regNext_27_0_stall_17;
  reg        [15:0]   io_in_r_bypass_regNext_27_1_data_17;
  reg                 io_in_r_bypass_regNext_27_1_load_store_17;
  reg                 io_in_r_bypass_regNext_27_1_df_is_ws_17;
  reg                 io_in_r_bypass_regNext_27_1_stall_17;
  reg        [15:0]   io_in_r_bypass_regNext_27_2_data_17;
  reg                 io_in_r_bypass_regNext_27_2_load_store_17;
  reg                 io_in_r_bypass_regNext_27_2_df_is_ws_17;
  reg                 io_in_r_bypass_regNext_27_2_stall_17;
  reg        [15:0]   io_in_r_bypass_regNext_27_3_data_17;
  reg                 io_in_r_bypass_regNext_27_3_load_store_17;
  reg                 io_in_r_bypass_regNext_27_3_df_is_ws_17;
  reg                 io_in_r_bypass_regNext_27_3_stall_17;
  reg        [15:0]   io_in_r_bypass_regNext_28_0_data_17;
  reg                 io_in_r_bypass_regNext_28_0_load_store_17;
  reg                 io_in_r_bypass_regNext_28_0_df_is_ws_17;
  reg                 io_in_r_bypass_regNext_28_0_stall_17;
  reg        [15:0]   io_in_r_bypass_regNext_28_1_data_17;
  reg                 io_in_r_bypass_regNext_28_1_load_store_17;
  reg                 io_in_r_bypass_regNext_28_1_df_is_ws_17;
  reg                 io_in_r_bypass_regNext_28_1_stall_17;
  reg        [15:0]   io_in_r_bypass_regNext_28_2_data_17;
  reg                 io_in_r_bypass_regNext_28_2_load_store_17;
  reg                 io_in_r_bypass_regNext_28_2_df_is_ws_17;
  reg                 io_in_r_bypass_regNext_28_2_stall_17;
  reg        [15:0]   io_in_r_bypass_regNext_28_3_data_17;
  reg                 io_in_r_bypass_regNext_28_3_load_store_17;
  reg                 io_in_r_bypass_regNext_28_3_df_is_ws_17;
  reg                 io_in_r_bypass_regNext_28_3_stall_17;
  reg        [15:0]   io_in_r_bypass_regNext_29_0_data_17;
  reg                 io_in_r_bypass_regNext_29_0_load_store_17;
  reg                 io_in_r_bypass_regNext_29_0_df_is_ws_17;
  reg                 io_in_r_bypass_regNext_29_0_stall_17;
  reg        [15:0]   io_in_r_bypass_regNext_29_1_data_17;
  reg                 io_in_r_bypass_regNext_29_1_load_store_17;
  reg                 io_in_r_bypass_regNext_29_1_df_is_ws_17;
  reg                 io_in_r_bypass_regNext_29_1_stall_17;
  reg        [15:0]   io_in_r_bypass_regNext_29_2_data_17;
  reg                 io_in_r_bypass_regNext_29_2_load_store_17;
  reg                 io_in_r_bypass_regNext_29_2_df_is_ws_17;
  reg                 io_in_r_bypass_regNext_29_2_stall_17;
  reg        [15:0]   io_in_r_bypass_regNext_29_3_data_17;
  reg                 io_in_r_bypass_regNext_29_3_load_store_17;
  reg                 io_in_r_bypass_regNext_29_3_df_is_ws_17;
  reg                 io_in_r_bypass_regNext_29_3_stall_17;
  reg        [15:0]   io_in_r_bypass_regNext_30_0_data_17;
  reg                 io_in_r_bypass_regNext_30_0_load_store_17;
  reg                 io_in_r_bypass_regNext_30_0_df_is_ws_17;
  reg                 io_in_r_bypass_regNext_30_0_stall_17;
  reg        [15:0]   io_in_r_bypass_regNext_30_1_data_17;
  reg                 io_in_r_bypass_regNext_30_1_load_store_17;
  reg                 io_in_r_bypass_regNext_30_1_df_is_ws_17;
  reg                 io_in_r_bypass_regNext_30_1_stall_17;
  reg        [15:0]   io_in_r_bypass_regNext_30_2_data_17;
  reg                 io_in_r_bypass_regNext_30_2_load_store_17;
  reg                 io_in_r_bypass_regNext_30_2_df_is_ws_17;
  reg                 io_in_r_bypass_regNext_30_2_stall_17;
  reg        [15:0]   io_in_r_bypass_regNext_30_3_data_17;
  reg                 io_in_r_bypass_regNext_30_3_load_store_17;
  reg                 io_in_r_bypass_regNext_30_3_df_is_ws_17;
  reg                 io_in_r_bypass_regNext_30_3_stall_17;
  reg        [15:0]   io_in_r_bypass_regNext_31_0_data_17;
  reg                 io_in_r_bypass_regNext_31_0_load_store_17;
  reg                 io_in_r_bypass_regNext_31_0_df_is_ws_17;
  reg                 io_in_r_bypass_regNext_31_0_stall_17;
  reg        [15:0]   io_in_r_bypass_regNext_31_1_data_17;
  reg                 io_in_r_bypass_regNext_31_1_load_store_17;
  reg                 io_in_r_bypass_regNext_31_1_df_is_ws_17;
  reg                 io_in_r_bypass_regNext_31_1_stall_17;
  reg        [15:0]   io_in_r_bypass_regNext_31_2_data_17;
  reg                 io_in_r_bypass_regNext_31_2_load_store_17;
  reg                 io_in_r_bypass_regNext_31_2_df_is_ws_17;
  reg                 io_in_r_bypass_regNext_31_2_stall_17;
  reg        [15:0]   io_in_r_bypass_regNext_31_3_data_17;
  reg                 io_in_r_bypass_regNext_31_3_load_store_17;
  reg                 io_in_r_bypass_regNext_31_3_df_is_ws_17;
  reg                 io_in_r_bypass_regNext_31_3_stall_17;
  reg        [15:0]   io_in_r_bypass_regNext_0_0_data_18;
  reg                 io_in_r_bypass_regNext_0_0_load_store_18;
  reg                 io_in_r_bypass_regNext_0_0_df_is_ws_18;
  reg                 io_in_r_bypass_regNext_0_0_stall_18;
  reg        [15:0]   io_in_r_bypass_regNext_0_1_data_18;
  reg                 io_in_r_bypass_regNext_0_1_load_store_18;
  reg                 io_in_r_bypass_regNext_0_1_df_is_ws_18;
  reg                 io_in_r_bypass_regNext_0_1_stall_18;
  reg        [15:0]   io_in_r_bypass_regNext_0_2_data_18;
  reg                 io_in_r_bypass_regNext_0_2_load_store_18;
  reg                 io_in_r_bypass_regNext_0_2_df_is_ws_18;
  reg                 io_in_r_bypass_regNext_0_2_stall_18;
  reg        [15:0]   io_in_r_bypass_regNext_0_3_data_18;
  reg                 io_in_r_bypass_regNext_0_3_load_store_18;
  reg                 io_in_r_bypass_regNext_0_3_df_is_ws_18;
  reg                 io_in_r_bypass_regNext_0_3_stall_18;
  reg        [15:0]   io_in_r_bypass_regNext_1_0_data_18;
  reg                 io_in_r_bypass_regNext_1_0_load_store_18;
  reg                 io_in_r_bypass_regNext_1_0_df_is_ws_18;
  reg                 io_in_r_bypass_regNext_1_0_stall_18;
  reg        [15:0]   io_in_r_bypass_regNext_1_1_data_18;
  reg                 io_in_r_bypass_regNext_1_1_load_store_18;
  reg                 io_in_r_bypass_regNext_1_1_df_is_ws_18;
  reg                 io_in_r_bypass_regNext_1_1_stall_18;
  reg        [15:0]   io_in_r_bypass_regNext_1_2_data_18;
  reg                 io_in_r_bypass_regNext_1_2_load_store_18;
  reg                 io_in_r_bypass_regNext_1_2_df_is_ws_18;
  reg                 io_in_r_bypass_regNext_1_2_stall_18;
  reg        [15:0]   io_in_r_bypass_regNext_1_3_data_18;
  reg                 io_in_r_bypass_regNext_1_3_load_store_18;
  reg                 io_in_r_bypass_regNext_1_3_df_is_ws_18;
  reg                 io_in_r_bypass_regNext_1_3_stall_18;
  reg        [15:0]   io_in_r_bypass_regNext_2_0_data_18;
  reg                 io_in_r_bypass_regNext_2_0_load_store_18;
  reg                 io_in_r_bypass_regNext_2_0_df_is_ws_18;
  reg                 io_in_r_bypass_regNext_2_0_stall_18;
  reg        [15:0]   io_in_r_bypass_regNext_2_1_data_18;
  reg                 io_in_r_bypass_regNext_2_1_load_store_18;
  reg                 io_in_r_bypass_regNext_2_1_df_is_ws_18;
  reg                 io_in_r_bypass_regNext_2_1_stall_18;
  reg        [15:0]   io_in_r_bypass_regNext_2_2_data_18;
  reg                 io_in_r_bypass_regNext_2_2_load_store_18;
  reg                 io_in_r_bypass_regNext_2_2_df_is_ws_18;
  reg                 io_in_r_bypass_regNext_2_2_stall_18;
  reg        [15:0]   io_in_r_bypass_regNext_2_3_data_18;
  reg                 io_in_r_bypass_regNext_2_3_load_store_18;
  reg                 io_in_r_bypass_regNext_2_3_df_is_ws_18;
  reg                 io_in_r_bypass_regNext_2_3_stall_18;
  reg        [15:0]   io_in_r_bypass_regNext_3_0_data_18;
  reg                 io_in_r_bypass_regNext_3_0_load_store_18;
  reg                 io_in_r_bypass_regNext_3_0_df_is_ws_18;
  reg                 io_in_r_bypass_regNext_3_0_stall_18;
  reg        [15:0]   io_in_r_bypass_regNext_3_1_data_18;
  reg                 io_in_r_bypass_regNext_3_1_load_store_18;
  reg                 io_in_r_bypass_regNext_3_1_df_is_ws_18;
  reg                 io_in_r_bypass_regNext_3_1_stall_18;
  reg        [15:0]   io_in_r_bypass_regNext_3_2_data_18;
  reg                 io_in_r_bypass_regNext_3_2_load_store_18;
  reg                 io_in_r_bypass_regNext_3_2_df_is_ws_18;
  reg                 io_in_r_bypass_regNext_3_2_stall_18;
  reg        [15:0]   io_in_r_bypass_regNext_3_3_data_18;
  reg                 io_in_r_bypass_regNext_3_3_load_store_18;
  reg                 io_in_r_bypass_regNext_3_3_df_is_ws_18;
  reg                 io_in_r_bypass_regNext_3_3_stall_18;
  reg        [15:0]   io_in_r_bypass_regNext_4_0_data_18;
  reg                 io_in_r_bypass_regNext_4_0_load_store_18;
  reg                 io_in_r_bypass_regNext_4_0_df_is_ws_18;
  reg                 io_in_r_bypass_regNext_4_0_stall_18;
  reg        [15:0]   io_in_r_bypass_regNext_4_1_data_18;
  reg                 io_in_r_bypass_regNext_4_1_load_store_18;
  reg                 io_in_r_bypass_regNext_4_1_df_is_ws_18;
  reg                 io_in_r_bypass_regNext_4_1_stall_18;
  reg        [15:0]   io_in_r_bypass_regNext_4_2_data_18;
  reg                 io_in_r_bypass_regNext_4_2_load_store_18;
  reg                 io_in_r_bypass_regNext_4_2_df_is_ws_18;
  reg                 io_in_r_bypass_regNext_4_2_stall_18;
  reg        [15:0]   io_in_r_bypass_regNext_4_3_data_18;
  reg                 io_in_r_bypass_regNext_4_3_load_store_18;
  reg                 io_in_r_bypass_regNext_4_3_df_is_ws_18;
  reg                 io_in_r_bypass_regNext_4_3_stall_18;
  reg        [15:0]   io_in_r_bypass_regNext_5_0_data_18;
  reg                 io_in_r_bypass_regNext_5_0_load_store_18;
  reg                 io_in_r_bypass_regNext_5_0_df_is_ws_18;
  reg                 io_in_r_bypass_regNext_5_0_stall_18;
  reg        [15:0]   io_in_r_bypass_regNext_5_1_data_18;
  reg                 io_in_r_bypass_regNext_5_1_load_store_18;
  reg                 io_in_r_bypass_regNext_5_1_df_is_ws_18;
  reg                 io_in_r_bypass_regNext_5_1_stall_18;
  reg        [15:0]   io_in_r_bypass_regNext_5_2_data_18;
  reg                 io_in_r_bypass_regNext_5_2_load_store_18;
  reg                 io_in_r_bypass_regNext_5_2_df_is_ws_18;
  reg                 io_in_r_bypass_regNext_5_2_stall_18;
  reg        [15:0]   io_in_r_bypass_regNext_5_3_data_18;
  reg                 io_in_r_bypass_regNext_5_3_load_store_18;
  reg                 io_in_r_bypass_regNext_5_3_df_is_ws_18;
  reg                 io_in_r_bypass_regNext_5_3_stall_18;
  reg        [15:0]   io_in_r_bypass_regNext_6_0_data_18;
  reg                 io_in_r_bypass_regNext_6_0_load_store_18;
  reg                 io_in_r_bypass_regNext_6_0_df_is_ws_18;
  reg                 io_in_r_bypass_regNext_6_0_stall_18;
  reg        [15:0]   io_in_r_bypass_regNext_6_1_data_18;
  reg                 io_in_r_bypass_regNext_6_1_load_store_18;
  reg                 io_in_r_bypass_regNext_6_1_df_is_ws_18;
  reg                 io_in_r_bypass_regNext_6_1_stall_18;
  reg        [15:0]   io_in_r_bypass_regNext_6_2_data_18;
  reg                 io_in_r_bypass_regNext_6_2_load_store_18;
  reg                 io_in_r_bypass_regNext_6_2_df_is_ws_18;
  reg                 io_in_r_bypass_regNext_6_2_stall_18;
  reg        [15:0]   io_in_r_bypass_regNext_6_3_data_18;
  reg                 io_in_r_bypass_regNext_6_3_load_store_18;
  reg                 io_in_r_bypass_regNext_6_3_df_is_ws_18;
  reg                 io_in_r_bypass_regNext_6_3_stall_18;
  reg        [15:0]   io_in_r_bypass_regNext_7_0_data_18;
  reg                 io_in_r_bypass_regNext_7_0_load_store_18;
  reg                 io_in_r_bypass_regNext_7_0_df_is_ws_18;
  reg                 io_in_r_bypass_regNext_7_0_stall_18;
  reg        [15:0]   io_in_r_bypass_regNext_7_1_data_18;
  reg                 io_in_r_bypass_regNext_7_1_load_store_18;
  reg                 io_in_r_bypass_regNext_7_1_df_is_ws_18;
  reg                 io_in_r_bypass_regNext_7_1_stall_18;
  reg        [15:0]   io_in_r_bypass_regNext_7_2_data_18;
  reg                 io_in_r_bypass_regNext_7_2_load_store_18;
  reg                 io_in_r_bypass_regNext_7_2_df_is_ws_18;
  reg                 io_in_r_bypass_regNext_7_2_stall_18;
  reg        [15:0]   io_in_r_bypass_regNext_7_3_data_18;
  reg                 io_in_r_bypass_regNext_7_3_load_store_18;
  reg                 io_in_r_bypass_regNext_7_3_df_is_ws_18;
  reg                 io_in_r_bypass_regNext_7_3_stall_18;
  reg        [15:0]   io_in_r_bypass_regNext_8_0_data_18;
  reg                 io_in_r_bypass_regNext_8_0_load_store_18;
  reg                 io_in_r_bypass_regNext_8_0_df_is_ws_18;
  reg                 io_in_r_bypass_regNext_8_0_stall_18;
  reg        [15:0]   io_in_r_bypass_regNext_8_1_data_18;
  reg                 io_in_r_bypass_regNext_8_1_load_store_18;
  reg                 io_in_r_bypass_regNext_8_1_df_is_ws_18;
  reg                 io_in_r_bypass_regNext_8_1_stall_18;
  reg        [15:0]   io_in_r_bypass_regNext_8_2_data_18;
  reg                 io_in_r_bypass_regNext_8_2_load_store_18;
  reg                 io_in_r_bypass_regNext_8_2_df_is_ws_18;
  reg                 io_in_r_bypass_regNext_8_2_stall_18;
  reg        [15:0]   io_in_r_bypass_regNext_8_3_data_18;
  reg                 io_in_r_bypass_regNext_8_3_load_store_18;
  reg                 io_in_r_bypass_regNext_8_3_df_is_ws_18;
  reg                 io_in_r_bypass_regNext_8_3_stall_18;
  reg        [15:0]   io_in_r_bypass_regNext_9_0_data_18;
  reg                 io_in_r_bypass_regNext_9_0_load_store_18;
  reg                 io_in_r_bypass_regNext_9_0_df_is_ws_18;
  reg                 io_in_r_bypass_regNext_9_0_stall_18;
  reg        [15:0]   io_in_r_bypass_regNext_9_1_data_18;
  reg                 io_in_r_bypass_regNext_9_1_load_store_18;
  reg                 io_in_r_bypass_regNext_9_1_df_is_ws_18;
  reg                 io_in_r_bypass_regNext_9_1_stall_18;
  reg        [15:0]   io_in_r_bypass_regNext_9_2_data_18;
  reg                 io_in_r_bypass_regNext_9_2_load_store_18;
  reg                 io_in_r_bypass_regNext_9_2_df_is_ws_18;
  reg                 io_in_r_bypass_regNext_9_2_stall_18;
  reg        [15:0]   io_in_r_bypass_regNext_9_3_data_18;
  reg                 io_in_r_bypass_regNext_9_3_load_store_18;
  reg                 io_in_r_bypass_regNext_9_3_df_is_ws_18;
  reg                 io_in_r_bypass_regNext_9_3_stall_18;
  reg        [15:0]   io_in_r_bypass_regNext_10_0_data_18;
  reg                 io_in_r_bypass_regNext_10_0_load_store_18;
  reg                 io_in_r_bypass_regNext_10_0_df_is_ws_18;
  reg                 io_in_r_bypass_regNext_10_0_stall_18;
  reg        [15:0]   io_in_r_bypass_regNext_10_1_data_18;
  reg                 io_in_r_bypass_regNext_10_1_load_store_18;
  reg                 io_in_r_bypass_regNext_10_1_df_is_ws_18;
  reg                 io_in_r_bypass_regNext_10_1_stall_18;
  reg        [15:0]   io_in_r_bypass_regNext_10_2_data_18;
  reg                 io_in_r_bypass_regNext_10_2_load_store_18;
  reg                 io_in_r_bypass_regNext_10_2_df_is_ws_18;
  reg                 io_in_r_bypass_regNext_10_2_stall_18;
  reg        [15:0]   io_in_r_bypass_regNext_10_3_data_18;
  reg                 io_in_r_bypass_regNext_10_3_load_store_18;
  reg                 io_in_r_bypass_regNext_10_3_df_is_ws_18;
  reg                 io_in_r_bypass_regNext_10_3_stall_18;
  reg        [15:0]   io_in_r_bypass_regNext_11_0_data_18;
  reg                 io_in_r_bypass_regNext_11_0_load_store_18;
  reg                 io_in_r_bypass_regNext_11_0_df_is_ws_18;
  reg                 io_in_r_bypass_regNext_11_0_stall_18;
  reg        [15:0]   io_in_r_bypass_regNext_11_1_data_18;
  reg                 io_in_r_bypass_regNext_11_1_load_store_18;
  reg                 io_in_r_bypass_regNext_11_1_df_is_ws_18;
  reg                 io_in_r_bypass_regNext_11_1_stall_18;
  reg        [15:0]   io_in_r_bypass_regNext_11_2_data_18;
  reg                 io_in_r_bypass_regNext_11_2_load_store_18;
  reg                 io_in_r_bypass_regNext_11_2_df_is_ws_18;
  reg                 io_in_r_bypass_regNext_11_2_stall_18;
  reg        [15:0]   io_in_r_bypass_regNext_11_3_data_18;
  reg                 io_in_r_bypass_regNext_11_3_load_store_18;
  reg                 io_in_r_bypass_regNext_11_3_df_is_ws_18;
  reg                 io_in_r_bypass_regNext_11_3_stall_18;
  reg        [15:0]   io_in_r_bypass_regNext_12_0_data_18;
  reg                 io_in_r_bypass_regNext_12_0_load_store_18;
  reg                 io_in_r_bypass_regNext_12_0_df_is_ws_18;
  reg                 io_in_r_bypass_regNext_12_0_stall_18;
  reg        [15:0]   io_in_r_bypass_regNext_12_1_data_18;
  reg                 io_in_r_bypass_regNext_12_1_load_store_18;
  reg                 io_in_r_bypass_regNext_12_1_df_is_ws_18;
  reg                 io_in_r_bypass_regNext_12_1_stall_18;
  reg        [15:0]   io_in_r_bypass_regNext_12_2_data_18;
  reg                 io_in_r_bypass_regNext_12_2_load_store_18;
  reg                 io_in_r_bypass_regNext_12_2_df_is_ws_18;
  reg                 io_in_r_bypass_regNext_12_2_stall_18;
  reg        [15:0]   io_in_r_bypass_regNext_12_3_data_18;
  reg                 io_in_r_bypass_regNext_12_3_load_store_18;
  reg                 io_in_r_bypass_regNext_12_3_df_is_ws_18;
  reg                 io_in_r_bypass_regNext_12_3_stall_18;
  reg        [15:0]   io_in_r_bypass_regNext_13_0_data_18;
  reg                 io_in_r_bypass_regNext_13_0_load_store_18;
  reg                 io_in_r_bypass_regNext_13_0_df_is_ws_18;
  reg                 io_in_r_bypass_regNext_13_0_stall_18;
  reg        [15:0]   io_in_r_bypass_regNext_13_1_data_18;
  reg                 io_in_r_bypass_regNext_13_1_load_store_18;
  reg                 io_in_r_bypass_regNext_13_1_df_is_ws_18;
  reg                 io_in_r_bypass_regNext_13_1_stall_18;
  reg        [15:0]   io_in_r_bypass_regNext_13_2_data_18;
  reg                 io_in_r_bypass_regNext_13_2_load_store_18;
  reg                 io_in_r_bypass_regNext_13_2_df_is_ws_18;
  reg                 io_in_r_bypass_regNext_13_2_stall_18;
  reg        [15:0]   io_in_r_bypass_regNext_13_3_data_18;
  reg                 io_in_r_bypass_regNext_13_3_load_store_18;
  reg                 io_in_r_bypass_regNext_13_3_df_is_ws_18;
  reg                 io_in_r_bypass_regNext_13_3_stall_18;
  reg        [15:0]   io_in_r_bypass_regNext_14_0_data_18;
  reg                 io_in_r_bypass_regNext_14_0_load_store_18;
  reg                 io_in_r_bypass_regNext_14_0_df_is_ws_18;
  reg                 io_in_r_bypass_regNext_14_0_stall_18;
  reg        [15:0]   io_in_r_bypass_regNext_14_1_data_18;
  reg                 io_in_r_bypass_regNext_14_1_load_store_18;
  reg                 io_in_r_bypass_regNext_14_1_df_is_ws_18;
  reg                 io_in_r_bypass_regNext_14_1_stall_18;
  reg        [15:0]   io_in_r_bypass_regNext_14_2_data_18;
  reg                 io_in_r_bypass_regNext_14_2_load_store_18;
  reg                 io_in_r_bypass_regNext_14_2_df_is_ws_18;
  reg                 io_in_r_bypass_regNext_14_2_stall_18;
  reg        [15:0]   io_in_r_bypass_regNext_14_3_data_18;
  reg                 io_in_r_bypass_regNext_14_3_load_store_18;
  reg                 io_in_r_bypass_regNext_14_3_df_is_ws_18;
  reg                 io_in_r_bypass_regNext_14_3_stall_18;
  reg        [15:0]   io_in_r_bypass_regNext_15_0_data_18;
  reg                 io_in_r_bypass_regNext_15_0_load_store_18;
  reg                 io_in_r_bypass_regNext_15_0_df_is_ws_18;
  reg                 io_in_r_bypass_regNext_15_0_stall_18;
  reg        [15:0]   io_in_r_bypass_regNext_15_1_data_18;
  reg                 io_in_r_bypass_regNext_15_1_load_store_18;
  reg                 io_in_r_bypass_regNext_15_1_df_is_ws_18;
  reg                 io_in_r_bypass_regNext_15_1_stall_18;
  reg        [15:0]   io_in_r_bypass_regNext_15_2_data_18;
  reg                 io_in_r_bypass_regNext_15_2_load_store_18;
  reg                 io_in_r_bypass_regNext_15_2_df_is_ws_18;
  reg                 io_in_r_bypass_regNext_15_2_stall_18;
  reg        [15:0]   io_in_r_bypass_regNext_15_3_data_18;
  reg                 io_in_r_bypass_regNext_15_3_load_store_18;
  reg                 io_in_r_bypass_regNext_15_3_df_is_ws_18;
  reg                 io_in_r_bypass_regNext_15_3_stall_18;
  reg        [15:0]   io_in_r_bypass_regNext_16_0_data_18;
  reg                 io_in_r_bypass_regNext_16_0_load_store_18;
  reg                 io_in_r_bypass_regNext_16_0_df_is_ws_18;
  reg                 io_in_r_bypass_regNext_16_0_stall_18;
  reg        [15:0]   io_in_r_bypass_regNext_16_1_data_18;
  reg                 io_in_r_bypass_regNext_16_1_load_store_18;
  reg                 io_in_r_bypass_regNext_16_1_df_is_ws_18;
  reg                 io_in_r_bypass_regNext_16_1_stall_18;
  reg        [15:0]   io_in_r_bypass_regNext_16_2_data_18;
  reg                 io_in_r_bypass_regNext_16_2_load_store_18;
  reg                 io_in_r_bypass_regNext_16_2_df_is_ws_18;
  reg                 io_in_r_bypass_regNext_16_2_stall_18;
  reg        [15:0]   io_in_r_bypass_regNext_16_3_data_18;
  reg                 io_in_r_bypass_regNext_16_3_load_store_18;
  reg                 io_in_r_bypass_regNext_16_3_df_is_ws_18;
  reg                 io_in_r_bypass_regNext_16_3_stall_18;
  reg        [15:0]   io_in_r_bypass_regNext_17_0_data_18;
  reg                 io_in_r_bypass_regNext_17_0_load_store_18;
  reg                 io_in_r_bypass_regNext_17_0_df_is_ws_18;
  reg                 io_in_r_bypass_regNext_17_0_stall_18;
  reg        [15:0]   io_in_r_bypass_regNext_17_1_data_18;
  reg                 io_in_r_bypass_regNext_17_1_load_store_18;
  reg                 io_in_r_bypass_regNext_17_1_df_is_ws_18;
  reg                 io_in_r_bypass_regNext_17_1_stall_18;
  reg        [15:0]   io_in_r_bypass_regNext_17_2_data_18;
  reg                 io_in_r_bypass_regNext_17_2_load_store_18;
  reg                 io_in_r_bypass_regNext_17_2_df_is_ws_18;
  reg                 io_in_r_bypass_regNext_17_2_stall_18;
  reg        [15:0]   io_in_r_bypass_regNext_17_3_data_18;
  reg                 io_in_r_bypass_regNext_17_3_load_store_18;
  reg                 io_in_r_bypass_regNext_17_3_df_is_ws_18;
  reg                 io_in_r_bypass_regNext_17_3_stall_18;
  reg        [15:0]   io_in_r_bypass_regNext_18_0_data_18;
  reg                 io_in_r_bypass_regNext_18_0_load_store_18;
  reg                 io_in_r_bypass_regNext_18_0_df_is_ws_18;
  reg                 io_in_r_bypass_regNext_18_0_stall_18;
  reg        [15:0]   io_in_r_bypass_regNext_18_1_data_18;
  reg                 io_in_r_bypass_regNext_18_1_load_store_18;
  reg                 io_in_r_bypass_regNext_18_1_df_is_ws_18;
  reg                 io_in_r_bypass_regNext_18_1_stall_18;
  reg        [15:0]   io_in_r_bypass_regNext_18_2_data_18;
  reg                 io_in_r_bypass_regNext_18_2_load_store_18;
  reg                 io_in_r_bypass_regNext_18_2_df_is_ws_18;
  reg                 io_in_r_bypass_regNext_18_2_stall_18;
  reg        [15:0]   io_in_r_bypass_regNext_18_3_data_18;
  reg                 io_in_r_bypass_regNext_18_3_load_store_18;
  reg                 io_in_r_bypass_regNext_18_3_df_is_ws_18;
  reg                 io_in_r_bypass_regNext_18_3_stall_18;
  reg        [15:0]   io_in_r_bypass_regNext_19_0_data_18;
  reg                 io_in_r_bypass_regNext_19_0_load_store_18;
  reg                 io_in_r_bypass_regNext_19_0_df_is_ws_18;
  reg                 io_in_r_bypass_regNext_19_0_stall_18;
  reg        [15:0]   io_in_r_bypass_regNext_19_1_data_18;
  reg                 io_in_r_bypass_regNext_19_1_load_store_18;
  reg                 io_in_r_bypass_regNext_19_1_df_is_ws_18;
  reg                 io_in_r_bypass_regNext_19_1_stall_18;
  reg        [15:0]   io_in_r_bypass_regNext_19_2_data_18;
  reg                 io_in_r_bypass_regNext_19_2_load_store_18;
  reg                 io_in_r_bypass_regNext_19_2_df_is_ws_18;
  reg                 io_in_r_bypass_regNext_19_2_stall_18;
  reg        [15:0]   io_in_r_bypass_regNext_19_3_data_18;
  reg                 io_in_r_bypass_regNext_19_3_load_store_18;
  reg                 io_in_r_bypass_regNext_19_3_df_is_ws_18;
  reg                 io_in_r_bypass_regNext_19_3_stall_18;
  reg        [15:0]   io_in_r_bypass_regNext_20_0_data_18;
  reg                 io_in_r_bypass_regNext_20_0_load_store_18;
  reg                 io_in_r_bypass_regNext_20_0_df_is_ws_18;
  reg                 io_in_r_bypass_regNext_20_0_stall_18;
  reg        [15:0]   io_in_r_bypass_regNext_20_1_data_18;
  reg                 io_in_r_bypass_regNext_20_1_load_store_18;
  reg                 io_in_r_bypass_regNext_20_1_df_is_ws_18;
  reg                 io_in_r_bypass_regNext_20_1_stall_18;
  reg        [15:0]   io_in_r_bypass_regNext_20_2_data_18;
  reg                 io_in_r_bypass_regNext_20_2_load_store_18;
  reg                 io_in_r_bypass_regNext_20_2_df_is_ws_18;
  reg                 io_in_r_bypass_regNext_20_2_stall_18;
  reg        [15:0]   io_in_r_bypass_regNext_20_3_data_18;
  reg                 io_in_r_bypass_regNext_20_3_load_store_18;
  reg                 io_in_r_bypass_regNext_20_3_df_is_ws_18;
  reg                 io_in_r_bypass_regNext_20_3_stall_18;
  reg        [15:0]   io_in_r_bypass_regNext_21_0_data_18;
  reg                 io_in_r_bypass_regNext_21_0_load_store_18;
  reg                 io_in_r_bypass_regNext_21_0_df_is_ws_18;
  reg                 io_in_r_bypass_regNext_21_0_stall_18;
  reg        [15:0]   io_in_r_bypass_regNext_21_1_data_18;
  reg                 io_in_r_bypass_regNext_21_1_load_store_18;
  reg                 io_in_r_bypass_regNext_21_1_df_is_ws_18;
  reg                 io_in_r_bypass_regNext_21_1_stall_18;
  reg        [15:0]   io_in_r_bypass_regNext_21_2_data_18;
  reg                 io_in_r_bypass_regNext_21_2_load_store_18;
  reg                 io_in_r_bypass_regNext_21_2_df_is_ws_18;
  reg                 io_in_r_bypass_regNext_21_2_stall_18;
  reg        [15:0]   io_in_r_bypass_regNext_21_3_data_18;
  reg                 io_in_r_bypass_regNext_21_3_load_store_18;
  reg                 io_in_r_bypass_regNext_21_3_df_is_ws_18;
  reg                 io_in_r_bypass_regNext_21_3_stall_18;
  reg        [15:0]   io_in_r_bypass_regNext_22_0_data_18;
  reg                 io_in_r_bypass_regNext_22_0_load_store_18;
  reg                 io_in_r_bypass_regNext_22_0_df_is_ws_18;
  reg                 io_in_r_bypass_regNext_22_0_stall_18;
  reg        [15:0]   io_in_r_bypass_regNext_22_1_data_18;
  reg                 io_in_r_bypass_regNext_22_1_load_store_18;
  reg                 io_in_r_bypass_regNext_22_1_df_is_ws_18;
  reg                 io_in_r_bypass_regNext_22_1_stall_18;
  reg        [15:0]   io_in_r_bypass_regNext_22_2_data_18;
  reg                 io_in_r_bypass_regNext_22_2_load_store_18;
  reg                 io_in_r_bypass_regNext_22_2_df_is_ws_18;
  reg                 io_in_r_bypass_regNext_22_2_stall_18;
  reg        [15:0]   io_in_r_bypass_regNext_22_3_data_18;
  reg                 io_in_r_bypass_regNext_22_3_load_store_18;
  reg                 io_in_r_bypass_regNext_22_3_df_is_ws_18;
  reg                 io_in_r_bypass_regNext_22_3_stall_18;
  reg        [15:0]   io_in_r_bypass_regNext_23_0_data_18;
  reg                 io_in_r_bypass_regNext_23_0_load_store_18;
  reg                 io_in_r_bypass_regNext_23_0_df_is_ws_18;
  reg                 io_in_r_bypass_regNext_23_0_stall_18;
  reg        [15:0]   io_in_r_bypass_regNext_23_1_data_18;
  reg                 io_in_r_bypass_regNext_23_1_load_store_18;
  reg                 io_in_r_bypass_regNext_23_1_df_is_ws_18;
  reg                 io_in_r_bypass_regNext_23_1_stall_18;
  reg        [15:0]   io_in_r_bypass_regNext_23_2_data_18;
  reg                 io_in_r_bypass_regNext_23_2_load_store_18;
  reg                 io_in_r_bypass_regNext_23_2_df_is_ws_18;
  reg                 io_in_r_bypass_regNext_23_2_stall_18;
  reg        [15:0]   io_in_r_bypass_regNext_23_3_data_18;
  reg                 io_in_r_bypass_regNext_23_3_load_store_18;
  reg                 io_in_r_bypass_regNext_23_3_df_is_ws_18;
  reg                 io_in_r_bypass_regNext_23_3_stall_18;
  reg        [15:0]   io_in_r_bypass_regNext_24_0_data_18;
  reg                 io_in_r_bypass_regNext_24_0_load_store_18;
  reg                 io_in_r_bypass_regNext_24_0_df_is_ws_18;
  reg                 io_in_r_bypass_regNext_24_0_stall_18;
  reg        [15:0]   io_in_r_bypass_regNext_24_1_data_18;
  reg                 io_in_r_bypass_regNext_24_1_load_store_18;
  reg                 io_in_r_bypass_regNext_24_1_df_is_ws_18;
  reg                 io_in_r_bypass_regNext_24_1_stall_18;
  reg        [15:0]   io_in_r_bypass_regNext_24_2_data_18;
  reg                 io_in_r_bypass_regNext_24_2_load_store_18;
  reg                 io_in_r_bypass_regNext_24_2_df_is_ws_18;
  reg                 io_in_r_bypass_regNext_24_2_stall_18;
  reg        [15:0]   io_in_r_bypass_regNext_24_3_data_18;
  reg                 io_in_r_bypass_regNext_24_3_load_store_18;
  reg                 io_in_r_bypass_regNext_24_3_df_is_ws_18;
  reg                 io_in_r_bypass_regNext_24_3_stall_18;
  reg        [15:0]   io_in_r_bypass_regNext_25_0_data_18;
  reg                 io_in_r_bypass_regNext_25_0_load_store_18;
  reg                 io_in_r_bypass_regNext_25_0_df_is_ws_18;
  reg                 io_in_r_bypass_regNext_25_0_stall_18;
  reg        [15:0]   io_in_r_bypass_regNext_25_1_data_18;
  reg                 io_in_r_bypass_regNext_25_1_load_store_18;
  reg                 io_in_r_bypass_regNext_25_1_df_is_ws_18;
  reg                 io_in_r_bypass_regNext_25_1_stall_18;
  reg        [15:0]   io_in_r_bypass_regNext_25_2_data_18;
  reg                 io_in_r_bypass_regNext_25_2_load_store_18;
  reg                 io_in_r_bypass_regNext_25_2_df_is_ws_18;
  reg                 io_in_r_bypass_regNext_25_2_stall_18;
  reg        [15:0]   io_in_r_bypass_regNext_25_3_data_18;
  reg                 io_in_r_bypass_regNext_25_3_load_store_18;
  reg                 io_in_r_bypass_regNext_25_3_df_is_ws_18;
  reg                 io_in_r_bypass_regNext_25_3_stall_18;
  reg        [15:0]   io_in_r_bypass_regNext_26_0_data_18;
  reg                 io_in_r_bypass_regNext_26_0_load_store_18;
  reg                 io_in_r_bypass_regNext_26_0_df_is_ws_18;
  reg                 io_in_r_bypass_regNext_26_0_stall_18;
  reg        [15:0]   io_in_r_bypass_regNext_26_1_data_18;
  reg                 io_in_r_bypass_regNext_26_1_load_store_18;
  reg                 io_in_r_bypass_regNext_26_1_df_is_ws_18;
  reg                 io_in_r_bypass_regNext_26_1_stall_18;
  reg        [15:0]   io_in_r_bypass_regNext_26_2_data_18;
  reg                 io_in_r_bypass_regNext_26_2_load_store_18;
  reg                 io_in_r_bypass_regNext_26_2_df_is_ws_18;
  reg                 io_in_r_bypass_regNext_26_2_stall_18;
  reg        [15:0]   io_in_r_bypass_regNext_26_3_data_18;
  reg                 io_in_r_bypass_regNext_26_3_load_store_18;
  reg                 io_in_r_bypass_regNext_26_3_df_is_ws_18;
  reg                 io_in_r_bypass_regNext_26_3_stall_18;
  reg        [15:0]   io_in_r_bypass_regNext_27_0_data_18;
  reg                 io_in_r_bypass_regNext_27_0_load_store_18;
  reg                 io_in_r_bypass_regNext_27_0_df_is_ws_18;
  reg                 io_in_r_bypass_regNext_27_0_stall_18;
  reg        [15:0]   io_in_r_bypass_regNext_27_1_data_18;
  reg                 io_in_r_bypass_regNext_27_1_load_store_18;
  reg                 io_in_r_bypass_regNext_27_1_df_is_ws_18;
  reg                 io_in_r_bypass_regNext_27_1_stall_18;
  reg        [15:0]   io_in_r_bypass_regNext_27_2_data_18;
  reg                 io_in_r_bypass_regNext_27_2_load_store_18;
  reg                 io_in_r_bypass_regNext_27_2_df_is_ws_18;
  reg                 io_in_r_bypass_regNext_27_2_stall_18;
  reg        [15:0]   io_in_r_bypass_regNext_27_3_data_18;
  reg                 io_in_r_bypass_regNext_27_3_load_store_18;
  reg                 io_in_r_bypass_regNext_27_3_df_is_ws_18;
  reg                 io_in_r_bypass_regNext_27_3_stall_18;
  reg        [15:0]   io_in_r_bypass_regNext_28_0_data_18;
  reg                 io_in_r_bypass_regNext_28_0_load_store_18;
  reg                 io_in_r_bypass_regNext_28_0_df_is_ws_18;
  reg                 io_in_r_bypass_regNext_28_0_stall_18;
  reg        [15:0]   io_in_r_bypass_regNext_28_1_data_18;
  reg                 io_in_r_bypass_regNext_28_1_load_store_18;
  reg                 io_in_r_bypass_regNext_28_1_df_is_ws_18;
  reg                 io_in_r_bypass_regNext_28_1_stall_18;
  reg        [15:0]   io_in_r_bypass_regNext_28_2_data_18;
  reg                 io_in_r_bypass_regNext_28_2_load_store_18;
  reg                 io_in_r_bypass_regNext_28_2_df_is_ws_18;
  reg                 io_in_r_bypass_regNext_28_2_stall_18;
  reg        [15:0]   io_in_r_bypass_regNext_28_3_data_18;
  reg                 io_in_r_bypass_regNext_28_3_load_store_18;
  reg                 io_in_r_bypass_regNext_28_3_df_is_ws_18;
  reg                 io_in_r_bypass_regNext_28_3_stall_18;
  reg        [15:0]   io_in_r_bypass_regNext_29_0_data_18;
  reg                 io_in_r_bypass_regNext_29_0_load_store_18;
  reg                 io_in_r_bypass_regNext_29_0_df_is_ws_18;
  reg                 io_in_r_bypass_regNext_29_0_stall_18;
  reg        [15:0]   io_in_r_bypass_regNext_29_1_data_18;
  reg                 io_in_r_bypass_regNext_29_1_load_store_18;
  reg                 io_in_r_bypass_regNext_29_1_df_is_ws_18;
  reg                 io_in_r_bypass_regNext_29_1_stall_18;
  reg        [15:0]   io_in_r_bypass_regNext_29_2_data_18;
  reg                 io_in_r_bypass_regNext_29_2_load_store_18;
  reg                 io_in_r_bypass_regNext_29_2_df_is_ws_18;
  reg                 io_in_r_bypass_regNext_29_2_stall_18;
  reg        [15:0]   io_in_r_bypass_regNext_29_3_data_18;
  reg                 io_in_r_bypass_regNext_29_3_load_store_18;
  reg                 io_in_r_bypass_regNext_29_3_df_is_ws_18;
  reg                 io_in_r_bypass_regNext_29_3_stall_18;
  reg        [15:0]   io_in_r_bypass_regNext_30_0_data_18;
  reg                 io_in_r_bypass_regNext_30_0_load_store_18;
  reg                 io_in_r_bypass_regNext_30_0_df_is_ws_18;
  reg                 io_in_r_bypass_regNext_30_0_stall_18;
  reg        [15:0]   io_in_r_bypass_regNext_30_1_data_18;
  reg                 io_in_r_bypass_regNext_30_1_load_store_18;
  reg                 io_in_r_bypass_regNext_30_1_df_is_ws_18;
  reg                 io_in_r_bypass_regNext_30_1_stall_18;
  reg        [15:0]   io_in_r_bypass_regNext_30_2_data_18;
  reg                 io_in_r_bypass_regNext_30_2_load_store_18;
  reg                 io_in_r_bypass_regNext_30_2_df_is_ws_18;
  reg                 io_in_r_bypass_regNext_30_2_stall_18;
  reg        [15:0]   io_in_r_bypass_regNext_30_3_data_18;
  reg                 io_in_r_bypass_regNext_30_3_load_store_18;
  reg                 io_in_r_bypass_regNext_30_3_df_is_ws_18;
  reg                 io_in_r_bypass_regNext_30_3_stall_18;
  reg        [15:0]   io_in_r_bypass_regNext_31_0_data_18;
  reg                 io_in_r_bypass_regNext_31_0_load_store_18;
  reg                 io_in_r_bypass_regNext_31_0_df_is_ws_18;
  reg                 io_in_r_bypass_regNext_31_0_stall_18;
  reg        [15:0]   io_in_r_bypass_regNext_31_1_data_18;
  reg                 io_in_r_bypass_regNext_31_1_load_store_18;
  reg                 io_in_r_bypass_regNext_31_1_df_is_ws_18;
  reg                 io_in_r_bypass_regNext_31_1_stall_18;
  reg        [15:0]   io_in_r_bypass_regNext_31_2_data_18;
  reg                 io_in_r_bypass_regNext_31_2_load_store_18;
  reg                 io_in_r_bypass_regNext_31_2_df_is_ws_18;
  reg                 io_in_r_bypass_regNext_31_2_stall_18;
  reg        [15:0]   io_in_r_bypass_regNext_31_3_data_18;
  reg                 io_in_r_bypass_regNext_31_3_load_store_18;
  reg                 io_in_r_bypass_regNext_31_3_df_is_ws_18;
  reg                 io_in_r_bypass_regNext_31_3_stall_18;
  reg        [15:0]   io_in_r_bypass_regNext_0_0_data_19;
  reg                 io_in_r_bypass_regNext_0_0_load_store_19;
  reg                 io_in_r_bypass_regNext_0_0_df_is_ws_19;
  reg                 io_in_r_bypass_regNext_0_0_stall_19;
  reg        [15:0]   io_in_r_bypass_regNext_0_1_data_19;
  reg                 io_in_r_bypass_regNext_0_1_load_store_19;
  reg                 io_in_r_bypass_regNext_0_1_df_is_ws_19;
  reg                 io_in_r_bypass_regNext_0_1_stall_19;
  reg        [15:0]   io_in_r_bypass_regNext_0_2_data_19;
  reg                 io_in_r_bypass_regNext_0_2_load_store_19;
  reg                 io_in_r_bypass_regNext_0_2_df_is_ws_19;
  reg                 io_in_r_bypass_regNext_0_2_stall_19;
  reg        [15:0]   io_in_r_bypass_regNext_0_3_data_19;
  reg                 io_in_r_bypass_regNext_0_3_load_store_19;
  reg                 io_in_r_bypass_regNext_0_3_df_is_ws_19;
  reg                 io_in_r_bypass_regNext_0_3_stall_19;
  reg        [15:0]   io_in_r_bypass_regNext_1_0_data_19;
  reg                 io_in_r_bypass_regNext_1_0_load_store_19;
  reg                 io_in_r_bypass_regNext_1_0_df_is_ws_19;
  reg                 io_in_r_bypass_regNext_1_0_stall_19;
  reg        [15:0]   io_in_r_bypass_regNext_1_1_data_19;
  reg                 io_in_r_bypass_regNext_1_1_load_store_19;
  reg                 io_in_r_bypass_regNext_1_1_df_is_ws_19;
  reg                 io_in_r_bypass_regNext_1_1_stall_19;
  reg        [15:0]   io_in_r_bypass_regNext_1_2_data_19;
  reg                 io_in_r_bypass_regNext_1_2_load_store_19;
  reg                 io_in_r_bypass_regNext_1_2_df_is_ws_19;
  reg                 io_in_r_bypass_regNext_1_2_stall_19;
  reg        [15:0]   io_in_r_bypass_regNext_1_3_data_19;
  reg                 io_in_r_bypass_regNext_1_3_load_store_19;
  reg                 io_in_r_bypass_regNext_1_3_df_is_ws_19;
  reg                 io_in_r_bypass_regNext_1_3_stall_19;
  reg        [15:0]   io_in_r_bypass_regNext_2_0_data_19;
  reg                 io_in_r_bypass_regNext_2_0_load_store_19;
  reg                 io_in_r_bypass_regNext_2_0_df_is_ws_19;
  reg                 io_in_r_bypass_regNext_2_0_stall_19;
  reg        [15:0]   io_in_r_bypass_regNext_2_1_data_19;
  reg                 io_in_r_bypass_regNext_2_1_load_store_19;
  reg                 io_in_r_bypass_regNext_2_1_df_is_ws_19;
  reg                 io_in_r_bypass_regNext_2_1_stall_19;
  reg        [15:0]   io_in_r_bypass_regNext_2_2_data_19;
  reg                 io_in_r_bypass_regNext_2_2_load_store_19;
  reg                 io_in_r_bypass_regNext_2_2_df_is_ws_19;
  reg                 io_in_r_bypass_regNext_2_2_stall_19;
  reg        [15:0]   io_in_r_bypass_regNext_2_3_data_19;
  reg                 io_in_r_bypass_regNext_2_3_load_store_19;
  reg                 io_in_r_bypass_regNext_2_3_df_is_ws_19;
  reg                 io_in_r_bypass_regNext_2_3_stall_19;
  reg        [15:0]   io_in_r_bypass_regNext_3_0_data_19;
  reg                 io_in_r_bypass_regNext_3_0_load_store_19;
  reg                 io_in_r_bypass_regNext_3_0_df_is_ws_19;
  reg                 io_in_r_bypass_regNext_3_0_stall_19;
  reg        [15:0]   io_in_r_bypass_regNext_3_1_data_19;
  reg                 io_in_r_bypass_regNext_3_1_load_store_19;
  reg                 io_in_r_bypass_regNext_3_1_df_is_ws_19;
  reg                 io_in_r_bypass_regNext_3_1_stall_19;
  reg        [15:0]   io_in_r_bypass_regNext_3_2_data_19;
  reg                 io_in_r_bypass_regNext_3_2_load_store_19;
  reg                 io_in_r_bypass_regNext_3_2_df_is_ws_19;
  reg                 io_in_r_bypass_regNext_3_2_stall_19;
  reg        [15:0]   io_in_r_bypass_regNext_3_3_data_19;
  reg                 io_in_r_bypass_regNext_3_3_load_store_19;
  reg                 io_in_r_bypass_regNext_3_3_df_is_ws_19;
  reg                 io_in_r_bypass_regNext_3_3_stall_19;
  reg        [15:0]   io_in_r_bypass_regNext_4_0_data_19;
  reg                 io_in_r_bypass_regNext_4_0_load_store_19;
  reg                 io_in_r_bypass_regNext_4_0_df_is_ws_19;
  reg                 io_in_r_bypass_regNext_4_0_stall_19;
  reg        [15:0]   io_in_r_bypass_regNext_4_1_data_19;
  reg                 io_in_r_bypass_regNext_4_1_load_store_19;
  reg                 io_in_r_bypass_regNext_4_1_df_is_ws_19;
  reg                 io_in_r_bypass_regNext_4_1_stall_19;
  reg        [15:0]   io_in_r_bypass_regNext_4_2_data_19;
  reg                 io_in_r_bypass_regNext_4_2_load_store_19;
  reg                 io_in_r_bypass_regNext_4_2_df_is_ws_19;
  reg                 io_in_r_bypass_regNext_4_2_stall_19;
  reg        [15:0]   io_in_r_bypass_regNext_4_3_data_19;
  reg                 io_in_r_bypass_regNext_4_3_load_store_19;
  reg                 io_in_r_bypass_regNext_4_3_df_is_ws_19;
  reg                 io_in_r_bypass_regNext_4_3_stall_19;
  reg        [15:0]   io_in_r_bypass_regNext_5_0_data_19;
  reg                 io_in_r_bypass_regNext_5_0_load_store_19;
  reg                 io_in_r_bypass_regNext_5_0_df_is_ws_19;
  reg                 io_in_r_bypass_regNext_5_0_stall_19;
  reg        [15:0]   io_in_r_bypass_regNext_5_1_data_19;
  reg                 io_in_r_bypass_regNext_5_1_load_store_19;
  reg                 io_in_r_bypass_regNext_5_1_df_is_ws_19;
  reg                 io_in_r_bypass_regNext_5_1_stall_19;
  reg        [15:0]   io_in_r_bypass_regNext_5_2_data_19;
  reg                 io_in_r_bypass_regNext_5_2_load_store_19;
  reg                 io_in_r_bypass_regNext_5_2_df_is_ws_19;
  reg                 io_in_r_bypass_regNext_5_2_stall_19;
  reg        [15:0]   io_in_r_bypass_regNext_5_3_data_19;
  reg                 io_in_r_bypass_regNext_5_3_load_store_19;
  reg                 io_in_r_bypass_regNext_5_3_df_is_ws_19;
  reg                 io_in_r_bypass_regNext_5_3_stall_19;
  reg        [15:0]   io_in_r_bypass_regNext_6_0_data_19;
  reg                 io_in_r_bypass_regNext_6_0_load_store_19;
  reg                 io_in_r_bypass_regNext_6_0_df_is_ws_19;
  reg                 io_in_r_bypass_regNext_6_0_stall_19;
  reg        [15:0]   io_in_r_bypass_regNext_6_1_data_19;
  reg                 io_in_r_bypass_regNext_6_1_load_store_19;
  reg                 io_in_r_bypass_regNext_6_1_df_is_ws_19;
  reg                 io_in_r_bypass_regNext_6_1_stall_19;
  reg        [15:0]   io_in_r_bypass_regNext_6_2_data_19;
  reg                 io_in_r_bypass_regNext_6_2_load_store_19;
  reg                 io_in_r_bypass_regNext_6_2_df_is_ws_19;
  reg                 io_in_r_bypass_regNext_6_2_stall_19;
  reg        [15:0]   io_in_r_bypass_regNext_6_3_data_19;
  reg                 io_in_r_bypass_regNext_6_3_load_store_19;
  reg                 io_in_r_bypass_regNext_6_3_df_is_ws_19;
  reg                 io_in_r_bypass_regNext_6_3_stall_19;
  reg        [15:0]   io_in_r_bypass_regNext_7_0_data_19;
  reg                 io_in_r_bypass_regNext_7_0_load_store_19;
  reg                 io_in_r_bypass_regNext_7_0_df_is_ws_19;
  reg                 io_in_r_bypass_regNext_7_0_stall_19;
  reg        [15:0]   io_in_r_bypass_regNext_7_1_data_19;
  reg                 io_in_r_bypass_regNext_7_1_load_store_19;
  reg                 io_in_r_bypass_regNext_7_1_df_is_ws_19;
  reg                 io_in_r_bypass_regNext_7_1_stall_19;
  reg        [15:0]   io_in_r_bypass_regNext_7_2_data_19;
  reg                 io_in_r_bypass_regNext_7_2_load_store_19;
  reg                 io_in_r_bypass_regNext_7_2_df_is_ws_19;
  reg                 io_in_r_bypass_regNext_7_2_stall_19;
  reg        [15:0]   io_in_r_bypass_regNext_7_3_data_19;
  reg                 io_in_r_bypass_regNext_7_3_load_store_19;
  reg                 io_in_r_bypass_regNext_7_3_df_is_ws_19;
  reg                 io_in_r_bypass_regNext_7_3_stall_19;
  reg        [15:0]   io_in_r_bypass_regNext_8_0_data_19;
  reg                 io_in_r_bypass_regNext_8_0_load_store_19;
  reg                 io_in_r_bypass_regNext_8_0_df_is_ws_19;
  reg                 io_in_r_bypass_regNext_8_0_stall_19;
  reg        [15:0]   io_in_r_bypass_regNext_8_1_data_19;
  reg                 io_in_r_bypass_regNext_8_1_load_store_19;
  reg                 io_in_r_bypass_regNext_8_1_df_is_ws_19;
  reg                 io_in_r_bypass_regNext_8_1_stall_19;
  reg        [15:0]   io_in_r_bypass_regNext_8_2_data_19;
  reg                 io_in_r_bypass_regNext_8_2_load_store_19;
  reg                 io_in_r_bypass_regNext_8_2_df_is_ws_19;
  reg                 io_in_r_bypass_regNext_8_2_stall_19;
  reg        [15:0]   io_in_r_bypass_regNext_8_3_data_19;
  reg                 io_in_r_bypass_regNext_8_3_load_store_19;
  reg                 io_in_r_bypass_regNext_8_3_df_is_ws_19;
  reg                 io_in_r_bypass_regNext_8_3_stall_19;
  reg        [15:0]   io_in_r_bypass_regNext_9_0_data_19;
  reg                 io_in_r_bypass_regNext_9_0_load_store_19;
  reg                 io_in_r_bypass_regNext_9_0_df_is_ws_19;
  reg                 io_in_r_bypass_regNext_9_0_stall_19;
  reg        [15:0]   io_in_r_bypass_regNext_9_1_data_19;
  reg                 io_in_r_bypass_regNext_9_1_load_store_19;
  reg                 io_in_r_bypass_regNext_9_1_df_is_ws_19;
  reg                 io_in_r_bypass_regNext_9_1_stall_19;
  reg        [15:0]   io_in_r_bypass_regNext_9_2_data_19;
  reg                 io_in_r_bypass_regNext_9_2_load_store_19;
  reg                 io_in_r_bypass_regNext_9_2_df_is_ws_19;
  reg                 io_in_r_bypass_regNext_9_2_stall_19;
  reg        [15:0]   io_in_r_bypass_regNext_9_3_data_19;
  reg                 io_in_r_bypass_regNext_9_3_load_store_19;
  reg                 io_in_r_bypass_regNext_9_3_df_is_ws_19;
  reg                 io_in_r_bypass_regNext_9_3_stall_19;
  reg        [15:0]   io_in_r_bypass_regNext_10_0_data_19;
  reg                 io_in_r_bypass_regNext_10_0_load_store_19;
  reg                 io_in_r_bypass_regNext_10_0_df_is_ws_19;
  reg                 io_in_r_bypass_regNext_10_0_stall_19;
  reg        [15:0]   io_in_r_bypass_regNext_10_1_data_19;
  reg                 io_in_r_bypass_regNext_10_1_load_store_19;
  reg                 io_in_r_bypass_regNext_10_1_df_is_ws_19;
  reg                 io_in_r_bypass_regNext_10_1_stall_19;
  reg        [15:0]   io_in_r_bypass_regNext_10_2_data_19;
  reg                 io_in_r_bypass_regNext_10_2_load_store_19;
  reg                 io_in_r_bypass_regNext_10_2_df_is_ws_19;
  reg                 io_in_r_bypass_regNext_10_2_stall_19;
  reg        [15:0]   io_in_r_bypass_regNext_10_3_data_19;
  reg                 io_in_r_bypass_regNext_10_3_load_store_19;
  reg                 io_in_r_bypass_regNext_10_3_df_is_ws_19;
  reg                 io_in_r_bypass_regNext_10_3_stall_19;
  reg        [15:0]   io_in_r_bypass_regNext_11_0_data_19;
  reg                 io_in_r_bypass_regNext_11_0_load_store_19;
  reg                 io_in_r_bypass_regNext_11_0_df_is_ws_19;
  reg                 io_in_r_bypass_regNext_11_0_stall_19;
  reg        [15:0]   io_in_r_bypass_regNext_11_1_data_19;
  reg                 io_in_r_bypass_regNext_11_1_load_store_19;
  reg                 io_in_r_bypass_regNext_11_1_df_is_ws_19;
  reg                 io_in_r_bypass_regNext_11_1_stall_19;
  reg        [15:0]   io_in_r_bypass_regNext_11_2_data_19;
  reg                 io_in_r_bypass_regNext_11_2_load_store_19;
  reg                 io_in_r_bypass_regNext_11_2_df_is_ws_19;
  reg                 io_in_r_bypass_regNext_11_2_stall_19;
  reg        [15:0]   io_in_r_bypass_regNext_11_3_data_19;
  reg                 io_in_r_bypass_regNext_11_3_load_store_19;
  reg                 io_in_r_bypass_regNext_11_3_df_is_ws_19;
  reg                 io_in_r_bypass_regNext_11_3_stall_19;
  reg        [15:0]   io_in_r_bypass_regNext_12_0_data_19;
  reg                 io_in_r_bypass_regNext_12_0_load_store_19;
  reg                 io_in_r_bypass_regNext_12_0_df_is_ws_19;
  reg                 io_in_r_bypass_regNext_12_0_stall_19;
  reg        [15:0]   io_in_r_bypass_regNext_12_1_data_19;
  reg                 io_in_r_bypass_regNext_12_1_load_store_19;
  reg                 io_in_r_bypass_regNext_12_1_df_is_ws_19;
  reg                 io_in_r_bypass_regNext_12_1_stall_19;
  reg        [15:0]   io_in_r_bypass_regNext_12_2_data_19;
  reg                 io_in_r_bypass_regNext_12_2_load_store_19;
  reg                 io_in_r_bypass_regNext_12_2_df_is_ws_19;
  reg                 io_in_r_bypass_regNext_12_2_stall_19;
  reg        [15:0]   io_in_r_bypass_regNext_12_3_data_19;
  reg                 io_in_r_bypass_regNext_12_3_load_store_19;
  reg                 io_in_r_bypass_regNext_12_3_df_is_ws_19;
  reg                 io_in_r_bypass_regNext_12_3_stall_19;
  reg        [15:0]   io_in_r_bypass_regNext_13_0_data_19;
  reg                 io_in_r_bypass_regNext_13_0_load_store_19;
  reg                 io_in_r_bypass_regNext_13_0_df_is_ws_19;
  reg                 io_in_r_bypass_regNext_13_0_stall_19;
  reg        [15:0]   io_in_r_bypass_regNext_13_1_data_19;
  reg                 io_in_r_bypass_regNext_13_1_load_store_19;
  reg                 io_in_r_bypass_regNext_13_1_df_is_ws_19;
  reg                 io_in_r_bypass_regNext_13_1_stall_19;
  reg        [15:0]   io_in_r_bypass_regNext_13_2_data_19;
  reg                 io_in_r_bypass_regNext_13_2_load_store_19;
  reg                 io_in_r_bypass_regNext_13_2_df_is_ws_19;
  reg                 io_in_r_bypass_regNext_13_2_stall_19;
  reg        [15:0]   io_in_r_bypass_regNext_13_3_data_19;
  reg                 io_in_r_bypass_regNext_13_3_load_store_19;
  reg                 io_in_r_bypass_regNext_13_3_df_is_ws_19;
  reg                 io_in_r_bypass_regNext_13_3_stall_19;
  reg        [15:0]   io_in_r_bypass_regNext_14_0_data_19;
  reg                 io_in_r_bypass_regNext_14_0_load_store_19;
  reg                 io_in_r_bypass_regNext_14_0_df_is_ws_19;
  reg                 io_in_r_bypass_regNext_14_0_stall_19;
  reg        [15:0]   io_in_r_bypass_regNext_14_1_data_19;
  reg                 io_in_r_bypass_regNext_14_1_load_store_19;
  reg                 io_in_r_bypass_regNext_14_1_df_is_ws_19;
  reg                 io_in_r_bypass_regNext_14_1_stall_19;
  reg        [15:0]   io_in_r_bypass_regNext_14_2_data_19;
  reg                 io_in_r_bypass_regNext_14_2_load_store_19;
  reg                 io_in_r_bypass_regNext_14_2_df_is_ws_19;
  reg                 io_in_r_bypass_regNext_14_2_stall_19;
  reg        [15:0]   io_in_r_bypass_regNext_14_3_data_19;
  reg                 io_in_r_bypass_regNext_14_3_load_store_19;
  reg                 io_in_r_bypass_regNext_14_3_df_is_ws_19;
  reg                 io_in_r_bypass_regNext_14_3_stall_19;
  reg        [15:0]   io_in_r_bypass_regNext_15_0_data_19;
  reg                 io_in_r_bypass_regNext_15_0_load_store_19;
  reg                 io_in_r_bypass_regNext_15_0_df_is_ws_19;
  reg                 io_in_r_bypass_regNext_15_0_stall_19;
  reg        [15:0]   io_in_r_bypass_regNext_15_1_data_19;
  reg                 io_in_r_bypass_regNext_15_1_load_store_19;
  reg                 io_in_r_bypass_regNext_15_1_df_is_ws_19;
  reg                 io_in_r_bypass_regNext_15_1_stall_19;
  reg        [15:0]   io_in_r_bypass_regNext_15_2_data_19;
  reg                 io_in_r_bypass_regNext_15_2_load_store_19;
  reg                 io_in_r_bypass_regNext_15_2_df_is_ws_19;
  reg                 io_in_r_bypass_regNext_15_2_stall_19;
  reg        [15:0]   io_in_r_bypass_regNext_15_3_data_19;
  reg                 io_in_r_bypass_regNext_15_3_load_store_19;
  reg                 io_in_r_bypass_regNext_15_3_df_is_ws_19;
  reg                 io_in_r_bypass_regNext_15_3_stall_19;
  reg        [15:0]   io_in_r_bypass_regNext_16_0_data_19;
  reg                 io_in_r_bypass_regNext_16_0_load_store_19;
  reg                 io_in_r_bypass_regNext_16_0_df_is_ws_19;
  reg                 io_in_r_bypass_regNext_16_0_stall_19;
  reg        [15:0]   io_in_r_bypass_regNext_16_1_data_19;
  reg                 io_in_r_bypass_regNext_16_1_load_store_19;
  reg                 io_in_r_bypass_regNext_16_1_df_is_ws_19;
  reg                 io_in_r_bypass_regNext_16_1_stall_19;
  reg        [15:0]   io_in_r_bypass_regNext_16_2_data_19;
  reg                 io_in_r_bypass_regNext_16_2_load_store_19;
  reg                 io_in_r_bypass_regNext_16_2_df_is_ws_19;
  reg                 io_in_r_bypass_regNext_16_2_stall_19;
  reg        [15:0]   io_in_r_bypass_regNext_16_3_data_19;
  reg                 io_in_r_bypass_regNext_16_3_load_store_19;
  reg                 io_in_r_bypass_regNext_16_3_df_is_ws_19;
  reg                 io_in_r_bypass_regNext_16_3_stall_19;
  reg        [15:0]   io_in_r_bypass_regNext_17_0_data_19;
  reg                 io_in_r_bypass_regNext_17_0_load_store_19;
  reg                 io_in_r_bypass_regNext_17_0_df_is_ws_19;
  reg                 io_in_r_bypass_regNext_17_0_stall_19;
  reg        [15:0]   io_in_r_bypass_regNext_17_1_data_19;
  reg                 io_in_r_bypass_regNext_17_1_load_store_19;
  reg                 io_in_r_bypass_regNext_17_1_df_is_ws_19;
  reg                 io_in_r_bypass_regNext_17_1_stall_19;
  reg        [15:0]   io_in_r_bypass_regNext_17_2_data_19;
  reg                 io_in_r_bypass_regNext_17_2_load_store_19;
  reg                 io_in_r_bypass_regNext_17_2_df_is_ws_19;
  reg                 io_in_r_bypass_regNext_17_2_stall_19;
  reg        [15:0]   io_in_r_bypass_regNext_17_3_data_19;
  reg                 io_in_r_bypass_regNext_17_3_load_store_19;
  reg                 io_in_r_bypass_regNext_17_3_df_is_ws_19;
  reg                 io_in_r_bypass_regNext_17_3_stall_19;
  reg        [15:0]   io_in_r_bypass_regNext_18_0_data_19;
  reg                 io_in_r_bypass_regNext_18_0_load_store_19;
  reg                 io_in_r_bypass_regNext_18_0_df_is_ws_19;
  reg                 io_in_r_bypass_regNext_18_0_stall_19;
  reg        [15:0]   io_in_r_bypass_regNext_18_1_data_19;
  reg                 io_in_r_bypass_regNext_18_1_load_store_19;
  reg                 io_in_r_bypass_regNext_18_1_df_is_ws_19;
  reg                 io_in_r_bypass_regNext_18_1_stall_19;
  reg        [15:0]   io_in_r_bypass_regNext_18_2_data_19;
  reg                 io_in_r_bypass_regNext_18_2_load_store_19;
  reg                 io_in_r_bypass_regNext_18_2_df_is_ws_19;
  reg                 io_in_r_bypass_regNext_18_2_stall_19;
  reg        [15:0]   io_in_r_bypass_regNext_18_3_data_19;
  reg                 io_in_r_bypass_regNext_18_3_load_store_19;
  reg                 io_in_r_bypass_regNext_18_3_df_is_ws_19;
  reg                 io_in_r_bypass_regNext_18_3_stall_19;
  reg        [15:0]   io_in_r_bypass_regNext_19_0_data_19;
  reg                 io_in_r_bypass_regNext_19_0_load_store_19;
  reg                 io_in_r_bypass_regNext_19_0_df_is_ws_19;
  reg                 io_in_r_bypass_regNext_19_0_stall_19;
  reg        [15:0]   io_in_r_bypass_regNext_19_1_data_19;
  reg                 io_in_r_bypass_regNext_19_1_load_store_19;
  reg                 io_in_r_bypass_regNext_19_1_df_is_ws_19;
  reg                 io_in_r_bypass_regNext_19_1_stall_19;
  reg        [15:0]   io_in_r_bypass_regNext_19_2_data_19;
  reg                 io_in_r_bypass_regNext_19_2_load_store_19;
  reg                 io_in_r_bypass_regNext_19_2_df_is_ws_19;
  reg                 io_in_r_bypass_regNext_19_2_stall_19;
  reg        [15:0]   io_in_r_bypass_regNext_19_3_data_19;
  reg                 io_in_r_bypass_regNext_19_3_load_store_19;
  reg                 io_in_r_bypass_regNext_19_3_df_is_ws_19;
  reg                 io_in_r_bypass_regNext_19_3_stall_19;
  reg        [15:0]   io_in_r_bypass_regNext_20_0_data_19;
  reg                 io_in_r_bypass_regNext_20_0_load_store_19;
  reg                 io_in_r_bypass_regNext_20_0_df_is_ws_19;
  reg                 io_in_r_bypass_regNext_20_0_stall_19;
  reg        [15:0]   io_in_r_bypass_regNext_20_1_data_19;
  reg                 io_in_r_bypass_regNext_20_1_load_store_19;
  reg                 io_in_r_bypass_regNext_20_1_df_is_ws_19;
  reg                 io_in_r_bypass_regNext_20_1_stall_19;
  reg        [15:0]   io_in_r_bypass_regNext_20_2_data_19;
  reg                 io_in_r_bypass_regNext_20_2_load_store_19;
  reg                 io_in_r_bypass_regNext_20_2_df_is_ws_19;
  reg                 io_in_r_bypass_regNext_20_2_stall_19;
  reg        [15:0]   io_in_r_bypass_regNext_20_3_data_19;
  reg                 io_in_r_bypass_regNext_20_3_load_store_19;
  reg                 io_in_r_bypass_regNext_20_3_df_is_ws_19;
  reg                 io_in_r_bypass_regNext_20_3_stall_19;
  reg        [15:0]   io_in_r_bypass_regNext_21_0_data_19;
  reg                 io_in_r_bypass_regNext_21_0_load_store_19;
  reg                 io_in_r_bypass_regNext_21_0_df_is_ws_19;
  reg                 io_in_r_bypass_regNext_21_0_stall_19;
  reg        [15:0]   io_in_r_bypass_regNext_21_1_data_19;
  reg                 io_in_r_bypass_regNext_21_1_load_store_19;
  reg                 io_in_r_bypass_regNext_21_1_df_is_ws_19;
  reg                 io_in_r_bypass_regNext_21_1_stall_19;
  reg        [15:0]   io_in_r_bypass_regNext_21_2_data_19;
  reg                 io_in_r_bypass_regNext_21_2_load_store_19;
  reg                 io_in_r_bypass_regNext_21_2_df_is_ws_19;
  reg                 io_in_r_bypass_regNext_21_2_stall_19;
  reg        [15:0]   io_in_r_bypass_regNext_21_3_data_19;
  reg                 io_in_r_bypass_regNext_21_3_load_store_19;
  reg                 io_in_r_bypass_regNext_21_3_df_is_ws_19;
  reg                 io_in_r_bypass_regNext_21_3_stall_19;
  reg        [15:0]   io_in_r_bypass_regNext_22_0_data_19;
  reg                 io_in_r_bypass_regNext_22_0_load_store_19;
  reg                 io_in_r_bypass_regNext_22_0_df_is_ws_19;
  reg                 io_in_r_bypass_regNext_22_0_stall_19;
  reg        [15:0]   io_in_r_bypass_regNext_22_1_data_19;
  reg                 io_in_r_bypass_regNext_22_1_load_store_19;
  reg                 io_in_r_bypass_regNext_22_1_df_is_ws_19;
  reg                 io_in_r_bypass_regNext_22_1_stall_19;
  reg        [15:0]   io_in_r_bypass_regNext_22_2_data_19;
  reg                 io_in_r_bypass_regNext_22_2_load_store_19;
  reg                 io_in_r_bypass_regNext_22_2_df_is_ws_19;
  reg                 io_in_r_bypass_regNext_22_2_stall_19;
  reg        [15:0]   io_in_r_bypass_regNext_22_3_data_19;
  reg                 io_in_r_bypass_regNext_22_3_load_store_19;
  reg                 io_in_r_bypass_regNext_22_3_df_is_ws_19;
  reg                 io_in_r_bypass_regNext_22_3_stall_19;
  reg        [15:0]   io_in_r_bypass_regNext_23_0_data_19;
  reg                 io_in_r_bypass_regNext_23_0_load_store_19;
  reg                 io_in_r_bypass_regNext_23_0_df_is_ws_19;
  reg                 io_in_r_bypass_regNext_23_0_stall_19;
  reg        [15:0]   io_in_r_bypass_regNext_23_1_data_19;
  reg                 io_in_r_bypass_regNext_23_1_load_store_19;
  reg                 io_in_r_bypass_regNext_23_1_df_is_ws_19;
  reg                 io_in_r_bypass_regNext_23_1_stall_19;
  reg        [15:0]   io_in_r_bypass_regNext_23_2_data_19;
  reg                 io_in_r_bypass_regNext_23_2_load_store_19;
  reg                 io_in_r_bypass_regNext_23_2_df_is_ws_19;
  reg                 io_in_r_bypass_regNext_23_2_stall_19;
  reg        [15:0]   io_in_r_bypass_regNext_23_3_data_19;
  reg                 io_in_r_bypass_regNext_23_3_load_store_19;
  reg                 io_in_r_bypass_regNext_23_3_df_is_ws_19;
  reg                 io_in_r_bypass_regNext_23_3_stall_19;
  reg        [15:0]   io_in_r_bypass_regNext_24_0_data_19;
  reg                 io_in_r_bypass_regNext_24_0_load_store_19;
  reg                 io_in_r_bypass_regNext_24_0_df_is_ws_19;
  reg                 io_in_r_bypass_regNext_24_0_stall_19;
  reg        [15:0]   io_in_r_bypass_regNext_24_1_data_19;
  reg                 io_in_r_bypass_regNext_24_1_load_store_19;
  reg                 io_in_r_bypass_regNext_24_1_df_is_ws_19;
  reg                 io_in_r_bypass_regNext_24_1_stall_19;
  reg        [15:0]   io_in_r_bypass_regNext_24_2_data_19;
  reg                 io_in_r_bypass_regNext_24_2_load_store_19;
  reg                 io_in_r_bypass_regNext_24_2_df_is_ws_19;
  reg                 io_in_r_bypass_regNext_24_2_stall_19;
  reg        [15:0]   io_in_r_bypass_regNext_24_3_data_19;
  reg                 io_in_r_bypass_regNext_24_3_load_store_19;
  reg                 io_in_r_bypass_regNext_24_3_df_is_ws_19;
  reg                 io_in_r_bypass_regNext_24_3_stall_19;
  reg        [15:0]   io_in_r_bypass_regNext_25_0_data_19;
  reg                 io_in_r_bypass_regNext_25_0_load_store_19;
  reg                 io_in_r_bypass_regNext_25_0_df_is_ws_19;
  reg                 io_in_r_bypass_regNext_25_0_stall_19;
  reg        [15:0]   io_in_r_bypass_regNext_25_1_data_19;
  reg                 io_in_r_bypass_regNext_25_1_load_store_19;
  reg                 io_in_r_bypass_regNext_25_1_df_is_ws_19;
  reg                 io_in_r_bypass_regNext_25_1_stall_19;
  reg        [15:0]   io_in_r_bypass_regNext_25_2_data_19;
  reg                 io_in_r_bypass_regNext_25_2_load_store_19;
  reg                 io_in_r_bypass_regNext_25_2_df_is_ws_19;
  reg                 io_in_r_bypass_regNext_25_2_stall_19;
  reg        [15:0]   io_in_r_bypass_regNext_25_3_data_19;
  reg                 io_in_r_bypass_regNext_25_3_load_store_19;
  reg                 io_in_r_bypass_regNext_25_3_df_is_ws_19;
  reg                 io_in_r_bypass_regNext_25_3_stall_19;
  reg        [15:0]   io_in_r_bypass_regNext_26_0_data_19;
  reg                 io_in_r_bypass_regNext_26_0_load_store_19;
  reg                 io_in_r_bypass_regNext_26_0_df_is_ws_19;
  reg                 io_in_r_bypass_regNext_26_0_stall_19;
  reg        [15:0]   io_in_r_bypass_regNext_26_1_data_19;
  reg                 io_in_r_bypass_regNext_26_1_load_store_19;
  reg                 io_in_r_bypass_regNext_26_1_df_is_ws_19;
  reg                 io_in_r_bypass_regNext_26_1_stall_19;
  reg        [15:0]   io_in_r_bypass_regNext_26_2_data_19;
  reg                 io_in_r_bypass_regNext_26_2_load_store_19;
  reg                 io_in_r_bypass_regNext_26_2_df_is_ws_19;
  reg                 io_in_r_bypass_regNext_26_2_stall_19;
  reg        [15:0]   io_in_r_bypass_regNext_26_3_data_19;
  reg                 io_in_r_bypass_regNext_26_3_load_store_19;
  reg                 io_in_r_bypass_regNext_26_3_df_is_ws_19;
  reg                 io_in_r_bypass_regNext_26_3_stall_19;
  reg        [15:0]   io_in_r_bypass_regNext_27_0_data_19;
  reg                 io_in_r_bypass_regNext_27_0_load_store_19;
  reg                 io_in_r_bypass_regNext_27_0_df_is_ws_19;
  reg                 io_in_r_bypass_regNext_27_0_stall_19;
  reg        [15:0]   io_in_r_bypass_regNext_27_1_data_19;
  reg                 io_in_r_bypass_regNext_27_1_load_store_19;
  reg                 io_in_r_bypass_regNext_27_1_df_is_ws_19;
  reg                 io_in_r_bypass_regNext_27_1_stall_19;
  reg        [15:0]   io_in_r_bypass_regNext_27_2_data_19;
  reg                 io_in_r_bypass_regNext_27_2_load_store_19;
  reg                 io_in_r_bypass_regNext_27_2_df_is_ws_19;
  reg                 io_in_r_bypass_regNext_27_2_stall_19;
  reg        [15:0]   io_in_r_bypass_regNext_27_3_data_19;
  reg                 io_in_r_bypass_regNext_27_3_load_store_19;
  reg                 io_in_r_bypass_regNext_27_3_df_is_ws_19;
  reg                 io_in_r_bypass_regNext_27_3_stall_19;
  reg        [15:0]   io_in_r_bypass_regNext_28_0_data_19;
  reg                 io_in_r_bypass_regNext_28_0_load_store_19;
  reg                 io_in_r_bypass_regNext_28_0_df_is_ws_19;
  reg                 io_in_r_bypass_regNext_28_0_stall_19;
  reg        [15:0]   io_in_r_bypass_regNext_28_1_data_19;
  reg                 io_in_r_bypass_regNext_28_1_load_store_19;
  reg                 io_in_r_bypass_regNext_28_1_df_is_ws_19;
  reg                 io_in_r_bypass_regNext_28_1_stall_19;
  reg        [15:0]   io_in_r_bypass_regNext_28_2_data_19;
  reg                 io_in_r_bypass_regNext_28_2_load_store_19;
  reg                 io_in_r_bypass_regNext_28_2_df_is_ws_19;
  reg                 io_in_r_bypass_regNext_28_2_stall_19;
  reg        [15:0]   io_in_r_bypass_regNext_28_3_data_19;
  reg                 io_in_r_bypass_regNext_28_3_load_store_19;
  reg                 io_in_r_bypass_regNext_28_3_df_is_ws_19;
  reg                 io_in_r_bypass_regNext_28_3_stall_19;
  reg        [15:0]   io_in_r_bypass_regNext_29_0_data_19;
  reg                 io_in_r_bypass_regNext_29_0_load_store_19;
  reg                 io_in_r_bypass_regNext_29_0_df_is_ws_19;
  reg                 io_in_r_bypass_regNext_29_0_stall_19;
  reg        [15:0]   io_in_r_bypass_regNext_29_1_data_19;
  reg                 io_in_r_bypass_regNext_29_1_load_store_19;
  reg                 io_in_r_bypass_regNext_29_1_df_is_ws_19;
  reg                 io_in_r_bypass_regNext_29_1_stall_19;
  reg        [15:0]   io_in_r_bypass_regNext_29_2_data_19;
  reg                 io_in_r_bypass_regNext_29_2_load_store_19;
  reg                 io_in_r_bypass_regNext_29_2_df_is_ws_19;
  reg                 io_in_r_bypass_regNext_29_2_stall_19;
  reg        [15:0]   io_in_r_bypass_regNext_29_3_data_19;
  reg                 io_in_r_bypass_regNext_29_3_load_store_19;
  reg                 io_in_r_bypass_regNext_29_3_df_is_ws_19;
  reg                 io_in_r_bypass_regNext_29_3_stall_19;
  reg        [15:0]   io_in_r_bypass_regNext_30_0_data_19;
  reg                 io_in_r_bypass_regNext_30_0_load_store_19;
  reg                 io_in_r_bypass_regNext_30_0_df_is_ws_19;
  reg                 io_in_r_bypass_regNext_30_0_stall_19;
  reg        [15:0]   io_in_r_bypass_regNext_30_1_data_19;
  reg                 io_in_r_bypass_regNext_30_1_load_store_19;
  reg                 io_in_r_bypass_regNext_30_1_df_is_ws_19;
  reg                 io_in_r_bypass_regNext_30_1_stall_19;
  reg        [15:0]   io_in_r_bypass_regNext_30_2_data_19;
  reg                 io_in_r_bypass_regNext_30_2_load_store_19;
  reg                 io_in_r_bypass_regNext_30_2_df_is_ws_19;
  reg                 io_in_r_bypass_regNext_30_2_stall_19;
  reg        [15:0]   io_in_r_bypass_regNext_30_3_data_19;
  reg                 io_in_r_bypass_regNext_30_3_load_store_19;
  reg                 io_in_r_bypass_regNext_30_3_df_is_ws_19;
  reg                 io_in_r_bypass_regNext_30_3_stall_19;
  reg        [15:0]   io_in_r_bypass_regNext_31_0_data_19;
  reg                 io_in_r_bypass_regNext_31_0_load_store_19;
  reg                 io_in_r_bypass_regNext_31_0_df_is_ws_19;
  reg                 io_in_r_bypass_regNext_31_0_stall_19;
  reg        [15:0]   io_in_r_bypass_regNext_31_1_data_19;
  reg                 io_in_r_bypass_regNext_31_1_load_store_19;
  reg                 io_in_r_bypass_regNext_31_1_df_is_ws_19;
  reg                 io_in_r_bypass_regNext_31_1_stall_19;
  reg        [15:0]   io_in_r_bypass_regNext_31_2_data_19;
  reg                 io_in_r_bypass_regNext_31_2_load_store_19;
  reg                 io_in_r_bypass_regNext_31_2_df_is_ws_19;
  reg                 io_in_r_bypass_regNext_31_2_stall_19;
  reg        [15:0]   io_in_r_bypass_regNext_31_3_data_19;
  reg                 io_in_r_bypass_regNext_31_3_load_store_19;
  reg                 io_in_r_bypass_regNext_31_3_df_is_ws_19;
  reg                 io_in_r_bypass_regNext_31_3_stall_19;
  reg        [15:0]   io_in_r_bypass_regNext_0_0_data_20;
  reg                 io_in_r_bypass_regNext_0_0_load_store_20;
  reg                 io_in_r_bypass_regNext_0_0_df_is_ws_20;
  reg                 io_in_r_bypass_regNext_0_0_stall_20;
  reg        [15:0]   io_in_r_bypass_regNext_0_1_data_20;
  reg                 io_in_r_bypass_regNext_0_1_load_store_20;
  reg                 io_in_r_bypass_regNext_0_1_df_is_ws_20;
  reg                 io_in_r_bypass_regNext_0_1_stall_20;
  reg        [15:0]   io_in_r_bypass_regNext_0_2_data_20;
  reg                 io_in_r_bypass_regNext_0_2_load_store_20;
  reg                 io_in_r_bypass_regNext_0_2_df_is_ws_20;
  reg                 io_in_r_bypass_regNext_0_2_stall_20;
  reg        [15:0]   io_in_r_bypass_regNext_0_3_data_20;
  reg                 io_in_r_bypass_regNext_0_3_load_store_20;
  reg                 io_in_r_bypass_regNext_0_3_df_is_ws_20;
  reg                 io_in_r_bypass_regNext_0_3_stall_20;
  reg        [15:0]   io_in_r_bypass_regNext_1_0_data_20;
  reg                 io_in_r_bypass_regNext_1_0_load_store_20;
  reg                 io_in_r_bypass_regNext_1_0_df_is_ws_20;
  reg                 io_in_r_bypass_regNext_1_0_stall_20;
  reg        [15:0]   io_in_r_bypass_regNext_1_1_data_20;
  reg                 io_in_r_bypass_regNext_1_1_load_store_20;
  reg                 io_in_r_bypass_regNext_1_1_df_is_ws_20;
  reg                 io_in_r_bypass_regNext_1_1_stall_20;
  reg        [15:0]   io_in_r_bypass_regNext_1_2_data_20;
  reg                 io_in_r_bypass_regNext_1_2_load_store_20;
  reg                 io_in_r_bypass_regNext_1_2_df_is_ws_20;
  reg                 io_in_r_bypass_regNext_1_2_stall_20;
  reg        [15:0]   io_in_r_bypass_regNext_1_3_data_20;
  reg                 io_in_r_bypass_regNext_1_3_load_store_20;
  reg                 io_in_r_bypass_regNext_1_3_df_is_ws_20;
  reg                 io_in_r_bypass_regNext_1_3_stall_20;
  reg        [15:0]   io_in_r_bypass_regNext_2_0_data_20;
  reg                 io_in_r_bypass_regNext_2_0_load_store_20;
  reg                 io_in_r_bypass_regNext_2_0_df_is_ws_20;
  reg                 io_in_r_bypass_regNext_2_0_stall_20;
  reg        [15:0]   io_in_r_bypass_regNext_2_1_data_20;
  reg                 io_in_r_bypass_regNext_2_1_load_store_20;
  reg                 io_in_r_bypass_regNext_2_1_df_is_ws_20;
  reg                 io_in_r_bypass_regNext_2_1_stall_20;
  reg        [15:0]   io_in_r_bypass_regNext_2_2_data_20;
  reg                 io_in_r_bypass_regNext_2_2_load_store_20;
  reg                 io_in_r_bypass_regNext_2_2_df_is_ws_20;
  reg                 io_in_r_bypass_regNext_2_2_stall_20;
  reg        [15:0]   io_in_r_bypass_regNext_2_3_data_20;
  reg                 io_in_r_bypass_regNext_2_3_load_store_20;
  reg                 io_in_r_bypass_regNext_2_3_df_is_ws_20;
  reg                 io_in_r_bypass_regNext_2_3_stall_20;
  reg        [15:0]   io_in_r_bypass_regNext_3_0_data_20;
  reg                 io_in_r_bypass_regNext_3_0_load_store_20;
  reg                 io_in_r_bypass_regNext_3_0_df_is_ws_20;
  reg                 io_in_r_bypass_regNext_3_0_stall_20;
  reg        [15:0]   io_in_r_bypass_regNext_3_1_data_20;
  reg                 io_in_r_bypass_regNext_3_1_load_store_20;
  reg                 io_in_r_bypass_regNext_3_1_df_is_ws_20;
  reg                 io_in_r_bypass_regNext_3_1_stall_20;
  reg        [15:0]   io_in_r_bypass_regNext_3_2_data_20;
  reg                 io_in_r_bypass_regNext_3_2_load_store_20;
  reg                 io_in_r_bypass_regNext_3_2_df_is_ws_20;
  reg                 io_in_r_bypass_regNext_3_2_stall_20;
  reg        [15:0]   io_in_r_bypass_regNext_3_3_data_20;
  reg                 io_in_r_bypass_regNext_3_3_load_store_20;
  reg                 io_in_r_bypass_regNext_3_3_df_is_ws_20;
  reg                 io_in_r_bypass_regNext_3_3_stall_20;
  reg        [15:0]   io_in_r_bypass_regNext_4_0_data_20;
  reg                 io_in_r_bypass_regNext_4_0_load_store_20;
  reg                 io_in_r_bypass_regNext_4_0_df_is_ws_20;
  reg                 io_in_r_bypass_regNext_4_0_stall_20;
  reg        [15:0]   io_in_r_bypass_regNext_4_1_data_20;
  reg                 io_in_r_bypass_regNext_4_1_load_store_20;
  reg                 io_in_r_bypass_regNext_4_1_df_is_ws_20;
  reg                 io_in_r_bypass_regNext_4_1_stall_20;
  reg        [15:0]   io_in_r_bypass_regNext_4_2_data_20;
  reg                 io_in_r_bypass_regNext_4_2_load_store_20;
  reg                 io_in_r_bypass_regNext_4_2_df_is_ws_20;
  reg                 io_in_r_bypass_regNext_4_2_stall_20;
  reg        [15:0]   io_in_r_bypass_regNext_4_3_data_20;
  reg                 io_in_r_bypass_regNext_4_3_load_store_20;
  reg                 io_in_r_bypass_regNext_4_3_df_is_ws_20;
  reg                 io_in_r_bypass_regNext_4_3_stall_20;
  reg        [15:0]   io_in_r_bypass_regNext_5_0_data_20;
  reg                 io_in_r_bypass_regNext_5_0_load_store_20;
  reg                 io_in_r_bypass_regNext_5_0_df_is_ws_20;
  reg                 io_in_r_bypass_regNext_5_0_stall_20;
  reg        [15:0]   io_in_r_bypass_regNext_5_1_data_20;
  reg                 io_in_r_bypass_regNext_5_1_load_store_20;
  reg                 io_in_r_bypass_regNext_5_1_df_is_ws_20;
  reg                 io_in_r_bypass_regNext_5_1_stall_20;
  reg        [15:0]   io_in_r_bypass_regNext_5_2_data_20;
  reg                 io_in_r_bypass_regNext_5_2_load_store_20;
  reg                 io_in_r_bypass_regNext_5_2_df_is_ws_20;
  reg                 io_in_r_bypass_regNext_5_2_stall_20;
  reg        [15:0]   io_in_r_bypass_regNext_5_3_data_20;
  reg                 io_in_r_bypass_regNext_5_3_load_store_20;
  reg                 io_in_r_bypass_regNext_5_3_df_is_ws_20;
  reg                 io_in_r_bypass_regNext_5_3_stall_20;
  reg        [15:0]   io_in_r_bypass_regNext_6_0_data_20;
  reg                 io_in_r_bypass_regNext_6_0_load_store_20;
  reg                 io_in_r_bypass_regNext_6_0_df_is_ws_20;
  reg                 io_in_r_bypass_regNext_6_0_stall_20;
  reg        [15:0]   io_in_r_bypass_regNext_6_1_data_20;
  reg                 io_in_r_bypass_regNext_6_1_load_store_20;
  reg                 io_in_r_bypass_regNext_6_1_df_is_ws_20;
  reg                 io_in_r_bypass_regNext_6_1_stall_20;
  reg        [15:0]   io_in_r_bypass_regNext_6_2_data_20;
  reg                 io_in_r_bypass_regNext_6_2_load_store_20;
  reg                 io_in_r_bypass_regNext_6_2_df_is_ws_20;
  reg                 io_in_r_bypass_regNext_6_2_stall_20;
  reg        [15:0]   io_in_r_bypass_regNext_6_3_data_20;
  reg                 io_in_r_bypass_regNext_6_3_load_store_20;
  reg                 io_in_r_bypass_regNext_6_3_df_is_ws_20;
  reg                 io_in_r_bypass_regNext_6_3_stall_20;
  reg        [15:0]   io_in_r_bypass_regNext_7_0_data_20;
  reg                 io_in_r_bypass_regNext_7_0_load_store_20;
  reg                 io_in_r_bypass_regNext_7_0_df_is_ws_20;
  reg                 io_in_r_bypass_regNext_7_0_stall_20;
  reg        [15:0]   io_in_r_bypass_regNext_7_1_data_20;
  reg                 io_in_r_bypass_regNext_7_1_load_store_20;
  reg                 io_in_r_bypass_regNext_7_1_df_is_ws_20;
  reg                 io_in_r_bypass_regNext_7_1_stall_20;
  reg        [15:0]   io_in_r_bypass_regNext_7_2_data_20;
  reg                 io_in_r_bypass_regNext_7_2_load_store_20;
  reg                 io_in_r_bypass_regNext_7_2_df_is_ws_20;
  reg                 io_in_r_bypass_regNext_7_2_stall_20;
  reg        [15:0]   io_in_r_bypass_regNext_7_3_data_20;
  reg                 io_in_r_bypass_regNext_7_3_load_store_20;
  reg                 io_in_r_bypass_regNext_7_3_df_is_ws_20;
  reg                 io_in_r_bypass_regNext_7_3_stall_20;
  reg        [15:0]   io_in_r_bypass_regNext_8_0_data_20;
  reg                 io_in_r_bypass_regNext_8_0_load_store_20;
  reg                 io_in_r_bypass_regNext_8_0_df_is_ws_20;
  reg                 io_in_r_bypass_regNext_8_0_stall_20;
  reg        [15:0]   io_in_r_bypass_regNext_8_1_data_20;
  reg                 io_in_r_bypass_regNext_8_1_load_store_20;
  reg                 io_in_r_bypass_regNext_8_1_df_is_ws_20;
  reg                 io_in_r_bypass_regNext_8_1_stall_20;
  reg        [15:0]   io_in_r_bypass_regNext_8_2_data_20;
  reg                 io_in_r_bypass_regNext_8_2_load_store_20;
  reg                 io_in_r_bypass_regNext_8_2_df_is_ws_20;
  reg                 io_in_r_bypass_regNext_8_2_stall_20;
  reg        [15:0]   io_in_r_bypass_regNext_8_3_data_20;
  reg                 io_in_r_bypass_regNext_8_3_load_store_20;
  reg                 io_in_r_bypass_regNext_8_3_df_is_ws_20;
  reg                 io_in_r_bypass_regNext_8_3_stall_20;
  reg        [15:0]   io_in_r_bypass_regNext_9_0_data_20;
  reg                 io_in_r_bypass_regNext_9_0_load_store_20;
  reg                 io_in_r_bypass_regNext_9_0_df_is_ws_20;
  reg                 io_in_r_bypass_regNext_9_0_stall_20;
  reg        [15:0]   io_in_r_bypass_regNext_9_1_data_20;
  reg                 io_in_r_bypass_regNext_9_1_load_store_20;
  reg                 io_in_r_bypass_regNext_9_1_df_is_ws_20;
  reg                 io_in_r_bypass_regNext_9_1_stall_20;
  reg        [15:0]   io_in_r_bypass_regNext_9_2_data_20;
  reg                 io_in_r_bypass_regNext_9_2_load_store_20;
  reg                 io_in_r_bypass_regNext_9_2_df_is_ws_20;
  reg                 io_in_r_bypass_regNext_9_2_stall_20;
  reg        [15:0]   io_in_r_bypass_regNext_9_3_data_20;
  reg                 io_in_r_bypass_regNext_9_3_load_store_20;
  reg                 io_in_r_bypass_regNext_9_3_df_is_ws_20;
  reg                 io_in_r_bypass_regNext_9_3_stall_20;
  reg        [15:0]   io_in_r_bypass_regNext_10_0_data_20;
  reg                 io_in_r_bypass_regNext_10_0_load_store_20;
  reg                 io_in_r_bypass_regNext_10_0_df_is_ws_20;
  reg                 io_in_r_bypass_regNext_10_0_stall_20;
  reg        [15:0]   io_in_r_bypass_regNext_10_1_data_20;
  reg                 io_in_r_bypass_regNext_10_1_load_store_20;
  reg                 io_in_r_bypass_regNext_10_1_df_is_ws_20;
  reg                 io_in_r_bypass_regNext_10_1_stall_20;
  reg        [15:0]   io_in_r_bypass_regNext_10_2_data_20;
  reg                 io_in_r_bypass_regNext_10_2_load_store_20;
  reg                 io_in_r_bypass_regNext_10_2_df_is_ws_20;
  reg                 io_in_r_bypass_regNext_10_2_stall_20;
  reg        [15:0]   io_in_r_bypass_regNext_10_3_data_20;
  reg                 io_in_r_bypass_regNext_10_3_load_store_20;
  reg                 io_in_r_bypass_regNext_10_3_df_is_ws_20;
  reg                 io_in_r_bypass_regNext_10_3_stall_20;
  reg        [15:0]   io_in_r_bypass_regNext_11_0_data_20;
  reg                 io_in_r_bypass_regNext_11_0_load_store_20;
  reg                 io_in_r_bypass_regNext_11_0_df_is_ws_20;
  reg                 io_in_r_bypass_regNext_11_0_stall_20;
  reg        [15:0]   io_in_r_bypass_regNext_11_1_data_20;
  reg                 io_in_r_bypass_regNext_11_1_load_store_20;
  reg                 io_in_r_bypass_regNext_11_1_df_is_ws_20;
  reg                 io_in_r_bypass_regNext_11_1_stall_20;
  reg        [15:0]   io_in_r_bypass_regNext_11_2_data_20;
  reg                 io_in_r_bypass_regNext_11_2_load_store_20;
  reg                 io_in_r_bypass_regNext_11_2_df_is_ws_20;
  reg                 io_in_r_bypass_regNext_11_2_stall_20;
  reg        [15:0]   io_in_r_bypass_regNext_11_3_data_20;
  reg                 io_in_r_bypass_regNext_11_3_load_store_20;
  reg                 io_in_r_bypass_regNext_11_3_df_is_ws_20;
  reg                 io_in_r_bypass_regNext_11_3_stall_20;
  reg        [15:0]   io_in_r_bypass_regNext_12_0_data_20;
  reg                 io_in_r_bypass_regNext_12_0_load_store_20;
  reg                 io_in_r_bypass_regNext_12_0_df_is_ws_20;
  reg                 io_in_r_bypass_regNext_12_0_stall_20;
  reg        [15:0]   io_in_r_bypass_regNext_12_1_data_20;
  reg                 io_in_r_bypass_regNext_12_1_load_store_20;
  reg                 io_in_r_bypass_regNext_12_1_df_is_ws_20;
  reg                 io_in_r_bypass_regNext_12_1_stall_20;
  reg        [15:0]   io_in_r_bypass_regNext_12_2_data_20;
  reg                 io_in_r_bypass_regNext_12_2_load_store_20;
  reg                 io_in_r_bypass_regNext_12_2_df_is_ws_20;
  reg                 io_in_r_bypass_regNext_12_2_stall_20;
  reg        [15:0]   io_in_r_bypass_regNext_12_3_data_20;
  reg                 io_in_r_bypass_regNext_12_3_load_store_20;
  reg                 io_in_r_bypass_regNext_12_3_df_is_ws_20;
  reg                 io_in_r_bypass_regNext_12_3_stall_20;
  reg        [15:0]   io_in_r_bypass_regNext_13_0_data_20;
  reg                 io_in_r_bypass_regNext_13_0_load_store_20;
  reg                 io_in_r_bypass_regNext_13_0_df_is_ws_20;
  reg                 io_in_r_bypass_regNext_13_0_stall_20;
  reg        [15:0]   io_in_r_bypass_regNext_13_1_data_20;
  reg                 io_in_r_bypass_regNext_13_1_load_store_20;
  reg                 io_in_r_bypass_regNext_13_1_df_is_ws_20;
  reg                 io_in_r_bypass_regNext_13_1_stall_20;
  reg        [15:0]   io_in_r_bypass_regNext_13_2_data_20;
  reg                 io_in_r_bypass_regNext_13_2_load_store_20;
  reg                 io_in_r_bypass_regNext_13_2_df_is_ws_20;
  reg                 io_in_r_bypass_regNext_13_2_stall_20;
  reg        [15:0]   io_in_r_bypass_regNext_13_3_data_20;
  reg                 io_in_r_bypass_regNext_13_3_load_store_20;
  reg                 io_in_r_bypass_regNext_13_3_df_is_ws_20;
  reg                 io_in_r_bypass_regNext_13_3_stall_20;
  reg        [15:0]   io_in_r_bypass_regNext_14_0_data_20;
  reg                 io_in_r_bypass_regNext_14_0_load_store_20;
  reg                 io_in_r_bypass_regNext_14_0_df_is_ws_20;
  reg                 io_in_r_bypass_regNext_14_0_stall_20;
  reg        [15:0]   io_in_r_bypass_regNext_14_1_data_20;
  reg                 io_in_r_bypass_regNext_14_1_load_store_20;
  reg                 io_in_r_bypass_regNext_14_1_df_is_ws_20;
  reg                 io_in_r_bypass_regNext_14_1_stall_20;
  reg        [15:0]   io_in_r_bypass_regNext_14_2_data_20;
  reg                 io_in_r_bypass_regNext_14_2_load_store_20;
  reg                 io_in_r_bypass_regNext_14_2_df_is_ws_20;
  reg                 io_in_r_bypass_regNext_14_2_stall_20;
  reg        [15:0]   io_in_r_bypass_regNext_14_3_data_20;
  reg                 io_in_r_bypass_regNext_14_3_load_store_20;
  reg                 io_in_r_bypass_regNext_14_3_df_is_ws_20;
  reg                 io_in_r_bypass_regNext_14_3_stall_20;
  reg        [15:0]   io_in_r_bypass_regNext_15_0_data_20;
  reg                 io_in_r_bypass_regNext_15_0_load_store_20;
  reg                 io_in_r_bypass_regNext_15_0_df_is_ws_20;
  reg                 io_in_r_bypass_regNext_15_0_stall_20;
  reg        [15:0]   io_in_r_bypass_regNext_15_1_data_20;
  reg                 io_in_r_bypass_regNext_15_1_load_store_20;
  reg                 io_in_r_bypass_regNext_15_1_df_is_ws_20;
  reg                 io_in_r_bypass_regNext_15_1_stall_20;
  reg        [15:0]   io_in_r_bypass_regNext_15_2_data_20;
  reg                 io_in_r_bypass_regNext_15_2_load_store_20;
  reg                 io_in_r_bypass_regNext_15_2_df_is_ws_20;
  reg                 io_in_r_bypass_regNext_15_2_stall_20;
  reg        [15:0]   io_in_r_bypass_regNext_15_3_data_20;
  reg                 io_in_r_bypass_regNext_15_3_load_store_20;
  reg                 io_in_r_bypass_regNext_15_3_df_is_ws_20;
  reg                 io_in_r_bypass_regNext_15_3_stall_20;
  reg        [15:0]   io_in_r_bypass_regNext_16_0_data_20;
  reg                 io_in_r_bypass_regNext_16_0_load_store_20;
  reg                 io_in_r_bypass_regNext_16_0_df_is_ws_20;
  reg                 io_in_r_bypass_regNext_16_0_stall_20;
  reg        [15:0]   io_in_r_bypass_regNext_16_1_data_20;
  reg                 io_in_r_bypass_regNext_16_1_load_store_20;
  reg                 io_in_r_bypass_regNext_16_1_df_is_ws_20;
  reg                 io_in_r_bypass_regNext_16_1_stall_20;
  reg        [15:0]   io_in_r_bypass_regNext_16_2_data_20;
  reg                 io_in_r_bypass_regNext_16_2_load_store_20;
  reg                 io_in_r_bypass_regNext_16_2_df_is_ws_20;
  reg                 io_in_r_bypass_regNext_16_2_stall_20;
  reg        [15:0]   io_in_r_bypass_regNext_16_3_data_20;
  reg                 io_in_r_bypass_regNext_16_3_load_store_20;
  reg                 io_in_r_bypass_regNext_16_3_df_is_ws_20;
  reg                 io_in_r_bypass_regNext_16_3_stall_20;
  reg        [15:0]   io_in_r_bypass_regNext_17_0_data_20;
  reg                 io_in_r_bypass_regNext_17_0_load_store_20;
  reg                 io_in_r_bypass_regNext_17_0_df_is_ws_20;
  reg                 io_in_r_bypass_regNext_17_0_stall_20;
  reg        [15:0]   io_in_r_bypass_regNext_17_1_data_20;
  reg                 io_in_r_bypass_regNext_17_1_load_store_20;
  reg                 io_in_r_bypass_regNext_17_1_df_is_ws_20;
  reg                 io_in_r_bypass_regNext_17_1_stall_20;
  reg        [15:0]   io_in_r_bypass_regNext_17_2_data_20;
  reg                 io_in_r_bypass_regNext_17_2_load_store_20;
  reg                 io_in_r_bypass_regNext_17_2_df_is_ws_20;
  reg                 io_in_r_bypass_regNext_17_2_stall_20;
  reg        [15:0]   io_in_r_bypass_regNext_17_3_data_20;
  reg                 io_in_r_bypass_regNext_17_3_load_store_20;
  reg                 io_in_r_bypass_regNext_17_3_df_is_ws_20;
  reg                 io_in_r_bypass_regNext_17_3_stall_20;
  reg        [15:0]   io_in_r_bypass_regNext_18_0_data_20;
  reg                 io_in_r_bypass_regNext_18_0_load_store_20;
  reg                 io_in_r_bypass_regNext_18_0_df_is_ws_20;
  reg                 io_in_r_bypass_regNext_18_0_stall_20;
  reg        [15:0]   io_in_r_bypass_regNext_18_1_data_20;
  reg                 io_in_r_bypass_regNext_18_1_load_store_20;
  reg                 io_in_r_bypass_regNext_18_1_df_is_ws_20;
  reg                 io_in_r_bypass_regNext_18_1_stall_20;
  reg        [15:0]   io_in_r_bypass_regNext_18_2_data_20;
  reg                 io_in_r_bypass_regNext_18_2_load_store_20;
  reg                 io_in_r_bypass_regNext_18_2_df_is_ws_20;
  reg                 io_in_r_bypass_regNext_18_2_stall_20;
  reg        [15:0]   io_in_r_bypass_regNext_18_3_data_20;
  reg                 io_in_r_bypass_regNext_18_3_load_store_20;
  reg                 io_in_r_bypass_regNext_18_3_df_is_ws_20;
  reg                 io_in_r_bypass_regNext_18_3_stall_20;
  reg        [15:0]   io_in_r_bypass_regNext_19_0_data_20;
  reg                 io_in_r_bypass_regNext_19_0_load_store_20;
  reg                 io_in_r_bypass_regNext_19_0_df_is_ws_20;
  reg                 io_in_r_bypass_regNext_19_0_stall_20;
  reg        [15:0]   io_in_r_bypass_regNext_19_1_data_20;
  reg                 io_in_r_bypass_regNext_19_1_load_store_20;
  reg                 io_in_r_bypass_regNext_19_1_df_is_ws_20;
  reg                 io_in_r_bypass_regNext_19_1_stall_20;
  reg        [15:0]   io_in_r_bypass_regNext_19_2_data_20;
  reg                 io_in_r_bypass_regNext_19_2_load_store_20;
  reg                 io_in_r_bypass_regNext_19_2_df_is_ws_20;
  reg                 io_in_r_bypass_regNext_19_2_stall_20;
  reg        [15:0]   io_in_r_bypass_regNext_19_3_data_20;
  reg                 io_in_r_bypass_regNext_19_3_load_store_20;
  reg                 io_in_r_bypass_regNext_19_3_df_is_ws_20;
  reg                 io_in_r_bypass_regNext_19_3_stall_20;
  reg        [15:0]   io_in_r_bypass_regNext_20_0_data_20;
  reg                 io_in_r_bypass_regNext_20_0_load_store_20;
  reg                 io_in_r_bypass_regNext_20_0_df_is_ws_20;
  reg                 io_in_r_bypass_regNext_20_0_stall_20;
  reg        [15:0]   io_in_r_bypass_regNext_20_1_data_20;
  reg                 io_in_r_bypass_regNext_20_1_load_store_20;
  reg                 io_in_r_bypass_regNext_20_1_df_is_ws_20;
  reg                 io_in_r_bypass_regNext_20_1_stall_20;
  reg        [15:0]   io_in_r_bypass_regNext_20_2_data_20;
  reg                 io_in_r_bypass_regNext_20_2_load_store_20;
  reg                 io_in_r_bypass_regNext_20_2_df_is_ws_20;
  reg                 io_in_r_bypass_regNext_20_2_stall_20;
  reg        [15:0]   io_in_r_bypass_regNext_20_3_data_20;
  reg                 io_in_r_bypass_regNext_20_3_load_store_20;
  reg                 io_in_r_bypass_regNext_20_3_df_is_ws_20;
  reg                 io_in_r_bypass_regNext_20_3_stall_20;
  reg        [15:0]   io_in_r_bypass_regNext_21_0_data_20;
  reg                 io_in_r_bypass_regNext_21_0_load_store_20;
  reg                 io_in_r_bypass_regNext_21_0_df_is_ws_20;
  reg                 io_in_r_bypass_regNext_21_0_stall_20;
  reg        [15:0]   io_in_r_bypass_regNext_21_1_data_20;
  reg                 io_in_r_bypass_regNext_21_1_load_store_20;
  reg                 io_in_r_bypass_regNext_21_1_df_is_ws_20;
  reg                 io_in_r_bypass_regNext_21_1_stall_20;
  reg        [15:0]   io_in_r_bypass_regNext_21_2_data_20;
  reg                 io_in_r_bypass_regNext_21_2_load_store_20;
  reg                 io_in_r_bypass_regNext_21_2_df_is_ws_20;
  reg                 io_in_r_bypass_regNext_21_2_stall_20;
  reg        [15:0]   io_in_r_bypass_regNext_21_3_data_20;
  reg                 io_in_r_bypass_regNext_21_3_load_store_20;
  reg                 io_in_r_bypass_regNext_21_3_df_is_ws_20;
  reg                 io_in_r_bypass_regNext_21_3_stall_20;
  reg        [15:0]   io_in_r_bypass_regNext_22_0_data_20;
  reg                 io_in_r_bypass_regNext_22_0_load_store_20;
  reg                 io_in_r_bypass_regNext_22_0_df_is_ws_20;
  reg                 io_in_r_bypass_regNext_22_0_stall_20;
  reg        [15:0]   io_in_r_bypass_regNext_22_1_data_20;
  reg                 io_in_r_bypass_regNext_22_1_load_store_20;
  reg                 io_in_r_bypass_regNext_22_1_df_is_ws_20;
  reg                 io_in_r_bypass_regNext_22_1_stall_20;
  reg        [15:0]   io_in_r_bypass_regNext_22_2_data_20;
  reg                 io_in_r_bypass_regNext_22_2_load_store_20;
  reg                 io_in_r_bypass_regNext_22_2_df_is_ws_20;
  reg                 io_in_r_bypass_regNext_22_2_stall_20;
  reg        [15:0]   io_in_r_bypass_regNext_22_3_data_20;
  reg                 io_in_r_bypass_regNext_22_3_load_store_20;
  reg                 io_in_r_bypass_regNext_22_3_df_is_ws_20;
  reg                 io_in_r_bypass_regNext_22_3_stall_20;
  reg        [15:0]   io_in_r_bypass_regNext_23_0_data_20;
  reg                 io_in_r_bypass_regNext_23_0_load_store_20;
  reg                 io_in_r_bypass_regNext_23_0_df_is_ws_20;
  reg                 io_in_r_bypass_regNext_23_0_stall_20;
  reg        [15:0]   io_in_r_bypass_regNext_23_1_data_20;
  reg                 io_in_r_bypass_regNext_23_1_load_store_20;
  reg                 io_in_r_bypass_regNext_23_1_df_is_ws_20;
  reg                 io_in_r_bypass_regNext_23_1_stall_20;
  reg        [15:0]   io_in_r_bypass_regNext_23_2_data_20;
  reg                 io_in_r_bypass_regNext_23_2_load_store_20;
  reg                 io_in_r_bypass_regNext_23_2_df_is_ws_20;
  reg                 io_in_r_bypass_regNext_23_2_stall_20;
  reg        [15:0]   io_in_r_bypass_regNext_23_3_data_20;
  reg                 io_in_r_bypass_regNext_23_3_load_store_20;
  reg                 io_in_r_bypass_regNext_23_3_df_is_ws_20;
  reg                 io_in_r_bypass_regNext_23_3_stall_20;
  reg        [15:0]   io_in_r_bypass_regNext_24_0_data_20;
  reg                 io_in_r_bypass_regNext_24_0_load_store_20;
  reg                 io_in_r_bypass_regNext_24_0_df_is_ws_20;
  reg                 io_in_r_bypass_regNext_24_0_stall_20;
  reg        [15:0]   io_in_r_bypass_regNext_24_1_data_20;
  reg                 io_in_r_bypass_regNext_24_1_load_store_20;
  reg                 io_in_r_bypass_regNext_24_1_df_is_ws_20;
  reg                 io_in_r_bypass_regNext_24_1_stall_20;
  reg        [15:0]   io_in_r_bypass_regNext_24_2_data_20;
  reg                 io_in_r_bypass_regNext_24_2_load_store_20;
  reg                 io_in_r_bypass_regNext_24_2_df_is_ws_20;
  reg                 io_in_r_bypass_regNext_24_2_stall_20;
  reg        [15:0]   io_in_r_bypass_regNext_24_3_data_20;
  reg                 io_in_r_bypass_regNext_24_3_load_store_20;
  reg                 io_in_r_bypass_regNext_24_3_df_is_ws_20;
  reg                 io_in_r_bypass_regNext_24_3_stall_20;
  reg        [15:0]   io_in_r_bypass_regNext_25_0_data_20;
  reg                 io_in_r_bypass_regNext_25_0_load_store_20;
  reg                 io_in_r_bypass_regNext_25_0_df_is_ws_20;
  reg                 io_in_r_bypass_regNext_25_0_stall_20;
  reg        [15:0]   io_in_r_bypass_regNext_25_1_data_20;
  reg                 io_in_r_bypass_regNext_25_1_load_store_20;
  reg                 io_in_r_bypass_regNext_25_1_df_is_ws_20;
  reg                 io_in_r_bypass_regNext_25_1_stall_20;
  reg        [15:0]   io_in_r_bypass_regNext_25_2_data_20;
  reg                 io_in_r_bypass_regNext_25_2_load_store_20;
  reg                 io_in_r_bypass_regNext_25_2_df_is_ws_20;
  reg                 io_in_r_bypass_regNext_25_2_stall_20;
  reg        [15:0]   io_in_r_bypass_regNext_25_3_data_20;
  reg                 io_in_r_bypass_regNext_25_3_load_store_20;
  reg                 io_in_r_bypass_regNext_25_3_df_is_ws_20;
  reg                 io_in_r_bypass_regNext_25_3_stall_20;
  reg        [15:0]   io_in_r_bypass_regNext_26_0_data_20;
  reg                 io_in_r_bypass_regNext_26_0_load_store_20;
  reg                 io_in_r_bypass_regNext_26_0_df_is_ws_20;
  reg                 io_in_r_bypass_regNext_26_0_stall_20;
  reg        [15:0]   io_in_r_bypass_regNext_26_1_data_20;
  reg                 io_in_r_bypass_regNext_26_1_load_store_20;
  reg                 io_in_r_bypass_regNext_26_1_df_is_ws_20;
  reg                 io_in_r_bypass_regNext_26_1_stall_20;
  reg        [15:0]   io_in_r_bypass_regNext_26_2_data_20;
  reg                 io_in_r_bypass_regNext_26_2_load_store_20;
  reg                 io_in_r_bypass_regNext_26_2_df_is_ws_20;
  reg                 io_in_r_bypass_regNext_26_2_stall_20;
  reg        [15:0]   io_in_r_bypass_regNext_26_3_data_20;
  reg                 io_in_r_bypass_regNext_26_3_load_store_20;
  reg                 io_in_r_bypass_regNext_26_3_df_is_ws_20;
  reg                 io_in_r_bypass_regNext_26_3_stall_20;
  reg        [15:0]   io_in_r_bypass_regNext_27_0_data_20;
  reg                 io_in_r_bypass_regNext_27_0_load_store_20;
  reg                 io_in_r_bypass_regNext_27_0_df_is_ws_20;
  reg                 io_in_r_bypass_regNext_27_0_stall_20;
  reg        [15:0]   io_in_r_bypass_regNext_27_1_data_20;
  reg                 io_in_r_bypass_regNext_27_1_load_store_20;
  reg                 io_in_r_bypass_regNext_27_1_df_is_ws_20;
  reg                 io_in_r_bypass_regNext_27_1_stall_20;
  reg        [15:0]   io_in_r_bypass_regNext_27_2_data_20;
  reg                 io_in_r_bypass_regNext_27_2_load_store_20;
  reg                 io_in_r_bypass_regNext_27_2_df_is_ws_20;
  reg                 io_in_r_bypass_regNext_27_2_stall_20;
  reg        [15:0]   io_in_r_bypass_regNext_27_3_data_20;
  reg                 io_in_r_bypass_regNext_27_3_load_store_20;
  reg                 io_in_r_bypass_regNext_27_3_df_is_ws_20;
  reg                 io_in_r_bypass_regNext_27_3_stall_20;
  reg        [15:0]   io_in_r_bypass_regNext_28_0_data_20;
  reg                 io_in_r_bypass_regNext_28_0_load_store_20;
  reg                 io_in_r_bypass_regNext_28_0_df_is_ws_20;
  reg                 io_in_r_bypass_regNext_28_0_stall_20;
  reg        [15:0]   io_in_r_bypass_regNext_28_1_data_20;
  reg                 io_in_r_bypass_regNext_28_1_load_store_20;
  reg                 io_in_r_bypass_regNext_28_1_df_is_ws_20;
  reg                 io_in_r_bypass_regNext_28_1_stall_20;
  reg        [15:0]   io_in_r_bypass_regNext_28_2_data_20;
  reg                 io_in_r_bypass_regNext_28_2_load_store_20;
  reg                 io_in_r_bypass_regNext_28_2_df_is_ws_20;
  reg                 io_in_r_bypass_regNext_28_2_stall_20;
  reg        [15:0]   io_in_r_bypass_regNext_28_3_data_20;
  reg                 io_in_r_bypass_regNext_28_3_load_store_20;
  reg                 io_in_r_bypass_regNext_28_3_df_is_ws_20;
  reg                 io_in_r_bypass_regNext_28_3_stall_20;
  reg        [15:0]   io_in_r_bypass_regNext_29_0_data_20;
  reg                 io_in_r_bypass_regNext_29_0_load_store_20;
  reg                 io_in_r_bypass_regNext_29_0_df_is_ws_20;
  reg                 io_in_r_bypass_regNext_29_0_stall_20;
  reg        [15:0]   io_in_r_bypass_regNext_29_1_data_20;
  reg                 io_in_r_bypass_regNext_29_1_load_store_20;
  reg                 io_in_r_bypass_regNext_29_1_df_is_ws_20;
  reg                 io_in_r_bypass_regNext_29_1_stall_20;
  reg        [15:0]   io_in_r_bypass_regNext_29_2_data_20;
  reg                 io_in_r_bypass_regNext_29_2_load_store_20;
  reg                 io_in_r_bypass_regNext_29_2_df_is_ws_20;
  reg                 io_in_r_bypass_regNext_29_2_stall_20;
  reg        [15:0]   io_in_r_bypass_regNext_29_3_data_20;
  reg                 io_in_r_bypass_regNext_29_3_load_store_20;
  reg                 io_in_r_bypass_regNext_29_3_df_is_ws_20;
  reg                 io_in_r_bypass_regNext_29_3_stall_20;
  reg        [15:0]   io_in_r_bypass_regNext_30_0_data_20;
  reg                 io_in_r_bypass_regNext_30_0_load_store_20;
  reg                 io_in_r_bypass_regNext_30_0_df_is_ws_20;
  reg                 io_in_r_bypass_regNext_30_0_stall_20;
  reg        [15:0]   io_in_r_bypass_regNext_30_1_data_20;
  reg                 io_in_r_bypass_regNext_30_1_load_store_20;
  reg                 io_in_r_bypass_regNext_30_1_df_is_ws_20;
  reg                 io_in_r_bypass_regNext_30_1_stall_20;
  reg        [15:0]   io_in_r_bypass_regNext_30_2_data_20;
  reg                 io_in_r_bypass_regNext_30_2_load_store_20;
  reg                 io_in_r_bypass_regNext_30_2_df_is_ws_20;
  reg                 io_in_r_bypass_regNext_30_2_stall_20;
  reg        [15:0]   io_in_r_bypass_regNext_30_3_data_20;
  reg                 io_in_r_bypass_regNext_30_3_load_store_20;
  reg                 io_in_r_bypass_regNext_30_3_df_is_ws_20;
  reg                 io_in_r_bypass_regNext_30_3_stall_20;
  reg        [15:0]   io_in_r_bypass_regNext_31_0_data_20;
  reg                 io_in_r_bypass_regNext_31_0_load_store_20;
  reg                 io_in_r_bypass_regNext_31_0_df_is_ws_20;
  reg                 io_in_r_bypass_regNext_31_0_stall_20;
  reg        [15:0]   io_in_r_bypass_regNext_31_1_data_20;
  reg                 io_in_r_bypass_regNext_31_1_load_store_20;
  reg                 io_in_r_bypass_regNext_31_1_df_is_ws_20;
  reg                 io_in_r_bypass_regNext_31_1_stall_20;
  reg        [15:0]   io_in_r_bypass_regNext_31_2_data_20;
  reg                 io_in_r_bypass_regNext_31_2_load_store_20;
  reg                 io_in_r_bypass_regNext_31_2_df_is_ws_20;
  reg                 io_in_r_bypass_regNext_31_2_stall_20;
  reg        [15:0]   io_in_r_bypass_regNext_31_3_data_20;
  reg                 io_in_r_bypass_regNext_31_3_load_store_20;
  reg                 io_in_r_bypass_regNext_31_3_df_is_ws_20;
  reg                 io_in_r_bypass_regNext_31_3_stall_20;
  reg        [15:0]   io_in_r_bypass_regNext_0_0_data_21;
  reg                 io_in_r_bypass_regNext_0_0_load_store_21;
  reg                 io_in_r_bypass_regNext_0_0_df_is_ws_21;
  reg                 io_in_r_bypass_regNext_0_0_stall_21;
  reg        [15:0]   io_in_r_bypass_regNext_0_1_data_21;
  reg                 io_in_r_bypass_regNext_0_1_load_store_21;
  reg                 io_in_r_bypass_regNext_0_1_df_is_ws_21;
  reg                 io_in_r_bypass_regNext_0_1_stall_21;
  reg        [15:0]   io_in_r_bypass_regNext_0_2_data_21;
  reg                 io_in_r_bypass_regNext_0_2_load_store_21;
  reg                 io_in_r_bypass_regNext_0_2_df_is_ws_21;
  reg                 io_in_r_bypass_regNext_0_2_stall_21;
  reg        [15:0]   io_in_r_bypass_regNext_0_3_data_21;
  reg                 io_in_r_bypass_regNext_0_3_load_store_21;
  reg                 io_in_r_bypass_regNext_0_3_df_is_ws_21;
  reg                 io_in_r_bypass_regNext_0_3_stall_21;
  reg        [15:0]   io_in_r_bypass_regNext_1_0_data_21;
  reg                 io_in_r_bypass_regNext_1_0_load_store_21;
  reg                 io_in_r_bypass_regNext_1_0_df_is_ws_21;
  reg                 io_in_r_bypass_regNext_1_0_stall_21;
  reg        [15:0]   io_in_r_bypass_regNext_1_1_data_21;
  reg                 io_in_r_bypass_regNext_1_1_load_store_21;
  reg                 io_in_r_bypass_regNext_1_1_df_is_ws_21;
  reg                 io_in_r_bypass_regNext_1_1_stall_21;
  reg        [15:0]   io_in_r_bypass_regNext_1_2_data_21;
  reg                 io_in_r_bypass_regNext_1_2_load_store_21;
  reg                 io_in_r_bypass_regNext_1_2_df_is_ws_21;
  reg                 io_in_r_bypass_regNext_1_2_stall_21;
  reg        [15:0]   io_in_r_bypass_regNext_1_3_data_21;
  reg                 io_in_r_bypass_regNext_1_3_load_store_21;
  reg                 io_in_r_bypass_regNext_1_3_df_is_ws_21;
  reg                 io_in_r_bypass_regNext_1_3_stall_21;
  reg        [15:0]   io_in_r_bypass_regNext_2_0_data_21;
  reg                 io_in_r_bypass_regNext_2_0_load_store_21;
  reg                 io_in_r_bypass_regNext_2_0_df_is_ws_21;
  reg                 io_in_r_bypass_regNext_2_0_stall_21;
  reg        [15:0]   io_in_r_bypass_regNext_2_1_data_21;
  reg                 io_in_r_bypass_regNext_2_1_load_store_21;
  reg                 io_in_r_bypass_regNext_2_1_df_is_ws_21;
  reg                 io_in_r_bypass_regNext_2_1_stall_21;
  reg        [15:0]   io_in_r_bypass_regNext_2_2_data_21;
  reg                 io_in_r_bypass_regNext_2_2_load_store_21;
  reg                 io_in_r_bypass_regNext_2_2_df_is_ws_21;
  reg                 io_in_r_bypass_regNext_2_2_stall_21;
  reg        [15:0]   io_in_r_bypass_regNext_2_3_data_21;
  reg                 io_in_r_bypass_regNext_2_3_load_store_21;
  reg                 io_in_r_bypass_regNext_2_3_df_is_ws_21;
  reg                 io_in_r_bypass_regNext_2_3_stall_21;
  reg        [15:0]   io_in_r_bypass_regNext_3_0_data_21;
  reg                 io_in_r_bypass_regNext_3_0_load_store_21;
  reg                 io_in_r_bypass_regNext_3_0_df_is_ws_21;
  reg                 io_in_r_bypass_regNext_3_0_stall_21;
  reg        [15:0]   io_in_r_bypass_regNext_3_1_data_21;
  reg                 io_in_r_bypass_regNext_3_1_load_store_21;
  reg                 io_in_r_bypass_regNext_3_1_df_is_ws_21;
  reg                 io_in_r_bypass_regNext_3_1_stall_21;
  reg        [15:0]   io_in_r_bypass_regNext_3_2_data_21;
  reg                 io_in_r_bypass_regNext_3_2_load_store_21;
  reg                 io_in_r_bypass_regNext_3_2_df_is_ws_21;
  reg                 io_in_r_bypass_regNext_3_2_stall_21;
  reg        [15:0]   io_in_r_bypass_regNext_3_3_data_21;
  reg                 io_in_r_bypass_regNext_3_3_load_store_21;
  reg                 io_in_r_bypass_regNext_3_3_df_is_ws_21;
  reg                 io_in_r_bypass_regNext_3_3_stall_21;
  reg        [15:0]   io_in_r_bypass_regNext_4_0_data_21;
  reg                 io_in_r_bypass_regNext_4_0_load_store_21;
  reg                 io_in_r_bypass_regNext_4_0_df_is_ws_21;
  reg                 io_in_r_bypass_regNext_4_0_stall_21;
  reg        [15:0]   io_in_r_bypass_regNext_4_1_data_21;
  reg                 io_in_r_bypass_regNext_4_1_load_store_21;
  reg                 io_in_r_bypass_regNext_4_1_df_is_ws_21;
  reg                 io_in_r_bypass_regNext_4_1_stall_21;
  reg        [15:0]   io_in_r_bypass_regNext_4_2_data_21;
  reg                 io_in_r_bypass_regNext_4_2_load_store_21;
  reg                 io_in_r_bypass_regNext_4_2_df_is_ws_21;
  reg                 io_in_r_bypass_regNext_4_2_stall_21;
  reg        [15:0]   io_in_r_bypass_regNext_4_3_data_21;
  reg                 io_in_r_bypass_regNext_4_3_load_store_21;
  reg                 io_in_r_bypass_regNext_4_3_df_is_ws_21;
  reg                 io_in_r_bypass_regNext_4_3_stall_21;
  reg        [15:0]   io_in_r_bypass_regNext_5_0_data_21;
  reg                 io_in_r_bypass_regNext_5_0_load_store_21;
  reg                 io_in_r_bypass_regNext_5_0_df_is_ws_21;
  reg                 io_in_r_bypass_regNext_5_0_stall_21;
  reg        [15:0]   io_in_r_bypass_regNext_5_1_data_21;
  reg                 io_in_r_bypass_regNext_5_1_load_store_21;
  reg                 io_in_r_bypass_regNext_5_1_df_is_ws_21;
  reg                 io_in_r_bypass_regNext_5_1_stall_21;
  reg        [15:0]   io_in_r_bypass_regNext_5_2_data_21;
  reg                 io_in_r_bypass_regNext_5_2_load_store_21;
  reg                 io_in_r_bypass_regNext_5_2_df_is_ws_21;
  reg                 io_in_r_bypass_regNext_5_2_stall_21;
  reg        [15:0]   io_in_r_bypass_regNext_5_3_data_21;
  reg                 io_in_r_bypass_regNext_5_3_load_store_21;
  reg                 io_in_r_bypass_regNext_5_3_df_is_ws_21;
  reg                 io_in_r_bypass_regNext_5_3_stall_21;
  reg        [15:0]   io_in_r_bypass_regNext_6_0_data_21;
  reg                 io_in_r_bypass_regNext_6_0_load_store_21;
  reg                 io_in_r_bypass_regNext_6_0_df_is_ws_21;
  reg                 io_in_r_bypass_regNext_6_0_stall_21;
  reg        [15:0]   io_in_r_bypass_regNext_6_1_data_21;
  reg                 io_in_r_bypass_regNext_6_1_load_store_21;
  reg                 io_in_r_bypass_regNext_6_1_df_is_ws_21;
  reg                 io_in_r_bypass_regNext_6_1_stall_21;
  reg        [15:0]   io_in_r_bypass_regNext_6_2_data_21;
  reg                 io_in_r_bypass_regNext_6_2_load_store_21;
  reg                 io_in_r_bypass_regNext_6_2_df_is_ws_21;
  reg                 io_in_r_bypass_regNext_6_2_stall_21;
  reg        [15:0]   io_in_r_bypass_regNext_6_3_data_21;
  reg                 io_in_r_bypass_regNext_6_3_load_store_21;
  reg                 io_in_r_bypass_regNext_6_3_df_is_ws_21;
  reg                 io_in_r_bypass_regNext_6_3_stall_21;
  reg        [15:0]   io_in_r_bypass_regNext_7_0_data_21;
  reg                 io_in_r_bypass_regNext_7_0_load_store_21;
  reg                 io_in_r_bypass_regNext_7_0_df_is_ws_21;
  reg                 io_in_r_bypass_regNext_7_0_stall_21;
  reg        [15:0]   io_in_r_bypass_regNext_7_1_data_21;
  reg                 io_in_r_bypass_regNext_7_1_load_store_21;
  reg                 io_in_r_bypass_regNext_7_1_df_is_ws_21;
  reg                 io_in_r_bypass_regNext_7_1_stall_21;
  reg        [15:0]   io_in_r_bypass_regNext_7_2_data_21;
  reg                 io_in_r_bypass_regNext_7_2_load_store_21;
  reg                 io_in_r_bypass_regNext_7_2_df_is_ws_21;
  reg                 io_in_r_bypass_regNext_7_2_stall_21;
  reg        [15:0]   io_in_r_bypass_regNext_7_3_data_21;
  reg                 io_in_r_bypass_regNext_7_3_load_store_21;
  reg                 io_in_r_bypass_regNext_7_3_df_is_ws_21;
  reg                 io_in_r_bypass_regNext_7_3_stall_21;
  reg        [15:0]   io_in_r_bypass_regNext_8_0_data_21;
  reg                 io_in_r_bypass_regNext_8_0_load_store_21;
  reg                 io_in_r_bypass_regNext_8_0_df_is_ws_21;
  reg                 io_in_r_bypass_regNext_8_0_stall_21;
  reg        [15:0]   io_in_r_bypass_regNext_8_1_data_21;
  reg                 io_in_r_bypass_regNext_8_1_load_store_21;
  reg                 io_in_r_bypass_regNext_8_1_df_is_ws_21;
  reg                 io_in_r_bypass_regNext_8_1_stall_21;
  reg        [15:0]   io_in_r_bypass_regNext_8_2_data_21;
  reg                 io_in_r_bypass_regNext_8_2_load_store_21;
  reg                 io_in_r_bypass_regNext_8_2_df_is_ws_21;
  reg                 io_in_r_bypass_regNext_8_2_stall_21;
  reg        [15:0]   io_in_r_bypass_regNext_8_3_data_21;
  reg                 io_in_r_bypass_regNext_8_3_load_store_21;
  reg                 io_in_r_bypass_regNext_8_3_df_is_ws_21;
  reg                 io_in_r_bypass_regNext_8_3_stall_21;
  reg        [15:0]   io_in_r_bypass_regNext_9_0_data_21;
  reg                 io_in_r_bypass_regNext_9_0_load_store_21;
  reg                 io_in_r_bypass_regNext_9_0_df_is_ws_21;
  reg                 io_in_r_bypass_regNext_9_0_stall_21;
  reg        [15:0]   io_in_r_bypass_regNext_9_1_data_21;
  reg                 io_in_r_bypass_regNext_9_1_load_store_21;
  reg                 io_in_r_bypass_regNext_9_1_df_is_ws_21;
  reg                 io_in_r_bypass_regNext_9_1_stall_21;
  reg        [15:0]   io_in_r_bypass_regNext_9_2_data_21;
  reg                 io_in_r_bypass_regNext_9_2_load_store_21;
  reg                 io_in_r_bypass_regNext_9_2_df_is_ws_21;
  reg                 io_in_r_bypass_regNext_9_2_stall_21;
  reg        [15:0]   io_in_r_bypass_regNext_9_3_data_21;
  reg                 io_in_r_bypass_regNext_9_3_load_store_21;
  reg                 io_in_r_bypass_regNext_9_3_df_is_ws_21;
  reg                 io_in_r_bypass_regNext_9_3_stall_21;
  reg        [15:0]   io_in_r_bypass_regNext_10_0_data_21;
  reg                 io_in_r_bypass_regNext_10_0_load_store_21;
  reg                 io_in_r_bypass_regNext_10_0_df_is_ws_21;
  reg                 io_in_r_bypass_regNext_10_0_stall_21;
  reg        [15:0]   io_in_r_bypass_regNext_10_1_data_21;
  reg                 io_in_r_bypass_regNext_10_1_load_store_21;
  reg                 io_in_r_bypass_regNext_10_1_df_is_ws_21;
  reg                 io_in_r_bypass_regNext_10_1_stall_21;
  reg        [15:0]   io_in_r_bypass_regNext_10_2_data_21;
  reg                 io_in_r_bypass_regNext_10_2_load_store_21;
  reg                 io_in_r_bypass_regNext_10_2_df_is_ws_21;
  reg                 io_in_r_bypass_regNext_10_2_stall_21;
  reg        [15:0]   io_in_r_bypass_regNext_10_3_data_21;
  reg                 io_in_r_bypass_regNext_10_3_load_store_21;
  reg                 io_in_r_bypass_regNext_10_3_df_is_ws_21;
  reg                 io_in_r_bypass_regNext_10_3_stall_21;
  reg        [15:0]   io_in_r_bypass_regNext_11_0_data_21;
  reg                 io_in_r_bypass_regNext_11_0_load_store_21;
  reg                 io_in_r_bypass_regNext_11_0_df_is_ws_21;
  reg                 io_in_r_bypass_regNext_11_0_stall_21;
  reg        [15:0]   io_in_r_bypass_regNext_11_1_data_21;
  reg                 io_in_r_bypass_regNext_11_1_load_store_21;
  reg                 io_in_r_bypass_regNext_11_1_df_is_ws_21;
  reg                 io_in_r_bypass_regNext_11_1_stall_21;
  reg        [15:0]   io_in_r_bypass_regNext_11_2_data_21;
  reg                 io_in_r_bypass_regNext_11_2_load_store_21;
  reg                 io_in_r_bypass_regNext_11_2_df_is_ws_21;
  reg                 io_in_r_bypass_regNext_11_2_stall_21;
  reg        [15:0]   io_in_r_bypass_regNext_11_3_data_21;
  reg                 io_in_r_bypass_regNext_11_3_load_store_21;
  reg                 io_in_r_bypass_regNext_11_3_df_is_ws_21;
  reg                 io_in_r_bypass_regNext_11_3_stall_21;
  reg        [15:0]   io_in_r_bypass_regNext_12_0_data_21;
  reg                 io_in_r_bypass_regNext_12_0_load_store_21;
  reg                 io_in_r_bypass_regNext_12_0_df_is_ws_21;
  reg                 io_in_r_bypass_regNext_12_0_stall_21;
  reg        [15:0]   io_in_r_bypass_regNext_12_1_data_21;
  reg                 io_in_r_bypass_regNext_12_1_load_store_21;
  reg                 io_in_r_bypass_regNext_12_1_df_is_ws_21;
  reg                 io_in_r_bypass_regNext_12_1_stall_21;
  reg        [15:0]   io_in_r_bypass_regNext_12_2_data_21;
  reg                 io_in_r_bypass_regNext_12_2_load_store_21;
  reg                 io_in_r_bypass_regNext_12_2_df_is_ws_21;
  reg                 io_in_r_bypass_regNext_12_2_stall_21;
  reg        [15:0]   io_in_r_bypass_regNext_12_3_data_21;
  reg                 io_in_r_bypass_regNext_12_3_load_store_21;
  reg                 io_in_r_bypass_regNext_12_3_df_is_ws_21;
  reg                 io_in_r_bypass_regNext_12_3_stall_21;
  reg        [15:0]   io_in_r_bypass_regNext_13_0_data_21;
  reg                 io_in_r_bypass_regNext_13_0_load_store_21;
  reg                 io_in_r_bypass_regNext_13_0_df_is_ws_21;
  reg                 io_in_r_bypass_regNext_13_0_stall_21;
  reg        [15:0]   io_in_r_bypass_regNext_13_1_data_21;
  reg                 io_in_r_bypass_regNext_13_1_load_store_21;
  reg                 io_in_r_bypass_regNext_13_1_df_is_ws_21;
  reg                 io_in_r_bypass_regNext_13_1_stall_21;
  reg        [15:0]   io_in_r_bypass_regNext_13_2_data_21;
  reg                 io_in_r_bypass_regNext_13_2_load_store_21;
  reg                 io_in_r_bypass_regNext_13_2_df_is_ws_21;
  reg                 io_in_r_bypass_regNext_13_2_stall_21;
  reg        [15:0]   io_in_r_bypass_regNext_13_3_data_21;
  reg                 io_in_r_bypass_regNext_13_3_load_store_21;
  reg                 io_in_r_bypass_regNext_13_3_df_is_ws_21;
  reg                 io_in_r_bypass_regNext_13_3_stall_21;
  reg        [15:0]   io_in_r_bypass_regNext_14_0_data_21;
  reg                 io_in_r_bypass_regNext_14_0_load_store_21;
  reg                 io_in_r_bypass_regNext_14_0_df_is_ws_21;
  reg                 io_in_r_bypass_regNext_14_0_stall_21;
  reg        [15:0]   io_in_r_bypass_regNext_14_1_data_21;
  reg                 io_in_r_bypass_regNext_14_1_load_store_21;
  reg                 io_in_r_bypass_regNext_14_1_df_is_ws_21;
  reg                 io_in_r_bypass_regNext_14_1_stall_21;
  reg        [15:0]   io_in_r_bypass_regNext_14_2_data_21;
  reg                 io_in_r_bypass_regNext_14_2_load_store_21;
  reg                 io_in_r_bypass_regNext_14_2_df_is_ws_21;
  reg                 io_in_r_bypass_regNext_14_2_stall_21;
  reg        [15:0]   io_in_r_bypass_regNext_14_3_data_21;
  reg                 io_in_r_bypass_regNext_14_3_load_store_21;
  reg                 io_in_r_bypass_regNext_14_3_df_is_ws_21;
  reg                 io_in_r_bypass_regNext_14_3_stall_21;
  reg        [15:0]   io_in_r_bypass_regNext_15_0_data_21;
  reg                 io_in_r_bypass_regNext_15_0_load_store_21;
  reg                 io_in_r_bypass_regNext_15_0_df_is_ws_21;
  reg                 io_in_r_bypass_regNext_15_0_stall_21;
  reg        [15:0]   io_in_r_bypass_regNext_15_1_data_21;
  reg                 io_in_r_bypass_regNext_15_1_load_store_21;
  reg                 io_in_r_bypass_regNext_15_1_df_is_ws_21;
  reg                 io_in_r_bypass_regNext_15_1_stall_21;
  reg        [15:0]   io_in_r_bypass_regNext_15_2_data_21;
  reg                 io_in_r_bypass_regNext_15_2_load_store_21;
  reg                 io_in_r_bypass_regNext_15_2_df_is_ws_21;
  reg                 io_in_r_bypass_regNext_15_2_stall_21;
  reg        [15:0]   io_in_r_bypass_regNext_15_3_data_21;
  reg                 io_in_r_bypass_regNext_15_3_load_store_21;
  reg                 io_in_r_bypass_regNext_15_3_df_is_ws_21;
  reg                 io_in_r_bypass_regNext_15_3_stall_21;
  reg        [15:0]   io_in_r_bypass_regNext_16_0_data_21;
  reg                 io_in_r_bypass_regNext_16_0_load_store_21;
  reg                 io_in_r_bypass_regNext_16_0_df_is_ws_21;
  reg                 io_in_r_bypass_regNext_16_0_stall_21;
  reg        [15:0]   io_in_r_bypass_regNext_16_1_data_21;
  reg                 io_in_r_bypass_regNext_16_1_load_store_21;
  reg                 io_in_r_bypass_regNext_16_1_df_is_ws_21;
  reg                 io_in_r_bypass_regNext_16_1_stall_21;
  reg        [15:0]   io_in_r_bypass_regNext_16_2_data_21;
  reg                 io_in_r_bypass_regNext_16_2_load_store_21;
  reg                 io_in_r_bypass_regNext_16_2_df_is_ws_21;
  reg                 io_in_r_bypass_regNext_16_2_stall_21;
  reg        [15:0]   io_in_r_bypass_regNext_16_3_data_21;
  reg                 io_in_r_bypass_regNext_16_3_load_store_21;
  reg                 io_in_r_bypass_regNext_16_3_df_is_ws_21;
  reg                 io_in_r_bypass_regNext_16_3_stall_21;
  reg        [15:0]   io_in_r_bypass_regNext_17_0_data_21;
  reg                 io_in_r_bypass_regNext_17_0_load_store_21;
  reg                 io_in_r_bypass_regNext_17_0_df_is_ws_21;
  reg                 io_in_r_bypass_regNext_17_0_stall_21;
  reg        [15:0]   io_in_r_bypass_regNext_17_1_data_21;
  reg                 io_in_r_bypass_regNext_17_1_load_store_21;
  reg                 io_in_r_bypass_regNext_17_1_df_is_ws_21;
  reg                 io_in_r_bypass_regNext_17_1_stall_21;
  reg        [15:0]   io_in_r_bypass_regNext_17_2_data_21;
  reg                 io_in_r_bypass_regNext_17_2_load_store_21;
  reg                 io_in_r_bypass_regNext_17_2_df_is_ws_21;
  reg                 io_in_r_bypass_regNext_17_2_stall_21;
  reg        [15:0]   io_in_r_bypass_regNext_17_3_data_21;
  reg                 io_in_r_bypass_regNext_17_3_load_store_21;
  reg                 io_in_r_bypass_regNext_17_3_df_is_ws_21;
  reg                 io_in_r_bypass_regNext_17_3_stall_21;
  reg        [15:0]   io_in_r_bypass_regNext_18_0_data_21;
  reg                 io_in_r_bypass_regNext_18_0_load_store_21;
  reg                 io_in_r_bypass_regNext_18_0_df_is_ws_21;
  reg                 io_in_r_bypass_regNext_18_0_stall_21;
  reg        [15:0]   io_in_r_bypass_regNext_18_1_data_21;
  reg                 io_in_r_bypass_regNext_18_1_load_store_21;
  reg                 io_in_r_bypass_regNext_18_1_df_is_ws_21;
  reg                 io_in_r_bypass_regNext_18_1_stall_21;
  reg        [15:0]   io_in_r_bypass_regNext_18_2_data_21;
  reg                 io_in_r_bypass_regNext_18_2_load_store_21;
  reg                 io_in_r_bypass_regNext_18_2_df_is_ws_21;
  reg                 io_in_r_bypass_regNext_18_2_stall_21;
  reg        [15:0]   io_in_r_bypass_regNext_18_3_data_21;
  reg                 io_in_r_bypass_regNext_18_3_load_store_21;
  reg                 io_in_r_bypass_regNext_18_3_df_is_ws_21;
  reg                 io_in_r_bypass_regNext_18_3_stall_21;
  reg        [15:0]   io_in_r_bypass_regNext_19_0_data_21;
  reg                 io_in_r_bypass_regNext_19_0_load_store_21;
  reg                 io_in_r_bypass_regNext_19_0_df_is_ws_21;
  reg                 io_in_r_bypass_regNext_19_0_stall_21;
  reg        [15:0]   io_in_r_bypass_regNext_19_1_data_21;
  reg                 io_in_r_bypass_regNext_19_1_load_store_21;
  reg                 io_in_r_bypass_regNext_19_1_df_is_ws_21;
  reg                 io_in_r_bypass_regNext_19_1_stall_21;
  reg        [15:0]   io_in_r_bypass_regNext_19_2_data_21;
  reg                 io_in_r_bypass_regNext_19_2_load_store_21;
  reg                 io_in_r_bypass_regNext_19_2_df_is_ws_21;
  reg                 io_in_r_bypass_regNext_19_2_stall_21;
  reg        [15:0]   io_in_r_bypass_regNext_19_3_data_21;
  reg                 io_in_r_bypass_regNext_19_3_load_store_21;
  reg                 io_in_r_bypass_regNext_19_3_df_is_ws_21;
  reg                 io_in_r_bypass_regNext_19_3_stall_21;
  reg        [15:0]   io_in_r_bypass_regNext_20_0_data_21;
  reg                 io_in_r_bypass_regNext_20_0_load_store_21;
  reg                 io_in_r_bypass_regNext_20_0_df_is_ws_21;
  reg                 io_in_r_bypass_regNext_20_0_stall_21;
  reg        [15:0]   io_in_r_bypass_regNext_20_1_data_21;
  reg                 io_in_r_bypass_regNext_20_1_load_store_21;
  reg                 io_in_r_bypass_regNext_20_1_df_is_ws_21;
  reg                 io_in_r_bypass_regNext_20_1_stall_21;
  reg        [15:0]   io_in_r_bypass_regNext_20_2_data_21;
  reg                 io_in_r_bypass_regNext_20_2_load_store_21;
  reg                 io_in_r_bypass_regNext_20_2_df_is_ws_21;
  reg                 io_in_r_bypass_regNext_20_2_stall_21;
  reg        [15:0]   io_in_r_bypass_regNext_20_3_data_21;
  reg                 io_in_r_bypass_regNext_20_3_load_store_21;
  reg                 io_in_r_bypass_regNext_20_3_df_is_ws_21;
  reg                 io_in_r_bypass_regNext_20_3_stall_21;
  reg        [15:0]   io_in_r_bypass_regNext_21_0_data_21;
  reg                 io_in_r_bypass_regNext_21_0_load_store_21;
  reg                 io_in_r_bypass_regNext_21_0_df_is_ws_21;
  reg                 io_in_r_bypass_regNext_21_0_stall_21;
  reg        [15:0]   io_in_r_bypass_regNext_21_1_data_21;
  reg                 io_in_r_bypass_regNext_21_1_load_store_21;
  reg                 io_in_r_bypass_regNext_21_1_df_is_ws_21;
  reg                 io_in_r_bypass_regNext_21_1_stall_21;
  reg        [15:0]   io_in_r_bypass_regNext_21_2_data_21;
  reg                 io_in_r_bypass_regNext_21_2_load_store_21;
  reg                 io_in_r_bypass_regNext_21_2_df_is_ws_21;
  reg                 io_in_r_bypass_regNext_21_2_stall_21;
  reg        [15:0]   io_in_r_bypass_regNext_21_3_data_21;
  reg                 io_in_r_bypass_regNext_21_3_load_store_21;
  reg                 io_in_r_bypass_regNext_21_3_df_is_ws_21;
  reg                 io_in_r_bypass_regNext_21_3_stall_21;
  reg        [15:0]   io_in_r_bypass_regNext_22_0_data_21;
  reg                 io_in_r_bypass_regNext_22_0_load_store_21;
  reg                 io_in_r_bypass_regNext_22_0_df_is_ws_21;
  reg                 io_in_r_bypass_regNext_22_0_stall_21;
  reg        [15:0]   io_in_r_bypass_regNext_22_1_data_21;
  reg                 io_in_r_bypass_regNext_22_1_load_store_21;
  reg                 io_in_r_bypass_regNext_22_1_df_is_ws_21;
  reg                 io_in_r_bypass_regNext_22_1_stall_21;
  reg        [15:0]   io_in_r_bypass_regNext_22_2_data_21;
  reg                 io_in_r_bypass_regNext_22_2_load_store_21;
  reg                 io_in_r_bypass_regNext_22_2_df_is_ws_21;
  reg                 io_in_r_bypass_regNext_22_2_stall_21;
  reg        [15:0]   io_in_r_bypass_regNext_22_3_data_21;
  reg                 io_in_r_bypass_regNext_22_3_load_store_21;
  reg                 io_in_r_bypass_regNext_22_3_df_is_ws_21;
  reg                 io_in_r_bypass_regNext_22_3_stall_21;
  reg        [15:0]   io_in_r_bypass_regNext_23_0_data_21;
  reg                 io_in_r_bypass_regNext_23_0_load_store_21;
  reg                 io_in_r_bypass_regNext_23_0_df_is_ws_21;
  reg                 io_in_r_bypass_regNext_23_0_stall_21;
  reg        [15:0]   io_in_r_bypass_regNext_23_1_data_21;
  reg                 io_in_r_bypass_regNext_23_1_load_store_21;
  reg                 io_in_r_bypass_regNext_23_1_df_is_ws_21;
  reg                 io_in_r_bypass_regNext_23_1_stall_21;
  reg        [15:0]   io_in_r_bypass_regNext_23_2_data_21;
  reg                 io_in_r_bypass_regNext_23_2_load_store_21;
  reg                 io_in_r_bypass_regNext_23_2_df_is_ws_21;
  reg                 io_in_r_bypass_regNext_23_2_stall_21;
  reg        [15:0]   io_in_r_bypass_regNext_23_3_data_21;
  reg                 io_in_r_bypass_regNext_23_3_load_store_21;
  reg                 io_in_r_bypass_regNext_23_3_df_is_ws_21;
  reg                 io_in_r_bypass_regNext_23_3_stall_21;
  reg        [15:0]   io_in_r_bypass_regNext_24_0_data_21;
  reg                 io_in_r_bypass_regNext_24_0_load_store_21;
  reg                 io_in_r_bypass_regNext_24_0_df_is_ws_21;
  reg                 io_in_r_bypass_regNext_24_0_stall_21;
  reg        [15:0]   io_in_r_bypass_regNext_24_1_data_21;
  reg                 io_in_r_bypass_regNext_24_1_load_store_21;
  reg                 io_in_r_bypass_regNext_24_1_df_is_ws_21;
  reg                 io_in_r_bypass_regNext_24_1_stall_21;
  reg        [15:0]   io_in_r_bypass_regNext_24_2_data_21;
  reg                 io_in_r_bypass_regNext_24_2_load_store_21;
  reg                 io_in_r_bypass_regNext_24_2_df_is_ws_21;
  reg                 io_in_r_bypass_regNext_24_2_stall_21;
  reg        [15:0]   io_in_r_bypass_regNext_24_3_data_21;
  reg                 io_in_r_bypass_regNext_24_3_load_store_21;
  reg                 io_in_r_bypass_regNext_24_3_df_is_ws_21;
  reg                 io_in_r_bypass_regNext_24_3_stall_21;
  reg        [15:0]   io_in_r_bypass_regNext_25_0_data_21;
  reg                 io_in_r_bypass_regNext_25_0_load_store_21;
  reg                 io_in_r_bypass_regNext_25_0_df_is_ws_21;
  reg                 io_in_r_bypass_regNext_25_0_stall_21;
  reg        [15:0]   io_in_r_bypass_regNext_25_1_data_21;
  reg                 io_in_r_bypass_regNext_25_1_load_store_21;
  reg                 io_in_r_bypass_regNext_25_1_df_is_ws_21;
  reg                 io_in_r_bypass_regNext_25_1_stall_21;
  reg        [15:0]   io_in_r_bypass_regNext_25_2_data_21;
  reg                 io_in_r_bypass_regNext_25_2_load_store_21;
  reg                 io_in_r_bypass_regNext_25_2_df_is_ws_21;
  reg                 io_in_r_bypass_regNext_25_2_stall_21;
  reg        [15:0]   io_in_r_bypass_regNext_25_3_data_21;
  reg                 io_in_r_bypass_regNext_25_3_load_store_21;
  reg                 io_in_r_bypass_regNext_25_3_df_is_ws_21;
  reg                 io_in_r_bypass_regNext_25_3_stall_21;
  reg        [15:0]   io_in_r_bypass_regNext_26_0_data_21;
  reg                 io_in_r_bypass_regNext_26_0_load_store_21;
  reg                 io_in_r_bypass_regNext_26_0_df_is_ws_21;
  reg                 io_in_r_bypass_regNext_26_0_stall_21;
  reg        [15:0]   io_in_r_bypass_regNext_26_1_data_21;
  reg                 io_in_r_bypass_regNext_26_1_load_store_21;
  reg                 io_in_r_bypass_regNext_26_1_df_is_ws_21;
  reg                 io_in_r_bypass_regNext_26_1_stall_21;
  reg        [15:0]   io_in_r_bypass_regNext_26_2_data_21;
  reg                 io_in_r_bypass_regNext_26_2_load_store_21;
  reg                 io_in_r_bypass_regNext_26_2_df_is_ws_21;
  reg                 io_in_r_bypass_regNext_26_2_stall_21;
  reg        [15:0]   io_in_r_bypass_regNext_26_3_data_21;
  reg                 io_in_r_bypass_regNext_26_3_load_store_21;
  reg                 io_in_r_bypass_regNext_26_3_df_is_ws_21;
  reg                 io_in_r_bypass_regNext_26_3_stall_21;
  reg        [15:0]   io_in_r_bypass_regNext_27_0_data_21;
  reg                 io_in_r_bypass_regNext_27_0_load_store_21;
  reg                 io_in_r_bypass_regNext_27_0_df_is_ws_21;
  reg                 io_in_r_bypass_regNext_27_0_stall_21;
  reg        [15:0]   io_in_r_bypass_regNext_27_1_data_21;
  reg                 io_in_r_bypass_regNext_27_1_load_store_21;
  reg                 io_in_r_bypass_regNext_27_1_df_is_ws_21;
  reg                 io_in_r_bypass_regNext_27_1_stall_21;
  reg        [15:0]   io_in_r_bypass_regNext_27_2_data_21;
  reg                 io_in_r_bypass_regNext_27_2_load_store_21;
  reg                 io_in_r_bypass_regNext_27_2_df_is_ws_21;
  reg                 io_in_r_bypass_regNext_27_2_stall_21;
  reg        [15:0]   io_in_r_bypass_regNext_27_3_data_21;
  reg                 io_in_r_bypass_regNext_27_3_load_store_21;
  reg                 io_in_r_bypass_regNext_27_3_df_is_ws_21;
  reg                 io_in_r_bypass_regNext_27_3_stall_21;
  reg        [15:0]   io_in_r_bypass_regNext_28_0_data_21;
  reg                 io_in_r_bypass_regNext_28_0_load_store_21;
  reg                 io_in_r_bypass_regNext_28_0_df_is_ws_21;
  reg                 io_in_r_bypass_regNext_28_0_stall_21;
  reg        [15:0]   io_in_r_bypass_regNext_28_1_data_21;
  reg                 io_in_r_bypass_regNext_28_1_load_store_21;
  reg                 io_in_r_bypass_regNext_28_1_df_is_ws_21;
  reg                 io_in_r_bypass_regNext_28_1_stall_21;
  reg        [15:0]   io_in_r_bypass_regNext_28_2_data_21;
  reg                 io_in_r_bypass_regNext_28_2_load_store_21;
  reg                 io_in_r_bypass_regNext_28_2_df_is_ws_21;
  reg                 io_in_r_bypass_regNext_28_2_stall_21;
  reg        [15:0]   io_in_r_bypass_regNext_28_3_data_21;
  reg                 io_in_r_bypass_regNext_28_3_load_store_21;
  reg                 io_in_r_bypass_regNext_28_3_df_is_ws_21;
  reg                 io_in_r_bypass_regNext_28_3_stall_21;
  reg        [15:0]   io_in_r_bypass_regNext_29_0_data_21;
  reg                 io_in_r_bypass_regNext_29_0_load_store_21;
  reg                 io_in_r_bypass_regNext_29_0_df_is_ws_21;
  reg                 io_in_r_bypass_regNext_29_0_stall_21;
  reg        [15:0]   io_in_r_bypass_regNext_29_1_data_21;
  reg                 io_in_r_bypass_regNext_29_1_load_store_21;
  reg                 io_in_r_bypass_regNext_29_1_df_is_ws_21;
  reg                 io_in_r_bypass_regNext_29_1_stall_21;
  reg        [15:0]   io_in_r_bypass_regNext_29_2_data_21;
  reg                 io_in_r_bypass_regNext_29_2_load_store_21;
  reg                 io_in_r_bypass_regNext_29_2_df_is_ws_21;
  reg                 io_in_r_bypass_regNext_29_2_stall_21;
  reg        [15:0]   io_in_r_bypass_regNext_29_3_data_21;
  reg                 io_in_r_bypass_regNext_29_3_load_store_21;
  reg                 io_in_r_bypass_regNext_29_3_df_is_ws_21;
  reg                 io_in_r_bypass_regNext_29_3_stall_21;
  reg        [15:0]   io_in_r_bypass_regNext_30_0_data_21;
  reg                 io_in_r_bypass_regNext_30_0_load_store_21;
  reg                 io_in_r_bypass_regNext_30_0_df_is_ws_21;
  reg                 io_in_r_bypass_regNext_30_0_stall_21;
  reg        [15:0]   io_in_r_bypass_regNext_30_1_data_21;
  reg                 io_in_r_bypass_regNext_30_1_load_store_21;
  reg                 io_in_r_bypass_regNext_30_1_df_is_ws_21;
  reg                 io_in_r_bypass_regNext_30_1_stall_21;
  reg        [15:0]   io_in_r_bypass_regNext_30_2_data_21;
  reg                 io_in_r_bypass_regNext_30_2_load_store_21;
  reg                 io_in_r_bypass_regNext_30_2_df_is_ws_21;
  reg                 io_in_r_bypass_regNext_30_2_stall_21;
  reg        [15:0]   io_in_r_bypass_regNext_30_3_data_21;
  reg                 io_in_r_bypass_regNext_30_3_load_store_21;
  reg                 io_in_r_bypass_regNext_30_3_df_is_ws_21;
  reg                 io_in_r_bypass_regNext_30_3_stall_21;
  reg        [15:0]   io_in_r_bypass_regNext_31_0_data_21;
  reg                 io_in_r_bypass_regNext_31_0_load_store_21;
  reg                 io_in_r_bypass_regNext_31_0_df_is_ws_21;
  reg                 io_in_r_bypass_regNext_31_0_stall_21;
  reg        [15:0]   io_in_r_bypass_regNext_31_1_data_21;
  reg                 io_in_r_bypass_regNext_31_1_load_store_21;
  reg                 io_in_r_bypass_regNext_31_1_df_is_ws_21;
  reg                 io_in_r_bypass_regNext_31_1_stall_21;
  reg        [15:0]   io_in_r_bypass_regNext_31_2_data_21;
  reg                 io_in_r_bypass_regNext_31_2_load_store_21;
  reg                 io_in_r_bypass_regNext_31_2_df_is_ws_21;
  reg                 io_in_r_bypass_regNext_31_2_stall_21;
  reg        [15:0]   io_in_r_bypass_regNext_31_3_data_21;
  reg                 io_in_r_bypass_regNext_31_3_load_store_21;
  reg                 io_in_r_bypass_regNext_31_3_df_is_ws_21;
  reg                 io_in_r_bypass_regNext_31_3_stall_21;
  reg        [15:0]   io_in_r_bypass_regNext_0_0_data_22;
  reg                 io_in_r_bypass_regNext_0_0_load_store_22;
  reg                 io_in_r_bypass_regNext_0_0_df_is_ws_22;
  reg                 io_in_r_bypass_regNext_0_0_stall_22;
  reg        [15:0]   io_in_r_bypass_regNext_0_1_data_22;
  reg                 io_in_r_bypass_regNext_0_1_load_store_22;
  reg                 io_in_r_bypass_regNext_0_1_df_is_ws_22;
  reg                 io_in_r_bypass_regNext_0_1_stall_22;
  reg        [15:0]   io_in_r_bypass_regNext_0_2_data_22;
  reg                 io_in_r_bypass_regNext_0_2_load_store_22;
  reg                 io_in_r_bypass_regNext_0_2_df_is_ws_22;
  reg                 io_in_r_bypass_regNext_0_2_stall_22;
  reg        [15:0]   io_in_r_bypass_regNext_0_3_data_22;
  reg                 io_in_r_bypass_regNext_0_3_load_store_22;
  reg                 io_in_r_bypass_regNext_0_3_df_is_ws_22;
  reg                 io_in_r_bypass_regNext_0_3_stall_22;
  reg        [15:0]   io_in_r_bypass_regNext_1_0_data_22;
  reg                 io_in_r_bypass_regNext_1_0_load_store_22;
  reg                 io_in_r_bypass_regNext_1_0_df_is_ws_22;
  reg                 io_in_r_bypass_regNext_1_0_stall_22;
  reg        [15:0]   io_in_r_bypass_regNext_1_1_data_22;
  reg                 io_in_r_bypass_regNext_1_1_load_store_22;
  reg                 io_in_r_bypass_regNext_1_1_df_is_ws_22;
  reg                 io_in_r_bypass_regNext_1_1_stall_22;
  reg        [15:0]   io_in_r_bypass_regNext_1_2_data_22;
  reg                 io_in_r_bypass_regNext_1_2_load_store_22;
  reg                 io_in_r_bypass_regNext_1_2_df_is_ws_22;
  reg                 io_in_r_bypass_regNext_1_2_stall_22;
  reg        [15:0]   io_in_r_bypass_regNext_1_3_data_22;
  reg                 io_in_r_bypass_regNext_1_3_load_store_22;
  reg                 io_in_r_bypass_regNext_1_3_df_is_ws_22;
  reg                 io_in_r_bypass_regNext_1_3_stall_22;
  reg        [15:0]   io_in_r_bypass_regNext_2_0_data_22;
  reg                 io_in_r_bypass_regNext_2_0_load_store_22;
  reg                 io_in_r_bypass_regNext_2_0_df_is_ws_22;
  reg                 io_in_r_bypass_regNext_2_0_stall_22;
  reg        [15:0]   io_in_r_bypass_regNext_2_1_data_22;
  reg                 io_in_r_bypass_regNext_2_1_load_store_22;
  reg                 io_in_r_bypass_regNext_2_1_df_is_ws_22;
  reg                 io_in_r_bypass_regNext_2_1_stall_22;
  reg        [15:0]   io_in_r_bypass_regNext_2_2_data_22;
  reg                 io_in_r_bypass_regNext_2_2_load_store_22;
  reg                 io_in_r_bypass_regNext_2_2_df_is_ws_22;
  reg                 io_in_r_bypass_regNext_2_2_stall_22;
  reg        [15:0]   io_in_r_bypass_regNext_2_3_data_22;
  reg                 io_in_r_bypass_regNext_2_3_load_store_22;
  reg                 io_in_r_bypass_regNext_2_3_df_is_ws_22;
  reg                 io_in_r_bypass_regNext_2_3_stall_22;
  reg        [15:0]   io_in_r_bypass_regNext_3_0_data_22;
  reg                 io_in_r_bypass_regNext_3_0_load_store_22;
  reg                 io_in_r_bypass_regNext_3_0_df_is_ws_22;
  reg                 io_in_r_bypass_regNext_3_0_stall_22;
  reg        [15:0]   io_in_r_bypass_regNext_3_1_data_22;
  reg                 io_in_r_bypass_regNext_3_1_load_store_22;
  reg                 io_in_r_bypass_regNext_3_1_df_is_ws_22;
  reg                 io_in_r_bypass_regNext_3_1_stall_22;
  reg        [15:0]   io_in_r_bypass_regNext_3_2_data_22;
  reg                 io_in_r_bypass_regNext_3_2_load_store_22;
  reg                 io_in_r_bypass_regNext_3_2_df_is_ws_22;
  reg                 io_in_r_bypass_regNext_3_2_stall_22;
  reg        [15:0]   io_in_r_bypass_regNext_3_3_data_22;
  reg                 io_in_r_bypass_regNext_3_3_load_store_22;
  reg                 io_in_r_bypass_regNext_3_3_df_is_ws_22;
  reg                 io_in_r_bypass_regNext_3_3_stall_22;
  reg        [15:0]   io_in_r_bypass_regNext_4_0_data_22;
  reg                 io_in_r_bypass_regNext_4_0_load_store_22;
  reg                 io_in_r_bypass_regNext_4_0_df_is_ws_22;
  reg                 io_in_r_bypass_regNext_4_0_stall_22;
  reg        [15:0]   io_in_r_bypass_regNext_4_1_data_22;
  reg                 io_in_r_bypass_regNext_4_1_load_store_22;
  reg                 io_in_r_bypass_regNext_4_1_df_is_ws_22;
  reg                 io_in_r_bypass_regNext_4_1_stall_22;
  reg        [15:0]   io_in_r_bypass_regNext_4_2_data_22;
  reg                 io_in_r_bypass_regNext_4_2_load_store_22;
  reg                 io_in_r_bypass_regNext_4_2_df_is_ws_22;
  reg                 io_in_r_bypass_regNext_4_2_stall_22;
  reg        [15:0]   io_in_r_bypass_regNext_4_3_data_22;
  reg                 io_in_r_bypass_regNext_4_3_load_store_22;
  reg                 io_in_r_bypass_regNext_4_3_df_is_ws_22;
  reg                 io_in_r_bypass_regNext_4_3_stall_22;
  reg        [15:0]   io_in_r_bypass_regNext_5_0_data_22;
  reg                 io_in_r_bypass_regNext_5_0_load_store_22;
  reg                 io_in_r_bypass_regNext_5_0_df_is_ws_22;
  reg                 io_in_r_bypass_regNext_5_0_stall_22;
  reg        [15:0]   io_in_r_bypass_regNext_5_1_data_22;
  reg                 io_in_r_bypass_regNext_5_1_load_store_22;
  reg                 io_in_r_bypass_regNext_5_1_df_is_ws_22;
  reg                 io_in_r_bypass_regNext_5_1_stall_22;
  reg        [15:0]   io_in_r_bypass_regNext_5_2_data_22;
  reg                 io_in_r_bypass_regNext_5_2_load_store_22;
  reg                 io_in_r_bypass_regNext_5_2_df_is_ws_22;
  reg                 io_in_r_bypass_regNext_5_2_stall_22;
  reg        [15:0]   io_in_r_bypass_regNext_5_3_data_22;
  reg                 io_in_r_bypass_regNext_5_3_load_store_22;
  reg                 io_in_r_bypass_regNext_5_3_df_is_ws_22;
  reg                 io_in_r_bypass_regNext_5_3_stall_22;
  reg        [15:0]   io_in_r_bypass_regNext_6_0_data_22;
  reg                 io_in_r_bypass_regNext_6_0_load_store_22;
  reg                 io_in_r_bypass_regNext_6_0_df_is_ws_22;
  reg                 io_in_r_bypass_regNext_6_0_stall_22;
  reg        [15:0]   io_in_r_bypass_regNext_6_1_data_22;
  reg                 io_in_r_bypass_regNext_6_1_load_store_22;
  reg                 io_in_r_bypass_regNext_6_1_df_is_ws_22;
  reg                 io_in_r_bypass_regNext_6_1_stall_22;
  reg        [15:0]   io_in_r_bypass_regNext_6_2_data_22;
  reg                 io_in_r_bypass_regNext_6_2_load_store_22;
  reg                 io_in_r_bypass_regNext_6_2_df_is_ws_22;
  reg                 io_in_r_bypass_regNext_6_2_stall_22;
  reg        [15:0]   io_in_r_bypass_regNext_6_3_data_22;
  reg                 io_in_r_bypass_regNext_6_3_load_store_22;
  reg                 io_in_r_bypass_regNext_6_3_df_is_ws_22;
  reg                 io_in_r_bypass_regNext_6_3_stall_22;
  reg        [15:0]   io_in_r_bypass_regNext_7_0_data_22;
  reg                 io_in_r_bypass_regNext_7_0_load_store_22;
  reg                 io_in_r_bypass_regNext_7_0_df_is_ws_22;
  reg                 io_in_r_bypass_regNext_7_0_stall_22;
  reg        [15:0]   io_in_r_bypass_regNext_7_1_data_22;
  reg                 io_in_r_bypass_regNext_7_1_load_store_22;
  reg                 io_in_r_bypass_regNext_7_1_df_is_ws_22;
  reg                 io_in_r_bypass_regNext_7_1_stall_22;
  reg        [15:0]   io_in_r_bypass_regNext_7_2_data_22;
  reg                 io_in_r_bypass_regNext_7_2_load_store_22;
  reg                 io_in_r_bypass_regNext_7_2_df_is_ws_22;
  reg                 io_in_r_bypass_regNext_7_2_stall_22;
  reg        [15:0]   io_in_r_bypass_regNext_7_3_data_22;
  reg                 io_in_r_bypass_regNext_7_3_load_store_22;
  reg                 io_in_r_bypass_regNext_7_3_df_is_ws_22;
  reg                 io_in_r_bypass_regNext_7_3_stall_22;
  reg        [15:0]   io_in_r_bypass_regNext_8_0_data_22;
  reg                 io_in_r_bypass_regNext_8_0_load_store_22;
  reg                 io_in_r_bypass_regNext_8_0_df_is_ws_22;
  reg                 io_in_r_bypass_regNext_8_0_stall_22;
  reg        [15:0]   io_in_r_bypass_regNext_8_1_data_22;
  reg                 io_in_r_bypass_regNext_8_1_load_store_22;
  reg                 io_in_r_bypass_regNext_8_1_df_is_ws_22;
  reg                 io_in_r_bypass_regNext_8_1_stall_22;
  reg        [15:0]   io_in_r_bypass_regNext_8_2_data_22;
  reg                 io_in_r_bypass_regNext_8_2_load_store_22;
  reg                 io_in_r_bypass_regNext_8_2_df_is_ws_22;
  reg                 io_in_r_bypass_regNext_8_2_stall_22;
  reg        [15:0]   io_in_r_bypass_regNext_8_3_data_22;
  reg                 io_in_r_bypass_regNext_8_3_load_store_22;
  reg                 io_in_r_bypass_regNext_8_3_df_is_ws_22;
  reg                 io_in_r_bypass_regNext_8_3_stall_22;
  reg        [15:0]   io_in_r_bypass_regNext_9_0_data_22;
  reg                 io_in_r_bypass_regNext_9_0_load_store_22;
  reg                 io_in_r_bypass_regNext_9_0_df_is_ws_22;
  reg                 io_in_r_bypass_regNext_9_0_stall_22;
  reg        [15:0]   io_in_r_bypass_regNext_9_1_data_22;
  reg                 io_in_r_bypass_regNext_9_1_load_store_22;
  reg                 io_in_r_bypass_regNext_9_1_df_is_ws_22;
  reg                 io_in_r_bypass_regNext_9_1_stall_22;
  reg        [15:0]   io_in_r_bypass_regNext_9_2_data_22;
  reg                 io_in_r_bypass_regNext_9_2_load_store_22;
  reg                 io_in_r_bypass_regNext_9_2_df_is_ws_22;
  reg                 io_in_r_bypass_regNext_9_2_stall_22;
  reg        [15:0]   io_in_r_bypass_regNext_9_3_data_22;
  reg                 io_in_r_bypass_regNext_9_3_load_store_22;
  reg                 io_in_r_bypass_regNext_9_3_df_is_ws_22;
  reg                 io_in_r_bypass_regNext_9_3_stall_22;
  reg        [15:0]   io_in_r_bypass_regNext_10_0_data_22;
  reg                 io_in_r_bypass_regNext_10_0_load_store_22;
  reg                 io_in_r_bypass_regNext_10_0_df_is_ws_22;
  reg                 io_in_r_bypass_regNext_10_0_stall_22;
  reg        [15:0]   io_in_r_bypass_regNext_10_1_data_22;
  reg                 io_in_r_bypass_regNext_10_1_load_store_22;
  reg                 io_in_r_bypass_regNext_10_1_df_is_ws_22;
  reg                 io_in_r_bypass_regNext_10_1_stall_22;
  reg        [15:0]   io_in_r_bypass_regNext_10_2_data_22;
  reg                 io_in_r_bypass_regNext_10_2_load_store_22;
  reg                 io_in_r_bypass_regNext_10_2_df_is_ws_22;
  reg                 io_in_r_bypass_regNext_10_2_stall_22;
  reg        [15:0]   io_in_r_bypass_regNext_10_3_data_22;
  reg                 io_in_r_bypass_regNext_10_3_load_store_22;
  reg                 io_in_r_bypass_regNext_10_3_df_is_ws_22;
  reg                 io_in_r_bypass_regNext_10_3_stall_22;
  reg        [15:0]   io_in_r_bypass_regNext_11_0_data_22;
  reg                 io_in_r_bypass_regNext_11_0_load_store_22;
  reg                 io_in_r_bypass_regNext_11_0_df_is_ws_22;
  reg                 io_in_r_bypass_regNext_11_0_stall_22;
  reg        [15:0]   io_in_r_bypass_regNext_11_1_data_22;
  reg                 io_in_r_bypass_regNext_11_1_load_store_22;
  reg                 io_in_r_bypass_regNext_11_1_df_is_ws_22;
  reg                 io_in_r_bypass_regNext_11_1_stall_22;
  reg        [15:0]   io_in_r_bypass_regNext_11_2_data_22;
  reg                 io_in_r_bypass_regNext_11_2_load_store_22;
  reg                 io_in_r_bypass_regNext_11_2_df_is_ws_22;
  reg                 io_in_r_bypass_regNext_11_2_stall_22;
  reg        [15:0]   io_in_r_bypass_regNext_11_3_data_22;
  reg                 io_in_r_bypass_regNext_11_3_load_store_22;
  reg                 io_in_r_bypass_regNext_11_3_df_is_ws_22;
  reg                 io_in_r_bypass_regNext_11_3_stall_22;
  reg        [15:0]   io_in_r_bypass_regNext_12_0_data_22;
  reg                 io_in_r_bypass_regNext_12_0_load_store_22;
  reg                 io_in_r_bypass_regNext_12_0_df_is_ws_22;
  reg                 io_in_r_bypass_regNext_12_0_stall_22;
  reg        [15:0]   io_in_r_bypass_regNext_12_1_data_22;
  reg                 io_in_r_bypass_regNext_12_1_load_store_22;
  reg                 io_in_r_bypass_regNext_12_1_df_is_ws_22;
  reg                 io_in_r_bypass_regNext_12_1_stall_22;
  reg        [15:0]   io_in_r_bypass_regNext_12_2_data_22;
  reg                 io_in_r_bypass_regNext_12_2_load_store_22;
  reg                 io_in_r_bypass_regNext_12_2_df_is_ws_22;
  reg                 io_in_r_bypass_regNext_12_2_stall_22;
  reg        [15:0]   io_in_r_bypass_regNext_12_3_data_22;
  reg                 io_in_r_bypass_regNext_12_3_load_store_22;
  reg                 io_in_r_bypass_regNext_12_3_df_is_ws_22;
  reg                 io_in_r_bypass_regNext_12_3_stall_22;
  reg        [15:0]   io_in_r_bypass_regNext_13_0_data_22;
  reg                 io_in_r_bypass_regNext_13_0_load_store_22;
  reg                 io_in_r_bypass_regNext_13_0_df_is_ws_22;
  reg                 io_in_r_bypass_regNext_13_0_stall_22;
  reg        [15:0]   io_in_r_bypass_regNext_13_1_data_22;
  reg                 io_in_r_bypass_regNext_13_1_load_store_22;
  reg                 io_in_r_bypass_regNext_13_1_df_is_ws_22;
  reg                 io_in_r_bypass_regNext_13_1_stall_22;
  reg        [15:0]   io_in_r_bypass_regNext_13_2_data_22;
  reg                 io_in_r_bypass_regNext_13_2_load_store_22;
  reg                 io_in_r_bypass_regNext_13_2_df_is_ws_22;
  reg                 io_in_r_bypass_regNext_13_2_stall_22;
  reg        [15:0]   io_in_r_bypass_regNext_13_3_data_22;
  reg                 io_in_r_bypass_regNext_13_3_load_store_22;
  reg                 io_in_r_bypass_regNext_13_3_df_is_ws_22;
  reg                 io_in_r_bypass_regNext_13_3_stall_22;
  reg        [15:0]   io_in_r_bypass_regNext_14_0_data_22;
  reg                 io_in_r_bypass_regNext_14_0_load_store_22;
  reg                 io_in_r_bypass_regNext_14_0_df_is_ws_22;
  reg                 io_in_r_bypass_regNext_14_0_stall_22;
  reg        [15:0]   io_in_r_bypass_regNext_14_1_data_22;
  reg                 io_in_r_bypass_regNext_14_1_load_store_22;
  reg                 io_in_r_bypass_regNext_14_1_df_is_ws_22;
  reg                 io_in_r_bypass_regNext_14_1_stall_22;
  reg        [15:0]   io_in_r_bypass_regNext_14_2_data_22;
  reg                 io_in_r_bypass_regNext_14_2_load_store_22;
  reg                 io_in_r_bypass_regNext_14_2_df_is_ws_22;
  reg                 io_in_r_bypass_regNext_14_2_stall_22;
  reg        [15:0]   io_in_r_bypass_regNext_14_3_data_22;
  reg                 io_in_r_bypass_regNext_14_3_load_store_22;
  reg                 io_in_r_bypass_regNext_14_3_df_is_ws_22;
  reg                 io_in_r_bypass_regNext_14_3_stall_22;
  reg        [15:0]   io_in_r_bypass_regNext_15_0_data_22;
  reg                 io_in_r_bypass_regNext_15_0_load_store_22;
  reg                 io_in_r_bypass_regNext_15_0_df_is_ws_22;
  reg                 io_in_r_bypass_regNext_15_0_stall_22;
  reg        [15:0]   io_in_r_bypass_regNext_15_1_data_22;
  reg                 io_in_r_bypass_regNext_15_1_load_store_22;
  reg                 io_in_r_bypass_regNext_15_1_df_is_ws_22;
  reg                 io_in_r_bypass_regNext_15_1_stall_22;
  reg        [15:0]   io_in_r_bypass_regNext_15_2_data_22;
  reg                 io_in_r_bypass_regNext_15_2_load_store_22;
  reg                 io_in_r_bypass_regNext_15_2_df_is_ws_22;
  reg                 io_in_r_bypass_regNext_15_2_stall_22;
  reg        [15:0]   io_in_r_bypass_regNext_15_3_data_22;
  reg                 io_in_r_bypass_regNext_15_3_load_store_22;
  reg                 io_in_r_bypass_regNext_15_3_df_is_ws_22;
  reg                 io_in_r_bypass_regNext_15_3_stall_22;
  reg        [15:0]   io_in_r_bypass_regNext_16_0_data_22;
  reg                 io_in_r_bypass_regNext_16_0_load_store_22;
  reg                 io_in_r_bypass_regNext_16_0_df_is_ws_22;
  reg                 io_in_r_bypass_regNext_16_0_stall_22;
  reg        [15:0]   io_in_r_bypass_regNext_16_1_data_22;
  reg                 io_in_r_bypass_regNext_16_1_load_store_22;
  reg                 io_in_r_bypass_regNext_16_1_df_is_ws_22;
  reg                 io_in_r_bypass_regNext_16_1_stall_22;
  reg        [15:0]   io_in_r_bypass_regNext_16_2_data_22;
  reg                 io_in_r_bypass_regNext_16_2_load_store_22;
  reg                 io_in_r_bypass_regNext_16_2_df_is_ws_22;
  reg                 io_in_r_bypass_regNext_16_2_stall_22;
  reg        [15:0]   io_in_r_bypass_regNext_16_3_data_22;
  reg                 io_in_r_bypass_regNext_16_3_load_store_22;
  reg                 io_in_r_bypass_regNext_16_3_df_is_ws_22;
  reg                 io_in_r_bypass_regNext_16_3_stall_22;
  reg        [15:0]   io_in_r_bypass_regNext_17_0_data_22;
  reg                 io_in_r_bypass_regNext_17_0_load_store_22;
  reg                 io_in_r_bypass_regNext_17_0_df_is_ws_22;
  reg                 io_in_r_bypass_regNext_17_0_stall_22;
  reg        [15:0]   io_in_r_bypass_regNext_17_1_data_22;
  reg                 io_in_r_bypass_regNext_17_1_load_store_22;
  reg                 io_in_r_bypass_regNext_17_1_df_is_ws_22;
  reg                 io_in_r_bypass_regNext_17_1_stall_22;
  reg        [15:0]   io_in_r_bypass_regNext_17_2_data_22;
  reg                 io_in_r_bypass_regNext_17_2_load_store_22;
  reg                 io_in_r_bypass_regNext_17_2_df_is_ws_22;
  reg                 io_in_r_bypass_regNext_17_2_stall_22;
  reg        [15:0]   io_in_r_bypass_regNext_17_3_data_22;
  reg                 io_in_r_bypass_regNext_17_3_load_store_22;
  reg                 io_in_r_bypass_regNext_17_3_df_is_ws_22;
  reg                 io_in_r_bypass_regNext_17_3_stall_22;
  reg        [15:0]   io_in_r_bypass_regNext_18_0_data_22;
  reg                 io_in_r_bypass_regNext_18_0_load_store_22;
  reg                 io_in_r_bypass_regNext_18_0_df_is_ws_22;
  reg                 io_in_r_bypass_regNext_18_0_stall_22;
  reg        [15:0]   io_in_r_bypass_regNext_18_1_data_22;
  reg                 io_in_r_bypass_regNext_18_1_load_store_22;
  reg                 io_in_r_bypass_regNext_18_1_df_is_ws_22;
  reg                 io_in_r_bypass_regNext_18_1_stall_22;
  reg        [15:0]   io_in_r_bypass_regNext_18_2_data_22;
  reg                 io_in_r_bypass_regNext_18_2_load_store_22;
  reg                 io_in_r_bypass_regNext_18_2_df_is_ws_22;
  reg                 io_in_r_bypass_regNext_18_2_stall_22;
  reg        [15:0]   io_in_r_bypass_regNext_18_3_data_22;
  reg                 io_in_r_bypass_regNext_18_3_load_store_22;
  reg                 io_in_r_bypass_regNext_18_3_df_is_ws_22;
  reg                 io_in_r_bypass_regNext_18_3_stall_22;
  reg        [15:0]   io_in_r_bypass_regNext_19_0_data_22;
  reg                 io_in_r_bypass_regNext_19_0_load_store_22;
  reg                 io_in_r_bypass_regNext_19_0_df_is_ws_22;
  reg                 io_in_r_bypass_regNext_19_0_stall_22;
  reg        [15:0]   io_in_r_bypass_regNext_19_1_data_22;
  reg                 io_in_r_bypass_regNext_19_1_load_store_22;
  reg                 io_in_r_bypass_regNext_19_1_df_is_ws_22;
  reg                 io_in_r_bypass_regNext_19_1_stall_22;
  reg        [15:0]   io_in_r_bypass_regNext_19_2_data_22;
  reg                 io_in_r_bypass_regNext_19_2_load_store_22;
  reg                 io_in_r_bypass_regNext_19_2_df_is_ws_22;
  reg                 io_in_r_bypass_regNext_19_2_stall_22;
  reg        [15:0]   io_in_r_bypass_regNext_19_3_data_22;
  reg                 io_in_r_bypass_regNext_19_3_load_store_22;
  reg                 io_in_r_bypass_regNext_19_3_df_is_ws_22;
  reg                 io_in_r_bypass_regNext_19_3_stall_22;
  reg        [15:0]   io_in_r_bypass_regNext_20_0_data_22;
  reg                 io_in_r_bypass_regNext_20_0_load_store_22;
  reg                 io_in_r_bypass_regNext_20_0_df_is_ws_22;
  reg                 io_in_r_bypass_regNext_20_0_stall_22;
  reg        [15:0]   io_in_r_bypass_regNext_20_1_data_22;
  reg                 io_in_r_bypass_regNext_20_1_load_store_22;
  reg                 io_in_r_bypass_regNext_20_1_df_is_ws_22;
  reg                 io_in_r_bypass_regNext_20_1_stall_22;
  reg        [15:0]   io_in_r_bypass_regNext_20_2_data_22;
  reg                 io_in_r_bypass_regNext_20_2_load_store_22;
  reg                 io_in_r_bypass_regNext_20_2_df_is_ws_22;
  reg                 io_in_r_bypass_regNext_20_2_stall_22;
  reg        [15:0]   io_in_r_bypass_regNext_20_3_data_22;
  reg                 io_in_r_bypass_regNext_20_3_load_store_22;
  reg                 io_in_r_bypass_regNext_20_3_df_is_ws_22;
  reg                 io_in_r_bypass_regNext_20_3_stall_22;
  reg        [15:0]   io_in_r_bypass_regNext_21_0_data_22;
  reg                 io_in_r_bypass_regNext_21_0_load_store_22;
  reg                 io_in_r_bypass_regNext_21_0_df_is_ws_22;
  reg                 io_in_r_bypass_regNext_21_0_stall_22;
  reg        [15:0]   io_in_r_bypass_regNext_21_1_data_22;
  reg                 io_in_r_bypass_regNext_21_1_load_store_22;
  reg                 io_in_r_bypass_regNext_21_1_df_is_ws_22;
  reg                 io_in_r_bypass_regNext_21_1_stall_22;
  reg        [15:0]   io_in_r_bypass_regNext_21_2_data_22;
  reg                 io_in_r_bypass_regNext_21_2_load_store_22;
  reg                 io_in_r_bypass_regNext_21_2_df_is_ws_22;
  reg                 io_in_r_bypass_regNext_21_2_stall_22;
  reg        [15:0]   io_in_r_bypass_regNext_21_3_data_22;
  reg                 io_in_r_bypass_regNext_21_3_load_store_22;
  reg                 io_in_r_bypass_regNext_21_3_df_is_ws_22;
  reg                 io_in_r_bypass_regNext_21_3_stall_22;
  reg        [15:0]   io_in_r_bypass_regNext_22_0_data_22;
  reg                 io_in_r_bypass_regNext_22_0_load_store_22;
  reg                 io_in_r_bypass_regNext_22_0_df_is_ws_22;
  reg                 io_in_r_bypass_regNext_22_0_stall_22;
  reg        [15:0]   io_in_r_bypass_regNext_22_1_data_22;
  reg                 io_in_r_bypass_regNext_22_1_load_store_22;
  reg                 io_in_r_bypass_regNext_22_1_df_is_ws_22;
  reg                 io_in_r_bypass_regNext_22_1_stall_22;
  reg        [15:0]   io_in_r_bypass_regNext_22_2_data_22;
  reg                 io_in_r_bypass_regNext_22_2_load_store_22;
  reg                 io_in_r_bypass_regNext_22_2_df_is_ws_22;
  reg                 io_in_r_bypass_regNext_22_2_stall_22;
  reg        [15:0]   io_in_r_bypass_regNext_22_3_data_22;
  reg                 io_in_r_bypass_regNext_22_3_load_store_22;
  reg                 io_in_r_bypass_regNext_22_3_df_is_ws_22;
  reg                 io_in_r_bypass_regNext_22_3_stall_22;
  reg        [15:0]   io_in_r_bypass_regNext_23_0_data_22;
  reg                 io_in_r_bypass_regNext_23_0_load_store_22;
  reg                 io_in_r_bypass_regNext_23_0_df_is_ws_22;
  reg                 io_in_r_bypass_regNext_23_0_stall_22;
  reg        [15:0]   io_in_r_bypass_regNext_23_1_data_22;
  reg                 io_in_r_bypass_regNext_23_1_load_store_22;
  reg                 io_in_r_bypass_regNext_23_1_df_is_ws_22;
  reg                 io_in_r_bypass_regNext_23_1_stall_22;
  reg        [15:0]   io_in_r_bypass_regNext_23_2_data_22;
  reg                 io_in_r_bypass_regNext_23_2_load_store_22;
  reg                 io_in_r_bypass_regNext_23_2_df_is_ws_22;
  reg                 io_in_r_bypass_regNext_23_2_stall_22;
  reg        [15:0]   io_in_r_bypass_regNext_23_3_data_22;
  reg                 io_in_r_bypass_regNext_23_3_load_store_22;
  reg                 io_in_r_bypass_regNext_23_3_df_is_ws_22;
  reg                 io_in_r_bypass_regNext_23_3_stall_22;
  reg        [15:0]   io_in_r_bypass_regNext_24_0_data_22;
  reg                 io_in_r_bypass_regNext_24_0_load_store_22;
  reg                 io_in_r_bypass_regNext_24_0_df_is_ws_22;
  reg                 io_in_r_bypass_regNext_24_0_stall_22;
  reg        [15:0]   io_in_r_bypass_regNext_24_1_data_22;
  reg                 io_in_r_bypass_regNext_24_1_load_store_22;
  reg                 io_in_r_bypass_regNext_24_1_df_is_ws_22;
  reg                 io_in_r_bypass_regNext_24_1_stall_22;
  reg        [15:0]   io_in_r_bypass_regNext_24_2_data_22;
  reg                 io_in_r_bypass_regNext_24_2_load_store_22;
  reg                 io_in_r_bypass_regNext_24_2_df_is_ws_22;
  reg                 io_in_r_bypass_regNext_24_2_stall_22;
  reg        [15:0]   io_in_r_bypass_regNext_24_3_data_22;
  reg                 io_in_r_bypass_regNext_24_3_load_store_22;
  reg                 io_in_r_bypass_regNext_24_3_df_is_ws_22;
  reg                 io_in_r_bypass_regNext_24_3_stall_22;
  reg        [15:0]   io_in_r_bypass_regNext_25_0_data_22;
  reg                 io_in_r_bypass_regNext_25_0_load_store_22;
  reg                 io_in_r_bypass_regNext_25_0_df_is_ws_22;
  reg                 io_in_r_bypass_regNext_25_0_stall_22;
  reg        [15:0]   io_in_r_bypass_regNext_25_1_data_22;
  reg                 io_in_r_bypass_regNext_25_1_load_store_22;
  reg                 io_in_r_bypass_regNext_25_1_df_is_ws_22;
  reg                 io_in_r_bypass_regNext_25_1_stall_22;
  reg        [15:0]   io_in_r_bypass_regNext_25_2_data_22;
  reg                 io_in_r_bypass_regNext_25_2_load_store_22;
  reg                 io_in_r_bypass_regNext_25_2_df_is_ws_22;
  reg                 io_in_r_bypass_regNext_25_2_stall_22;
  reg        [15:0]   io_in_r_bypass_regNext_25_3_data_22;
  reg                 io_in_r_bypass_regNext_25_3_load_store_22;
  reg                 io_in_r_bypass_regNext_25_3_df_is_ws_22;
  reg                 io_in_r_bypass_regNext_25_3_stall_22;
  reg        [15:0]   io_in_r_bypass_regNext_26_0_data_22;
  reg                 io_in_r_bypass_regNext_26_0_load_store_22;
  reg                 io_in_r_bypass_regNext_26_0_df_is_ws_22;
  reg                 io_in_r_bypass_regNext_26_0_stall_22;
  reg        [15:0]   io_in_r_bypass_regNext_26_1_data_22;
  reg                 io_in_r_bypass_regNext_26_1_load_store_22;
  reg                 io_in_r_bypass_regNext_26_1_df_is_ws_22;
  reg                 io_in_r_bypass_regNext_26_1_stall_22;
  reg        [15:0]   io_in_r_bypass_regNext_26_2_data_22;
  reg                 io_in_r_bypass_regNext_26_2_load_store_22;
  reg                 io_in_r_bypass_regNext_26_2_df_is_ws_22;
  reg                 io_in_r_bypass_regNext_26_2_stall_22;
  reg        [15:0]   io_in_r_bypass_regNext_26_3_data_22;
  reg                 io_in_r_bypass_regNext_26_3_load_store_22;
  reg                 io_in_r_bypass_regNext_26_3_df_is_ws_22;
  reg                 io_in_r_bypass_regNext_26_3_stall_22;
  reg        [15:0]   io_in_r_bypass_regNext_27_0_data_22;
  reg                 io_in_r_bypass_regNext_27_0_load_store_22;
  reg                 io_in_r_bypass_regNext_27_0_df_is_ws_22;
  reg                 io_in_r_bypass_regNext_27_0_stall_22;
  reg        [15:0]   io_in_r_bypass_regNext_27_1_data_22;
  reg                 io_in_r_bypass_regNext_27_1_load_store_22;
  reg                 io_in_r_bypass_regNext_27_1_df_is_ws_22;
  reg                 io_in_r_bypass_regNext_27_1_stall_22;
  reg        [15:0]   io_in_r_bypass_regNext_27_2_data_22;
  reg                 io_in_r_bypass_regNext_27_2_load_store_22;
  reg                 io_in_r_bypass_regNext_27_2_df_is_ws_22;
  reg                 io_in_r_bypass_regNext_27_2_stall_22;
  reg        [15:0]   io_in_r_bypass_regNext_27_3_data_22;
  reg                 io_in_r_bypass_regNext_27_3_load_store_22;
  reg                 io_in_r_bypass_regNext_27_3_df_is_ws_22;
  reg                 io_in_r_bypass_regNext_27_3_stall_22;
  reg        [15:0]   io_in_r_bypass_regNext_28_0_data_22;
  reg                 io_in_r_bypass_regNext_28_0_load_store_22;
  reg                 io_in_r_bypass_regNext_28_0_df_is_ws_22;
  reg                 io_in_r_bypass_regNext_28_0_stall_22;
  reg        [15:0]   io_in_r_bypass_regNext_28_1_data_22;
  reg                 io_in_r_bypass_regNext_28_1_load_store_22;
  reg                 io_in_r_bypass_regNext_28_1_df_is_ws_22;
  reg                 io_in_r_bypass_regNext_28_1_stall_22;
  reg        [15:0]   io_in_r_bypass_regNext_28_2_data_22;
  reg                 io_in_r_bypass_regNext_28_2_load_store_22;
  reg                 io_in_r_bypass_regNext_28_2_df_is_ws_22;
  reg                 io_in_r_bypass_regNext_28_2_stall_22;
  reg        [15:0]   io_in_r_bypass_regNext_28_3_data_22;
  reg                 io_in_r_bypass_regNext_28_3_load_store_22;
  reg                 io_in_r_bypass_regNext_28_3_df_is_ws_22;
  reg                 io_in_r_bypass_regNext_28_3_stall_22;
  reg        [15:0]   io_in_r_bypass_regNext_29_0_data_22;
  reg                 io_in_r_bypass_regNext_29_0_load_store_22;
  reg                 io_in_r_bypass_regNext_29_0_df_is_ws_22;
  reg                 io_in_r_bypass_regNext_29_0_stall_22;
  reg        [15:0]   io_in_r_bypass_regNext_29_1_data_22;
  reg                 io_in_r_bypass_regNext_29_1_load_store_22;
  reg                 io_in_r_bypass_regNext_29_1_df_is_ws_22;
  reg                 io_in_r_bypass_regNext_29_1_stall_22;
  reg        [15:0]   io_in_r_bypass_regNext_29_2_data_22;
  reg                 io_in_r_bypass_regNext_29_2_load_store_22;
  reg                 io_in_r_bypass_regNext_29_2_df_is_ws_22;
  reg                 io_in_r_bypass_regNext_29_2_stall_22;
  reg        [15:0]   io_in_r_bypass_regNext_29_3_data_22;
  reg                 io_in_r_bypass_regNext_29_3_load_store_22;
  reg                 io_in_r_bypass_regNext_29_3_df_is_ws_22;
  reg                 io_in_r_bypass_regNext_29_3_stall_22;
  reg        [15:0]   io_in_r_bypass_regNext_30_0_data_22;
  reg                 io_in_r_bypass_regNext_30_0_load_store_22;
  reg                 io_in_r_bypass_regNext_30_0_df_is_ws_22;
  reg                 io_in_r_bypass_regNext_30_0_stall_22;
  reg        [15:0]   io_in_r_bypass_regNext_30_1_data_22;
  reg                 io_in_r_bypass_regNext_30_1_load_store_22;
  reg                 io_in_r_bypass_regNext_30_1_df_is_ws_22;
  reg                 io_in_r_bypass_regNext_30_1_stall_22;
  reg        [15:0]   io_in_r_bypass_regNext_30_2_data_22;
  reg                 io_in_r_bypass_regNext_30_2_load_store_22;
  reg                 io_in_r_bypass_regNext_30_2_df_is_ws_22;
  reg                 io_in_r_bypass_regNext_30_2_stall_22;
  reg        [15:0]   io_in_r_bypass_regNext_30_3_data_22;
  reg                 io_in_r_bypass_regNext_30_3_load_store_22;
  reg                 io_in_r_bypass_regNext_30_3_df_is_ws_22;
  reg                 io_in_r_bypass_regNext_30_3_stall_22;
  reg        [15:0]   io_in_r_bypass_regNext_31_0_data_22;
  reg                 io_in_r_bypass_regNext_31_0_load_store_22;
  reg                 io_in_r_bypass_regNext_31_0_df_is_ws_22;
  reg                 io_in_r_bypass_regNext_31_0_stall_22;
  reg        [15:0]   io_in_r_bypass_regNext_31_1_data_22;
  reg                 io_in_r_bypass_regNext_31_1_load_store_22;
  reg                 io_in_r_bypass_regNext_31_1_df_is_ws_22;
  reg                 io_in_r_bypass_regNext_31_1_stall_22;
  reg        [15:0]   io_in_r_bypass_regNext_31_2_data_22;
  reg                 io_in_r_bypass_regNext_31_2_load_store_22;
  reg                 io_in_r_bypass_regNext_31_2_df_is_ws_22;
  reg                 io_in_r_bypass_regNext_31_2_stall_22;
  reg        [15:0]   io_in_r_bypass_regNext_31_3_data_22;
  reg                 io_in_r_bypass_regNext_31_3_load_store_22;
  reg                 io_in_r_bypass_regNext_31_3_df_is_ws_22;
  reg                 io_in_r_bypass_regNext_31_3_stall_22;
  reg        [15:0]   io_in_r_bypass_regNext_0_0_data_23;
  reg                 io_in_r_bypass_regNext_0_0_load_store_23;
  reg                 io_in_r_bypass_regNext_0_0_df_is_ws_23;
  reg                 io_in_r_bypass_regNext_0_0_stall_23;
  reg        [15:0]   io_in_r_bypass_regNext_0_1_data_23;
  reg                 io_in_r_bypass_regNext_0_1_load_store_23;
  reg                 io_in_r_bypass_regNext_0_1_df_is_ws_23;
  reg                 io_in_r_bypass_regNext_0_1_stall_23;
  reg        [15:0]   io_in_r_bypass_regNext_0_2_data_23;
  reg                 io_in_r_bypass_regNext_0_2_load_store_23;
  reg                 io_in_r_bypass_regNext_0_2_df_is_ws_23;
  reg                 io_in_r_bypass_regNext_0_2_stall_23;
  reg        [15:0]   io_in_r_bypass_regNext_0_3_data_23;
  reg                 io_in_r_bypass_regNext_0_3_load_store_23;
  reg                 io_in_r_bypass_regNext_0_3_df_is_ws_23;
  reg                 io_in_r_bypass_regNext_0_3_stall_23;
  reg        [15:0]   io_in_r_bypass_regNext_1_0_data_23;
  reg                 io_in_r_bypass_regNext_1_0_load_store_23;
  reg                 io_in_r_bypass_regNext_1_0_df_is_ws_23;
  reg                 io_in_r_bypass_regNext_1_0_stall_23;
  reg        [15:0]   io_in_r_bypass_regNext_1_1_data_23;
  reg                 io_in_r_bypass_regNext_1_1_load_store_23;
  reg                 io_in_r_bypass_regNext_1_1_df_is_ws_23;
  reg                 io_in_r_bypass_regNext_1_1_stall_23;
  reg        [15:0]   io_in_r_bypass_regNext_1_2_data_23;
  reg                 io_in_r_bypass_regNext_1_2_load_store_23;
  reg                 io_in_r_bypass_regNext_1_2_df_is_ws_23;
  reg                 io_in_r_bypass_regNext_1_2_stall_23;
  reg        [15:0]   io_in_r_bypass_regNext_1_3_data_23;
  reg                 io_in_r_bypass_regNext_1_3_load_store_23;
  reg                 io_in_r_bypass_regNext_1_3_df_is_ws_23;
  reg                 io_in_r_bypass_regNext_1_3_stall_23;
  reg        [15:0]   io_in_r_bypass_regNext_2_0_data_23;
  reg                 io_in_r_bypass_regNext_2_0_load_store_23;
  reg                 io_in_r_bypass_regNext_2_0_df_is_ws_23;
  reg                 io_in_r_bypass_regNext_2_0_stall_23;
  reg        [15:0]   io_in_r_bypass_regNext_2_1_data_23;
  reg                 io_in_r_bypass_regNext_2_1_load_store_23;
  reg                 io_in_r_bypass_regNext_2_1_df_is_ws_23;
  reg                 io_in_r_bypass_regNext_2_1_stall_23;
  reg        [15:0]   io_in_r_bypass_regNext_2_2_data_23;
  reg                 io_in_r_bypass_regNext_2_2_load_store_23;
  reg                 io_in_r_bypass_regNext_2_2_df_is_ws_23;
  reg                 io_in_r_bypass_regNext_2_2_stall_23;
  reg        [15:0]   io_in_r_bypass_regNext_2_3_data_23;
  reg                 io_in_r_bypass_regNext_2_3_load_store_23;
  reg                 io_in_r_bypass_regNext_2_3_df_is_ws_23;
  reg                 io_in_r_bypass_regNext_2_3_stall_23;
  reg        [15:0]   io_in_r_bypass_regNext_3_0_data_23;
  reg                 io_in_r_bypass_regNext_3_0_load_store_23;
  reg                 io_in_r_bypass_regNext_3_0_df_is_ws_23;
  reg                 io_in_r_bypass_regNext_3_0_stall_23;
  reg        [15:0]   io_in_r_bypass_regNext_3_1_data_23;
  reg                 io_in_r_bypass_regNext_3_1_load_store_23;
  reg                 io_in_r_bypass_regNext_3_1_df_is_ws_23;
  reg                 io_in_r_bypass_regNext_3_1_stall_23;
  reg        [15:0]   io_in_r_bypass_regNext_3_2_data_23;
  reg                 io_in_r_bypass_regNext_3_2_load_store_23;
  reg                 io_in_r_bypass_regNext_3_2_df_is_ws_23;
  reg                 io_in_r_bypass_regNext_3_2_stall_23;
  reg        [15:0]   io_in_r_bypass_regNext_3_3_data_23;
  reg                 io_in_r_bypass_regNext_3_3_load_store_23;
  reg                 io_in_r_bypass_regNext_3_3_df_is_ws_23;
  reg                 io_in_r_bypass_regNext_3_3_stall_23;
  reg        [15:0]   io_in_r_bypass_regNext_4_0_data_23;
  reg                 io_in_r_bypass_regNext_4_0_load_store_23;
  reg                 io_in_r_bypass_regNext_4_0_df_is_ws_23;
  reg                 io_in_r_bypass_regNext_4_0_stall_23;
  reg        [15:0]   io_in_r_bypass_regNext_4_1_data_23;
  reg                 io_in_r_bypass_regNext_4_1_load_store_23;
  reg                 io_in_r_bypass_regNext_4_1_df_is_ws_23;
  reg                 io_in_r_bypass_regNext_4_1_stall_23;
  reg        [15:0]   io_in_r_bypass_regNext_4_2_data_23;
  reg                 io_in_r_bypass_regNext_4_2_load_store_23;
  reg                 io_in_r_bypass_regNext_4_2_df_is_ws_23;
  reg                 io_in_r_bypass_regNext_4_2_stall_23;
  reg        [15:0]   io_in_r_bypass_regNext_4_3_data_23;
  reg                 io_in_r_bypass_regNext_4_3_load_store_23;
  reg                 io_in_r_bypass_regNext_4_3_df_is_ws_23;
  reg                 io_in_r_bypass_regNext_4_3_stall_23;
  reg        [15:0]   io_in_r_bypass_regNext_5_0_data_23;
  reg                 io_in_r_bypass_regNext_5_0_load_store_23;
  reg                 io_in_r_bypass_regNext_5_0_df_is_ws_23;
  reg                 io_in_r_bypass_regNext_5_0_stall_23;
  reg        [15:0]   io_in_r_bypass_regNext_5_1_data_23;
  reg                 io_in_r_bypass_regNext_5_1_load_store_23;
  reg                 io_in_r_bypass_regNext_5_1_df_is_ws_23;
  reg                 io_in_r_bypass_regNext_5_1_stall_23;
  reg        [15:0]   io_in_r_bypass_regNext_5_2_data_23;
  reg                 io_in_r_bypass_regNext_5_2_load_store_23;
  reg                 io_in_r_bypass_regNext_5_2_df_is_ws_23;
  reg                 io_in_r_bypass_regNext_5_2_stall_23;
  reg        [15:0]   io_in_r_bypass_regNext_5_3_data_23;
  reg                 io_in_r_bypass_regNext_5_3_load_store_23;
  reg                 io_in_r_bypass_regNext_5_3_df_is_ws_23;
  reg                 io_in_r_bypass_regNext_5_3_stall_23;
  reg        [15:0]   io_in_r_bypass_regNext_6_0_data_23;
  reg                 io_in_r_bypass_regNext_6_0_load_store_23;
  reg                 io_in_r_bypass_regNext_6_0_df_is_ws_23;
  reg                 io_in_r_bypass_regNext_6_0_stall_23;
  reg        [15:0]   io_in_r_bypass_regNext_6_1_data_23;
  reg                 io_in_r_bypass_regNext_6_1_load_store_23;
  reg                 io_in_r_bypass_regNext_6_1_df_is_ws_23;
  reg                 io_in_r_bypass_regNext_6_1_stall_23;
  reg        [15:0]   io_in_r_bypass_regNext_6_2_data_23;
  reg                 io_in_r_bypass_regNext_6_2_load_store_23;
  reg                 io_in_r_bypass_regNext_6_2_df_is_ws_23;
  reg                 io_in_r_bypass_regNext_6_2_stall_23;
  reg        [15:0]   io_in_r_bypass_regNext_6_3_data_23;
  reg                 io_in_r_bypass_regNext_6_3_load_store_23;
  reg                 io_in_r_bypass_regNext_6_3_df_is_ws_23;
  reg                 io_in_r_bypass_regNext_6_3_stall_23;
  reg        [15:0]   io_in_r_bypass_regNext_7_0_data_23;
  reg                 io_in_r_bypass_regNext_7_0_load_store_23;
  reg                 io_in_r_bypass_regNext_7_0_df_is_ws_23;
  reg                 io_in_r_bypass_regNext_7_0_stall_23;
  reg        [15:0]   io_in_r_bypass_regNext_7_1_data_23;
  reg                 io_in_r_bypass_regNext_7_1_load_store_23;
  reg                 io_in_r_bypass_regNext_7_1_df_is_ws_23;
  reg                 io_in_r_bypass_regNext_7_1_stall_23;
  reg        [15:0]   io_in_r_bypass_regNext_7_2_data_23;
  reg                 io_in_r_bypass_regNext_7_2_load_store_23;
  reg                 io_in_r_bypass_regNext_7_2_df_is_ws_23;
  reg                 io_in_r_bypass_regNext_7_2_stall_23;
  reg        [15:0]   io_in_r_bypass_regNext_7_3_data_23;
  reg                 io_in_r_bypass_regNext_7_3_load_store_23;
  reg                 io_in_r_bypass_regNext_7_3_df_is_ws_23;
  reg                 io_in_r_bypass_regNext_7_3_stall_23;
  reg        [15:0]   io_in_r_bypass_regNext_8_0_data_23;
  reg                 io_in_r_bypass_regNext_8_0_load_store_23;
  reg                 io_in_r_bypass_regNext_8_0_df_is_ws_23;
  reg                 io_in_r_bypass_regNext_8_0_stall_23;
  reg        [15:0]   io_in_r_bypass_regNext_8_1_data_23;
  reg                 io_in_r_bypass_regNext_8_1_load_store_23;
  reg                 io_in_r_bypass_regNext_8_1_df_is_ws_23;
  reg                 io_in_r_bypass_regNext_8_1_stall_23;
  reg        [15:0]   io_in_r_bypass_regNext_8_2_data_23;
  reg                 io_in_r_bypass_regNext_8_2_load_store_23;
  reg                 io_in_r_bypass_regNext_8_2_df_is_ws_23;
  reg                 io_in_r_bypass_regNext_8_2_stall_23;
  reg        [15:0]   io_in_r_bypass_regNext_8_3_data_23;
  reg                 io_in_r_bypass_regNext_8_3_load_store_23;
  reg                 io_in_r_bypass_regNext_8_3_df_is_ws_23;
  reg                 io_in_r_bypass_regNext_8_3_stall_23;
  reg        [15:0]   io_in_r_bypass_regNext_9_0_data_23;
  reg                 io_in_r_bypass_regNext_9_0_load_store_23;
  reg                 io_in_r_bypass_regNext_9_0_df_is_ws_23;
  reg                 io_in_r_bypass_regNext_9_0_stall_23;
  reg        [15:0]   io_in_r_bypass_regNext_9_1_data_23;
  reg                 io_in_r_bypass_regNext_9_1_load_store_23;
  reg                 io_in_r_bypass_regNext_9_1_df_is_ws_23;
  reg                 io_in_r_bypass_regNext_9_1_stall_23;
  reg        [15:0]   io_in_r_bypass_regNext_9_2_data_23;
  reg                 io_in_r_bypass_regNext_9_2_load_store_23;
  reg                 io_in_r_bypass_regNext_9_2_df_is_ws_23;
  reg                 io_in_r_bypass_regNext_9_2_stall_23;
  reg        [15:0]   io_in_r_bypass_regNext_9_3_data_23;
  reg                 io_in_r_bypass_regNext_9_3_load_store_23;
  reg                 io_in_r_bypass_regNext_9_3_df_is_ws_23;
  reg                 io_in_r_bypass_regNext_9_3_stall_23;
  reg        [15:0]   io_in_r_bypass_regNext_10_0_data_23;
  reg                 io_in_r_bypass_regNext_10_0_load_store_23;
  reg                 io_in_r_bypass_regNext_10_0_df_is_ws_23;
  reg                 io_in_r_bypass_regNext_10_0_stall_23;
  reg        [15:0]   io_in_r_bypass_regNext_10_1_data_23;
  reg                 io_in_r_bypass_regNext_10_1_load_store_23;
  reg                 io_in_r_bypass_regNext_10_1_df_is_ws_23;
  reg                 io_in_r_bypass_regNext_10_1_stall_23;
  reg        [15:0]   io_in_r_bypass_regNext_10_2_data_23;
  reg                 io_in_r_bypass_regNext_10_2_load_store_23;
  reg                 io_in_r_bypass_regNext_10_2_df_is_ws_23;
  reg                 io_in_r_bypass_regNext_10_2_stall_23;
  reg        [15:0]   io_in_r_bypass_regNext_10_3_data_23;
  reg                 io_in_r_bypass_regNext_10_3_load_store_23;
  reg                 io_in_r_bypass_regNext_10_3_df_is_ws_23;
  reg                 io_in_r_bypass_regNext_10_3_stall_23;
  reg        [15:0]   io_in_r_bypass_regNext_11_0_data_23;
  reg                 io_in_r_bypass_regNext_11_0_load_store_23;
  reg                 io_in_r_bypass_regNext_11_0_df_is_ws_23;
  reg                 io_in_r_bypass_regNext_11_0_stall_23;
  reg        [15:0]   io_in_r_bypass_regNext_11_1_data_23;
  reg                 io_in_r_bypass_regNext_11_1_load_store_23;
  reg                 io_in_r_bypass_regNext_11_1_df_is_ws_23;
  reg                 io_in_r_bypass_regNext_11_1_stall_23;
  reg        [15:0]   io_in_r_bypass_regNext_11_2_data_23;
  reg                 io_in_r_bypass_regNext_11_2_load_store_23;
  reg                 io_in_r_bypass_regNext_11_2_df_is_ws_23;
  reg                 io_in_r_bypass_regNext_11_2_stall_23;
  reg        [15:0]   io_in_r_bypass_regNext_11_3_data_23;
  reg                 io_in_r_bypass_regNext_11_3_load_store_23;
  reg                 io_in_r_bypass_regNext_11_3_df_is_ws_23;
  reg                 io_in_r_bypass_regNext_11_3_stall_23;
  reg        [15:0]   io_in_r_bypass_regNext_12_0_data_23;
  reg                 io_in_r_bypass_regNext_12_0_load_store_23;
  reg                 io_in_r_bypass_regNext_12_0_df_is_ws_23;
  reg                 io_in_r_bypass_regNext_12_0_stall_23;
  reg        [15:0]   io_in_r_bypass_regNext_12_1_data_23;
  reg                 io_in_r_bypass_regNext_12_1_load_store_23;
  reg                 io_in_r_bypass_regNext_12_1_df_is_ws_23;
  reg                 io_in_r_bypass_regNext_12_1_stall_23;
  reg        [15:0]   io_in_r_bypass_regNext_12_2_data_23;
  reg                 io_in_r_bypass_regNext_12_2_load_store_23;
  reg                 io_in_r_bypass_regNext_12_2_df_is_ws_23;
  reg                 io_in_r_bypass_regNext_12_2_stall_23;
  reg        [15:0]   io_in_r_bypass_regNext_12_3_data_23;
  reg                 io_in_r_bypass_regNext_12_3_load_store_23;
  reg                 io_in_r_bypass_regNext_12_3_df_is_ws_23;
  reg                 io_in_r_bypass_regNext_12_3_stall_23;
  reg        [15:0]   io_in_r_bypass_regNext_13_0_data_23;
  reg                 io_in_r_bypass_regNext_13_0_load_store_23;
  reg                 io_in_r_bypass_regNext_13_0_df_is_ws_23;
  reg                 io_in_r_bypass_regNext_13_0_stall_23;
  reg        [15:0]   io_in_r_bypass_regNext_13_1_data_23;
  reg                 io_in_r_bypass_regNext_13_1_load_store_23;
  reg                 io_in_r_bypass_regNext_13_1_df_is_ws_23;
  reg                 io_in_r_bypass_regNext_13_1_stall_23;
  reg        [15:0]   io_in_r_bypass_regNext_13_2_data_23;
  reg                 io_in_r_bypass_regNext_13_2_load_store_23;
  reg                 io_in_r_bypass_regNext_13_2_df_is_ws_23;
  reg                 io_in_r_bypass_regNext_13_2_stall_23;
  reg        [15:0]   io_in_r_bypass_regNext_13_3_data_23;
  reg                 io_in_r_bypass_regNext_13_3_load_store_23;
  reg                 io_in_r_bypass_regNext_13_3_df_is_ws_23;
  reg                 io_in_r_bypass_regNext_13_3_stall_23;
  reg        [15:0]   io_in_r_bypass_regNext_14_0_data_23;
  reg                 io_in_r_bypass_regNext_14_0_load_store_23;
  reg                 io_in_r_bypass_regNext_14_0_df_is_ws_23;
  reg                 io_in_r_bypass_regNext_14_0_stall_23;
  reg        [15:0]   io_in_r_bypass_regNext_14_1_data_23;
  reg                 io_in_r_bypass_regNext_14_1_load_store_23;
  reg                 io_in_r_bypass_regNext_14_1_df_is_ws_23;
  reg                 io_in_r_bypass_regNext_14_1_stall_23;
  reg        [15:0]   io_in_r_bypass_regNext_14_2_data_23;
  reg                 io_in_r_bypass_regNext_14_2_load_store_23;
  reg                 io_in_r_bypass_regNext_14_2_df_is_ws_23;
  reg                 io_in_r_bypass_regNext_14_2_stall_23;
  reg        [15:0]   io_in_r_bypass_regNext_14_3_data_23;
  reg                 io_in_r_bypass_regNext_14_3_load_store_23;
  reg                 io_in_r_bypass_regNext_14_3_df_is_ws_23;
  reg                 io_in_r_bypass_regNext_14_3_stall_23;
  reg        [15:0]   io_in_r_bypass_regNext_15_0_data_23;
  reg                 io_in_r_bypass_regNext_15_0_load_store_23;
  reg                 io_in_r_bypass_regNext_15_0_df_is_ws_23;
  reg                 io_in_r_bypass_regNext_15_0_stall_23;
  reg        [15:0]   io_in_r_bypass_regNext_15_1_data_23;
  reg                 io_in_r_bypass_regNext_15_1_load_store_23;
  reg                 io_in_r_bypass_regNext_15_1_df_is_ws_23;
  reg                 io_in_r_bypass_regNext_15_1_stall_23;
  reg        [15:0]   io_in_r_bypass_regNext_15_2_data_23;
  reg                 io_in_r_bypass_regNext_15_2_load_store_23;
  reg                 io_in_r_bypass_regNext_15_2_df_is_ws_23;
  reg                 io_in_r_bypass_regNext_15_2_stall_23;
  reg        [15:0]   io_in_r_bypass_regNext_15_3_data_23;
  reg                 io_in_r_bypass_regNext_15_3_load_store_23;
  reg                 io_in_r_bypass_regNext_15_3_df_is_ws_23;
  reg                 io_in_r_bypass_regNext_15_3_stall_23;
  reg        [15:0]   io_in_r_bypass_regNext_16_0_data_23;
  reg                 io_in_r_bypass_regNext_16_0_load_store_23;
  reg                 io_in_r_bypass_regNext_16_0_df_is_ws_23;
  reg                 io_in_r_bypass_regNext_16_0_stall_23;
  reg        [15:0]   io_in_r_bypass_regNext_16_1_data_23;
  reg                 io_in_r_bypass_regNext_16_1_load_store_23;
  reg                 io_in_r_bypass_regNext_16_1_df_is_ws_23;
  reg                 io_in_r_bypass_regNext_16_1_stall_23;
  reg        [15:0]   io_in_r_bypass_regNext_16_2_data_23;
  reg                 io_in_r_bypass_regNext_16_2_load_store_23;
  reg                 io_in_r_bypass_regNext_16_2_df_is_ws_23;
  reg                 io_in_r_bypass_regNext_16_2_stall_23;
  reg        [15:0]   io_in_r_bypass_regNext_16_3_data_23;
  reg                 io_in_r_bypass_regNext_16_3_load_store_23;
  reg                 io_in_r_bypass_regNext_16_3_df_is_ws_23;
  reg                 io_in_r_bypass_regNext_16_3_stall_23;
  reg        [15:0]   io_in_r_bypass_regNext_17_0_data_23;
  reg                 io_in_r_bypass_regNext_17_0_load_store_23;
  reg                 io_in_r_bypass_regNext_17_0_df_is_ws_23;
  reg                 io_in_r_bypass_regNext_17_0_stall_23;
  reg        [15:0]   io_in_r_bypass_regNext_17_1_data_23;
  reg                 io_in_r_bypass_regNext_17_1_load_store_23;
  reg                 io_in_r_bypass_regNext_17_1_df_is_ws_23;
  reg                 io_in_r_bypass_regNext_17_1_stall_23;
  reg        [15:0]   io_in_r_bypass_regNext_17_2_data_23;
  reg                 io_in_r_bypass_regNext_17_2_load_store_23;
  reg                 io_in_r_bypass_regNext_17_2_df_is_ws_23;
  reg                 io_in_r_bypass_regNext_17_2_stall_23;
  reg        [15:0]   io_in_r_bypass_regNext_17_3_data_23;
  reg                 io_in_r_bypass_regNext_17_3_load_store_23;
  reg                 io_in_r_bypass_regNext_17_3_df_is_ws_23;
  reg                 io_in_r_bypass_regNext_17_3_stall_23;
  reg        [15:0]   io_in_r_bypass_regNext_18_0_data_23;
  reg                 io_in_r_bypass_regNext_18_0_load_store_23;
  reg                 io_in_r_bypass_regNext_18_0_df_is_ws_23;
  reg                 io_in_r_bypass_regNext_18_0_stall_23;
  reg        [15:0]   io_in_r_bypass_regNext_18_1_data_23;
  reg                 io_in_r_bypass_regNext_18_1_load_store_23;
  reg                 io_in_r_bypass_regNext_18_1_df_is_ws_23;
  reg                 io_in_r_bypass_regNext_18_1_stall_23;
  reg        [15:0]   io_in_r_bypass_regNext_18_2_data_23;
  reg                 io_in_r_bypass_regNext_18_2_load_store_23;
  reg                 io_in_r_bypass_regNext_18_2_df_is_ws_23;
  reg                 io_in_r_bypass_regNext_18_2_stall_23;
  reg        [15:0]   io_in_r_bypass_regNext_18_3_data_23;
  reg                 io_in_r_bypass_regNext_18_3_load_store_23;
  reg                 io_in_r_bypass_regNext_18_3_df_is_ws_23;
  reg                 io_in_r_bypass_regNext_18_3_stall_23;
  reg        [15:0]   io_in_r_bypass_regNext_19_0_data_23;
  reg                 io_in_r_bypass_regNext_19_0_load_store_23;
  reg                 io_in_r_bypass_regNext_19_0_df_is_ws_23;
  reg                 io_in_r_bypass_regNext_19_0_stall_23;
  reg        [15:0]   io_in_r_bypass_regNext_19_1_data_23;
  reg                 io_in_r_bypass_regNext_19_1_load_store_23;
  reg                 io_in_r_bypass_regNext_19_1_df_is_ws_23;
  reg                 io_in_r_bypass_regNext_19_1_stall_23;
  reg        [15:0]   io_in_r_bypass_regNext_19_2_data_23;
  reg                 io_in_r_bypass_regNext_19_2_load_store_23;
  reg                 io_in_r_bypass_regNext_19_2_df_is_ws_23;
  reg                 io_in_r_bypass_regNext_19_2_stall_23;
  reg        [15:0]   io_in_r_bypass_regNext_19_3_data_23;
  reg                 io_in_r_bypass_regNext_19_3_load_store_23;
  reg                 io_in_r_bypass_regNext_19_3_df_is_ws_23;
  reg                 io_in_r_bypass_regNext_19_3_stall_23;
  reg        [15:0]   io_in_r_bypass_regNext_20_0_data_23;
  reg                 io_in_r_bypass_regNext_20_0_load_store_23;
  reg                 io_in_r_bypass_regNext_20_0_df_is_ws_23;
  reg                 io_in_r_bypass_regNext_20_0_stall_23;
  reg        [15:0]   io_in_r_bypass_regNext_20_1_data_23;
  reg                 io_in_r_bypass_regNext_20_1_load_store_23;
  reg                 io_in_r_bypass_regNext_20_1_df_is_ws_23;
  reg                 io_in_r_bypass_regNext_20_1_stall_23;
  reg        [15:0]   io_in_r_bypass_regNext_20_2_data_23;
  reg                 io_in_r_bypass_regNext_20_2_load_store_23;
  reg                 io_in_r_bypass_regNext_20_2_df_is_ws_23;
  reg                 io_in_r_bypass_regNext_20_2_stall_23;
  reg        [15:0]   io_in_r_bypass_regNext_20_3_data_23;
  reg                 io_in_r_bypass_regNext_20_3_load_store_23;
  reg                 io_in_r_bypass_regNext_20_3_df_is_ws_23;
  reg                 io_in_r_bypass_regNext_20_3_stall_23;
  reg        [15:0]   io_in_r_bypass_regNext_21_0_data_23;
  reg                 io_in_r_bypass_regNext_21_0_load_store_23;
  reg                 io_in_r_bypass_regNext_21_0_df_is_ws_23;
  reg                 io_in_r_bypass_regNext_21_0_stall_23;
  reg        [15:0]   io_in_r_bypass_regNext_21_1_data_23;
  reg                 io_in_r_bypass_regNext_21_1_load_store_23;
  reg                 io_in_r_bypass_regNext_21_1_df_is_ws_23;
  reg                 io_in_r_bypass_regNext_21_1_stall_23;
  reg        [15:0]   io_in_r_bypass_regNext_21_2_data_23;
  reg                 io_in_r_bypass_regNext_21_2_load_store_23;
  reg                 io_in_r_bypass_regNext_21_2_df_is_ws_23;
  reg                 io_in_r_bypass_regNext_21_2_stall_23;
  reg        [15:0]   io_in_r_bypass_regNext_21_3_data_23;
  reg                 io_in_r_bypass_regNext_21_3_load_store_23;
  reg                 io_in_r_bypass_regNext_21_3_df_is_ws_23;
  reg                 io_in_r_bypass_regNext_21_3_stall_23;
  reg        [15:0]   io_in_r_bypass_regNext_22_0_data_23;
  reg                 io_in_r_bypass_regNext_22_0_load_store_23;
  reg                 io_in_r_bypass_regNext_22_0_df_is_ws_23;
  reg                 io_in_r_bypass_regNext_22_0_stall_23;
  reg        [15:0]   io_in_r_bypass_regNext_22_1_data_23;
  reg                 io_in_r_bypass_regNext_22_1_load_store_23;
  reg                 io_in_r_bypass_regNext_22_1_df_is_ws_23;
  reg                 io_in_r_bypass_regNext_22_1_stall_23;
  reg        [15:0]   io_in_r_bypass_regNext_22_2_data_23;
  reg                 io_in_r_bypass_regNext_22_2_load_store_23;
  reg                 io_in_r_bypass_regNext_22_2_df_is_ws_23;
  reg                 io_in_r_bypass_regNext_22_2_stall_23;
  reg        [15:0]   io_in_r_bypass_regNext_22_3_data_23;
  reg                 io_in_r_bypass_regNext_22_3_load_store_23;
  reg                 io_in_r_bypass_regNext_22_3_df_is_ws_23;
  reg                 io_in_r_bypass_regNext_22_3_stall_23;
  reg        [15:0]   io_in_r_bypass_regNext_23_0_data_23;
  reg                 io_in_r_bypass_regNext_23_0_load_store_23;
  reg                 io_in_r_bypass_regNext_23_0_df_is_ws_23;
  reg                 io_in_r_bypass_regNext_23_0_stall_23;
  reg        [15:0]   io_in_r_bypass_regNext_23_1_data_23;
  reg                 io_in_r_bypass_regNext_23_1_load_store_23;
  reg                 io_in_r_bypass_regNext_23_1_df_is_ws_23;
  reg                 io_in_r_bypass_regNext_23_1_stall_23;
  reg        [15:0]   io_in_r_bypass_regNext_23_2_data_23;
  reg                 io_in_r_bypass_regNext_23_2_load_store_23;
  reg                 io_in_r_bypass_regNext_23_2_df_is_ws_23;
  reg                 io_in_r_bypass_regNext_23_2_stall_23;
  reg        [15:0]   io_in_r_bypass_regNext_23_3_data_23;
  reg                 io_in_r_bypass_regNext_23_3_load_store_23;
  reg                 io_in_r_bypass_regNext_23_3_df_is_ws_23;
  reg                 io_in_r_bypass_regNext_23_3_stall_23;
  reg        [15:0]   io_in_r_bypass_regNext_24_0_data_23;
  reg                 io_in_r_bypass_regNext_24_0_load_store_23;
  reg                 io_in_r_bypass_regNext_24_0_df_is_ws_23;
  reg                 io_in_r_bypass_regNext_24_0_stall_23;
  reg        [15:0]   io_in_r_bypass_regNext_24_1_data_23;
  reg                 io_in_r_bypass_regNext_24_1_load_store_23;
  reg                 io_in_r_bypass_regNext_24_1_df_is_ws_23;
  reg                 io_in_r_bypass_regNext_24_1_stall_23;
  reg        [15:0]   io_in_r_bypass_regNext_24_2_data_23;
  reg                 io_in_r_bypass_regNext_24_2_load_store_23;
  reg                 io_in_r_bypass_regNext_24_2_df_is_ws_23;
  reg                 io_in_r_bypass_regNext_24_2_stall_23;
  reg        [15:0]   io_in_r_bypass_regNext_24_3_data_23;
  reg                 io_in_r_bypass_regNext_24_3_load_store_23;
  reg                 io_in_r_bypass_regNext_24_3_df_is_ws_23;
  reg                 io_in_r_bypass_regNext_24_3_stall_23;
  reg        [15:0]   io_in_r_bypass_regNext_25_0_data_23;
  reg                 io_in_r_bypass_regNext_25_0_load_store_23;
  reg                 io_in_r_bypass_regNext_25_0_df_is_ws_23;
  reg                 io_in_r_bypass_regNext_25_0_stall_23;
  reg        [15:0]   io_in_r_bypass_regNext_25_1_data_23;
  reg                 io_in_r_bypass_regNext_25_1_load_store_23;
  reg                 io_in_r_bypass_regNext_25_1_df_is_ws_23;
  reg                 io_in_r_bypass_regNext_25_1_stall_23;
  reg        [15:0]   io_in_r_bypass_regNext_25_2_data_23;
  reg                 io_in_r_bypass_regNext_25_2_load_store_23;
  reg                 io_in_r_bypass_regNext_25_2_df_is_ws_23;
  reg                 io_in_r_bypass_regNext_25_2_stall_23;
  reg        [15:0]   io_in_r_bypass_regNext_25_3_data_23;
  reg                 io_in_r_bypass_regNext_25_3_load_store_23;
  reg                 io_in_r_bypass_regNext_25_3_df_is_ws_23;
  reg                 io_in_r_bypass_regNext_25_3_stall_23;
  reg        [15:0]   io_in_r_bypass_regNext_26_0_data_23;
  reg                 io_in_r_bypass_regNext_26_0_load_store_23;
  reg                 io_in_r_bypass_regNext_26_0_df_is_ws_23;
  reg                 io_in_r_bypass_regNext_26_0_stall_23;
  reg        [15:0]   io_in_r_bypass_regNext_26_1_data_23;
  reg                 io_in_r_bypass_regNext_26_1_load_store_23;
  reg                 io_in_r_bypass_regNext_26_1_df_is_ws_23;
  reg                 io_in_r_bypass_regNext_26_1_stall_23;
  reg        [15:0]   io_in_r_bypass_regNext_26_2_data_23;
  reg                 io_in_r_bypass_regNext_26_2_load_store_23;
  reg                 io_in_r_bypass_regNext_26_2_df_is_ws_23;
  reg                 io_in_r_bypass_regNext_26_2_stall_23;
  reg        [15:0]   io_in_r_bypass_regNext_26_3_data_23;
  reg                 io_in_r_bypass_regNext_26_3_load_store_23;
  reg                 io_in_r_bypass_regNext_26_3_df_is_ws_23;
  reg                 io_in_r_bypass_regNext_26_3_stall_23;
  reg        [15:0]   io_in_r_bypass_regNext_27_0_data_23;
  reg                 io_in_r_bypass_regNext_27_0_load_store_23;
  reg                 io_in_r_bypass_regNext_27_0_df_is_ws_23;
  reg                 io_in_r_bypass_regNext_27_0_stall_23;
  reg        [15:0]   io_in_r_bypass_regNext_27_1_data_23;
  reg                 io_in_r_bypass_regNext_27_1_load_store_23;
  reg                 io_in_r_bypass_regNext_27_1_df_is_ws_23;
  reg                 io_in_r_bypass_regNext_27_1_stall_23;
  reg        [15:0]   io_in_r_bypass_regNext_27_2_data_23;
  reg                 io_in_r_bypass_regNext_27_2_load_store_23;
  reg                 io_in_r_bypass_regNext_27_2_df_is_ws_23;
  reg                 io_in_r_bypass_regNext_27_2_stall_23;
  reg        [15:0]   io_in_r_bypass_regNext_27_3_data_23;
  reg                 io_in_r_bypass_regNext_27_3_load_store_23;
  reg                 io_in_r_bypass_regNext_27_3_df_is_ws_23;
  reg                 io_in_r_bypass_regNext_27_3_stall_23;
  reg        [15:0]   io_in_r_bypass_regNext_28_0_data_23;
  reg                 io_in_r_bypass_regNext_28_0_load_store_23;
  reg                 io_in_r_bypass_regNext_28_0_df_is_ws_23;
  reg                 io_in_r_bypass_regNext_28_0_stall_23;
  reg        [15:0]   io_in_r_bypass_regNext_28_1_data_23;
  reg                 io_in_r_bypass_regNext_28_1_load_store_23;
  reg                 io_in_r_bypass_regNext_28_1_df_is_ws_23;
  reg                 io_in_r_bypass_regNext_28_1_stall_23;
  reg        [15:0]   io_in_r_bypass_regNext_28_2_data_23;
  reg                 io_in_r_bypass_regNext_28_2_load_store_23;
  reg                 io_in_r_bypass_regNext_28_2_df_is_ws_23;
  reg                 io_in_r_bypass_regNext_28_2_stall_23;
  reg        [15:0]   io_in_r_bypass_regNext_28_3_data_23;
  reg                 io_in_r_bypass_regNext_28_3_load_store_23;
  reg                 io_in_r_bypass_regNext_28_3_df_is_ws_23;
  reg                 io_in_r_bypass_regNext_28_3_stall_23;
  reg        [15:0]   io_in_r_bypass_regNext_29_0_data_23;
  reg                 io_in_r_bypass_regNext_29_0_load_store_23;
  reg                 io_in_r_bypass_regNext_29_0_df_is_ws_23;
  reg                 io_in_r_bypass_regNext_29_0_stall_23;
  reg        [15:0]   io_in_r_bypass_regNext_29_1_data_23;
  reg                 io_in_r_bypass_regNext_29_1_load_store_23;
  reg                 io_in_r_bypass_regNext_29_1_df_is_ws_23;
  reg                 io_in_r_bypass_regNext_29_1_stall_23;
  reg        [15:0]   io_in_r_bypass_regNext_29_2_data_23;
  reg                 io_in_r_bypass_regNext_29_2_load_store_23;
  reg                 io_in_r_bypass_regNext_29_2_df_is_ws_23;
  reg                 io_in_r_bypass_regNext_29_2_stall_23;
  reg        [15:0]   io_in_r_bypass_regNext_29_3_data_23;
  reg                 io_in_r_bypass_regNext_29_3_load_store_23;
  reg                 io_in_r_bypass_regNext_29_3_df_is_ws_23;
  reg                 io_in_r_bypass_regNext_29_3_stall_23;
  reg        [15:0]   io_in_r_bypass_regNext_30_0_data_23;
  reg                 io_in_r_bypass_regNext_30_0_load_store_23;
  reg                 io_in_r_bypass_regNext_30_0_df_is_ws_23;
  reg                 io_in_r_bypass_regNext_30_0_stall_23;
  reg        [15:0]   io_in_r_bypass_regNext_30_1_data_23;
  reg                 io_in_r_bypass_regNext_30_1_load_store_23;
  reg                 io_in_r_bypass_regNext_30_1_df_is_ws_23;
  reg                 io_in_r_bypass_regNext_30_1_stall_23;
  reg        [15:0]   io_in_r_bypass_regNext_30_2_data_23;
  reg                 io_in_r_bypass_regNext_30_2_load_store_23;
  reg                 io_in_r_bypass_regNext_30_2_df_is_ws_23;
  reg                 io_in_r_bypass_regNext_30_2_stall_23;
  reg        [15:0]   io_in_r_bypass_regNext_30_3_data_23;
  reg                 io_in_r_bypass_regNext_30_3_load_store_23;
  reg                 io_in_r_bypass_regNext_30_3_df_is_ws_23;
  reg                 io_in_r_bypass_regNext_30_3_stall_23;
  reg        [15:0]   io_in_r_bypass_regNext_31_0_data_23;
  reg                 io_in_r_bypass_regNext_31_0_load_store_23;
  reg                 io_in_r_bypass_regNext_31_0_df_is_ws_23;
  reg                 io_in_r_bypass_regNext_31_0_stall_23;
  reg        [15:0]   io_in_r_bypass_regNext_31_1_data_23;
  reg                 io_in_r_bypass_regNext_31_1_load_store_23;
  reg                 io_in_r_bypass_regNext_31_1_df_is_ws_23;
  reg                 io_in_r_bypass_regNext_31_1_stall_23;
  reg        [15:0]   io_in_r_bypass_regNext_31_2_data_23;
  reg                 io_in_r_bypass_regNext_31_2_load_store_23;
  reg                 io_in_r_bypass_regNext_31_2_df_is_ws_23;
  reg                 io_in_r_bypass_regNext_31_2_stall_23;
  reg        [15:0]   io_in_r_bypass_regNext_31_3_data_23;
  reg                 io_in_r_bypass_regNext_31_3_load_store_23;
  reg                 io_in_r_bypass_regNext_31_3_df_is_ws_23;
  reg                 io_in_r_bypass_regNext_31_3_stall_23;
  reg        [15:0]   io_in_r_bypass_regNext_0_0_data_24;
  reg                 io_in_r_bypass_regNext_0_0_load_store_24;
  reg                 io_in_r_bypass_regNext_0_0_df_is_ws_24;
  reg                 io_in_r_bypass_regNext_0_0_stall_24;
  reg        [15:0]   io_in_r_bypass_regNext_0_1_data_24;
  reg                 io_in_r_bypass_regNext_0_1_load_store_24;
  reg                 io_in_r_bypass_regNext_0_1_df_is_ws_24;
  reg                 io_in_r_bypass_regNext_0_1_stall_24;
  reg        [15:0]   io_in_r_bypass_regNext_0_2_data_24;
  reg                 io_in_r_bypass_regNext_0_2_load_store_24;
  reg                 io_in_r_bypass_regNext_0_2_df_is_ws_24;
  reg                 io_in_r_bypass_regNext_0_2_stall_24;
  reg        [15:0]   io_in_r_bypass_regNext_0_3_data_24;
  reg                 io_in_r_bypass_regNext_0_3_load_store_24;
  reg                 io_in_r_bypass_regNext_0_3_df_is_ws_24;
  reg                 io_in_r_bypass_regNext_0_3_stall_24;
  reg        [15:0]   io_in_r_bypass_regNext_1_0_data_24;
  reg                 io_in_r_bypass_regNext_1_0_load_store_24;
  reg                 io_in_r_bypass_regNext_1_0_df_is_ws_24;
  reg                 io_in_r_bypass_regNext_1_0_stall_24;
  reg        [15:0]   io_in_r_bypass_regNext_1_1_data_24;
  reg                 io_in_r_bypass_regNext_1_1_load_store_24;
  reg                 io_in_r_bypass_regNext_1_1_df_is_ws_24;
  reg                 io_in_r_bypass_regNext_1_1_stall_24;
  reg        [15:0]   io_in_r_bypass_regNext_1_2_data_24;
  reg                 io_in_r_bypass_regNext_1_2_load_store_24;
  reg                 io_in_r_bypass_regNext_1_2_df_is_ws_24;
  reg                 io_in_r_bypass_regNext_1_2_stall_24;
  reg        [15:0]   io_in_r_bypass_regNext_1_3_data_24;
  reg                 io_in_r_bypass_regNext_1_3_load_store_24;
  reg                 io_in_r_bypass_regNext_1_3_df_is_ws_24;
  reg                 io_in_r_bypass_regNext_1_3_stall_24;
  reg        [15:0]   io_in_r_bypass_regNext_2_0_data_24;
  reg                 io_in_r_bypass_regNext_2_0_load_store_24;
  reg                 io_in_r_bypass_regNext_2_0_df_is_ws_24;
  reg                 io_in_r_bypass_regNext_2_0_stall_24;
  reg        [15:0]   io_in_r_bypass_regNext_2_1_data_24;
  reg                 io_in_r_bypass_regNext_2_1_load_store_24;
  reg                 io_in_r_bypass_regNext_2_1_df_is_ws_24;
  reg                 io_in_r_bypass_regNext_2_1_stall_24;
  reg        [15:0]   io_in_r_bypass_regNext_2_2_data_24;
  reg                 io_in_r_bypass_regNext_2_2_load_store_24;
  reg                 io_in_r_bypass_regNext_2_2_df_is_ws_24;
  reg                 io_in_r_bypass_regNext_2_2_stall_24;
  reg        [15:0]   io_in_r_bypass_regNext_2_3_data_24;
  reg                 io_in_r_bypass_regNext_2_3_load_store_24;
  reg                 io_in_r_bypass_regNext_2_3_df_is_ws_24;
  reg                 io_in_r_bypass_regNext_2_3_stall_24;
  reg        [15:0]   io_in_r_bypass_regNext_3_0_data_24;
  reg                 io_in_r_bypass_regNext_3_0_load_store_24;
  reg                 io_in_r_bypass_regNext_3_0_df_is_ws_24;
  reg                 io_in_r_bypass_regNext_3_0_stall_24;
  reg        [15:0]   io_in_r_bypass_regNext_3_1_data_24;
  reg                 io_in_r_bypass_regNext_3_1_load_store_24;
  reg                 io_in_r_bypass_regNext_3_1_df_is_ws_24;
  reg                 io_in_r_bypass_regNext_3_1_stall_24;
  reg        [15:0]   io_in_r_bypass_regNext_3_2_data_24;
  reg                 io_in_r_bypass_regNext_3_2_load_store_24;
  reg                 io_in_r_bypass_regNext_3_2_df_is_ws_24;
  reg                 io_in_r_bypass_regNext_3_2_stall_24;
  reg        [15:0]   io_in_r_bypass_regNext_3_3_data_24;
  reg                 io_in_r_bypass_regNext_3_3_load_store_24;
  reg                 io_in_r_bypass_regNext_3_3_df_is_ws_24;
  reg                 io_in_r_bypass_regNext_3_3_stall_24;
  reg        [15:0]   io_in_r_bypass_regNext_4_0_data_24;
  reg                 io_in_r_bypass_regNext_4_0_load_store_24;
  reg                 io_in_r_bypass_regNext_4_0_df_is_ws_24;
  reg                 io_in_r_bypass_regNext_4_0_stall_24;
  reg        [15:0]   io_in_r_bypass_regNext_4_1_data_24;
  reg                 io_in_r_bypass_regNext_4_1_load_store_24;
  reg                 io_in_r_bypass_regNext_4_1_df_is_ws_24;
  reg                 io_in_r_bypass_regNext_4_1_stall_24;
  reg        [15:0]   io_in_r_bypass_regNext_4_2_data_24;
  reg                 io_in_r_bypass_regNext_4_2_load_store_24;
  reg                 io_in_r_bypass_regNext_4_2_df_is_ws_24;
  reg                 io_in_r_bypass_regNext_4_2_stall_24;
  reg        [15:0]   io_in_r_bypass_regNext_4_3_data_24;
  reg                 io_in_r_bypass_regNext_4_3_load_store_24;
  reg                 io_in_r_bypass_regNext_4_3_df_is_ws_24;
  reg                 io_in_r_bypass_regNext_4_3_stall_24;
  reg        [15:0]   io_in_r_bypass_regNext_5_0_data_24;
  reg                 io_in_r_bypass_regNext_5_0_load_store_24;
  reg                 io_in_r_bypass_regNext_5_0_df_is_ws_24;
  reg                 io_in_r_bypass_regNext_5_0_stall_24;
  reg        [15:0]   io_in_r_bypass_regNext_5_1_data_24;
  reg                 io_in_r_bypass_regNext_5_1_load_store_24;
  reg                 io_in_r_bypass_regNext_5_1_df_is_ws_24;
  reg                 io_in_r_bypass_regNext_5_1_stall_24;
  reg        [15:0]   io_in_r_bypass_regNext_5_2_data_24;
  reg                 io_in_r_bypass_regNext_5_2_load_store_24;
  reg                 io_in_r_bypass_regNext_5_2_df_is_ws_24;
  reg                 io_in_r_bypass_regNext_5_2_stall_24;
  reg        [15:0]   io_in_r_bypass_regNext_5_3_data_24;
  reg                 io_in_r_bypass_regNext_5_3_load_store_24;
  reg                 io_in_r_bypass_regNext_5_3_df_is_ws_24;
  reg                 io_in_r_bypass_regNext_5_3_stall_24;
  reg        [15:0]   io_in_r_bypass_regNext_6_0_data_24;
  reg                 io_in_r_bypass_regNext_6_0_load_store_24;
  reg                 io_in_r_bypass_regNext_6_0_df_is_ws_24;
  reg                 io_in_r_bypass_regNext_6_0_stall_24;
  reg        [15:0]   io_in_r_bypass_regNext_6_1_data_24;
  reg                 io_in_r_bypass_regNext_6_1_load_store_24;
  reg                 io_in_r_bypass_regNext_6_1_df_is_ws_24;
  reg                 io_in_r_bypass_regNext_6_1_stall_24;
  reg        [15:0]   io_in_r_bypass_regNext_6_2_data_24;
  reg                 io_in_r_bypass_regNext_6_2_load_store_24;
  reg                 io_in_r_bypass_regNext_6_2_df_is_ws_24;
  reg                 io_in_r_bypass_regNext_6_2_stall_24;
  reg        [15:0]   io_in_r_bypass_regNext_6_3_data_24;
  reg                 io_in_r_bypass_regNext_6_3_load_store_24;
  reg                 io_in_r_bypass_regNext_6_3_df_is_ws_24;
  reg                 io_in_r_bypass_regNext_6_3_stall_24;
  reg        [15:0]   io_in_r_bypass_regNext_7_0_data_24;
  reg                 io_in_r_bypass_regNext_7_0_load_store_24;
  reg                 io_in_r_bypass_regNext_7_0_df_is_ws_24;
  reg                 io_in_r_bypass_regNext_7_0_stall_24;
  reg        [15:0]   io_in_r_bypass_regNext_7_1_data_24;
  reg                 io_in_r_bypass_regNext_7_1_load_store_24;
  reg                 io_in_r_bypass_regNext_7_1_df_is_ws_24;
  reg                 io_in_r_bypass_regNext_7_1_stall_24;
  reg        [15:0]   io_in_r_bypass_regNext_7_2_data_24;
  reg                 io_in_r_bypass_regNext_7_2_load_store_24;
  reg                 io_in_r_bypass_regNext_7_2_df_is_ws_24;
  reg                 io_in_r_bypass_regNext_7_2_stall_24;
  reg        [15:0]   io_in_r_bypass_regNext_7_3_data_24;
  reg                 io_in_r_bypass_regNext_7_3_load_store_24;
  reg                 io_in_r_bypass_regNext_7_3_df_is_ws_24;
  reg                 io_in_r_bypass_regNext_7_3_stall_24;
  reg        [15:0]   io_in_r_bypass_regNext_8_0_data_24;
  reg                 io_in_r_bypass_regNext_8_0_load_store_24;
  reg                 io_in_r_bypass_regNext_8_0_df_is_ws_24;
  reg                 io_in_r_bypass_regNext_8_0_stall_24;
  reg        [15:0]   io_in_r_bypass_regNext_8_1_data_24;
  reg                 io_in_r_bypass_regNext_8_1_load_store_24;
  reg                 io_in_r_bypass_regNext_8_1_df_is_ws_24;
  reg                 io_in_r_bypass_regNext_8_1_stall_24;
  reg        [15:0]   io_in_r_bypass_regNext_8_2_data_24;
  reg                 io_in_r_bypass_regNext_8_2_load_store_24;
  reg                 io_in_r_bypass_regNext_8_2_df_is_ws_24;
  reg                 io_in_r_bypass_regNext_8_2_stall_24;
  reg        [15:0]   io_in_r_bypass_regNext_8_3_data_24;
  reg                 io_in_r_bypass_regNext_8_3_load_store_24;
  reg                 io_in_r_bypass_regNext_8_3_df_is_ws_24;
  reg                 io_in_r_bypass_regNext_8_3_stall_24;
  reg        [15:0]   io_in_r_bypass_regNext_9_0_data_24;
  reg                 io_in_r_bypass_regNext_9_0_load_store_24;
  reg                 io_in_r_bypass_regNext_9_0_df_is_ws_24;
  reg                 io_in_r_bypass_regNext_9_0_stall_24;
  reg        [15:0]   io_in_r_bypass_regNext_9_1_data_24;
  reg                 io_in_r_bypass_regNext_9_1_load_store_24;
  reg                 io_in_r_bypass_regNext_9_1_df_is_ws_24;
  reg                 io_in_r_bypass_regNext_9_1_stall_24;
  reg        [15:0]   io_in_r_bypass_regNext_9_2_data_24;
  reg                 io_in_r_bypass_regNext_9_2_load_store_24;
  reg                 io_in_r_bypass_regNext_9_2_df_is_ws_24;
  reg                 io_in_r_bypass_regNext_9_2_stall_24;
  reg        [15:0]   io_in_r_bypass_regNext_9_3_data_24;
  reg                 io_in_r_bypass_regNext_9_3_load_store_24;
  reg                 io_in_r_bypass_regNext_9_3_df_is_ws_24;
  reg                 io_in_r_bypass_regNext_9_3_stall_24;
  reg        [15:0]   io_in_r_bypass_regNext_10_0_data_24;
  reg                 io_in_r_bypass_regNext_10_0_load_store_24;
  reg                 io_in_r_bypass_regNext_10_0_df_is_ws_24;
  reg                 io_in_r_bypass_regNext_10_0_stall_24;
  reg        [15:0]   io_in_r_bypass_regNext_10_1_data_24;
  reg                 io_in_r_bypass_regNext_10_1_load_store_24;
  reg                 io_in_r_bypass_regNext_10_1_df_is_ws_24;
  reg                 io_in_r_bypass_regNext_10_1_stall_24;
  reg        [15:0]   io_in_r_bypass_regNext_10_2_data_24;
  reg                 io_in_r_bypass_regNext_10_2_load_store_24;
  reg                 io_in_r_bypass_regNext_10_2_df_is_ws_24;
  reg                 io_in_r_bypass_regNext_10_2_stall_24;
  reg        [15:0]   io_in_r_bypass_regNext_10_3_data_24;
  reg                 io_in_r_bypass_regNext_10_3_load_store_24;
  reg                 io_in_r_bypass_regNext_10_3_df_is_ws_24;
  reg                 io_in_r_bypass_regNext_10_3_stall_24;
  reg        [15:0]   io_in_r_bypass_regNext_11_0_data_24;
  reg                 io_in_r_bypass_regNext_11_0_load_store_24;
  reg                 io_in_r_bypass_regNext_11_0_df_is_ws_24;
  reg                 io_in_r_bypass_regNext_11_0_stall_24;
  reg        [15:0]   io_in_r_bypass_regNext_11_1_data_24;
  reg                 io_in_r_bypass_regNext_11_1_load_store_24;
  reg                 io_in_r_bypass_regNext_11_1_df_is_ws_24;
  reg                 io_in_r_bypass_regNext_11_1_stall_24;
  reg        [15:0]   io_in_r_bypass_regNext_11_2_data_24;
  reg                 io_in_r_bypass_regNext_11_2_load_store_24;
  reg                 io_in_r_bypass_regNext_11_2_df_is_ws_24;
  reg                 io_in_r_bypass_regNext_11_2_stall_24;
  reg        [15:0]   io_in_r_bypass_regNext_11_3_data_24;
  reg                 io_in_r_bypass_regNext_11_3_load_store_24;
  reg                 io_in_r_bypass_regNext_11_3_df_is_ws_24;
  reg                 io_in_r_bypass_regNext_11_3_stall_24;
  reg        [15:0]   io_in_r_bypass_regNext_12_0_data_24;
  reg                 io_in_r_bypass_regNext_12_0_load_store_24;
  reg                 io_in_r_bypass_regNext_12_0_df_is_ws_24;
  reg                 io_in_r_bypass_regNext_12_0_stall_24;
  reg        [15:0]   io_in_r_bypass_regNext_12_1_data_24;
  reg                 io_in_r_bypass_regNext_12_1_load_store_24;
  reg                 io_in_r_bypass_regNext_12_1_df_is_ws_24;
  reg                 io_in_r_bypass_regNext_12_1_stall_24;
  reg        [15:0]   io_in_r_bypass_regNext_12_2_data_24;
  reg                 io_in_r_bypass_regNext_12_2_load_store_24;
  reg                 io_in_r_bypass_regNext_12_2_df_is_ws_24;
  reg                 io_in_r_bypass_regNext_12_2_stall_24;
  reg        [15:0]   io_in_r_bypass_regNext_12_3_data_24;
  reg                 io_in_r_bypass_regNext_12_3_load_store_24;
  reg                 io_in_r_bypass_regNext_12_3_df_is_ws_24;
  reg                 io_in_r_bypass_regNext_12_3_stall_24;
  reg        [15:0]   io_in_r_bypass_regNext_13_0_data_24;
  reg                 io_in_r_bypass_regNext_13_0_load_store_24;
  reg                 io_in_r_bypass_regNext_13_0_df_is_ws_24;
  reg                 io_in_r_bypass_regNext_13_0_stall_24;
  reg        [15:0]   io_in_r_bypass_regNext_13_1_data_24;
  reg                 io_in_r_bypass_regNext_13_1_load_store_24;
  reg                 io_in_r_bypass_regNext_13_1_df_is_ws_24;
  reg                 io_in_r_bypass_regNext_13_1_stall_24;
  reg        [15:0]   io_in_r_bypass_regNext_13_2_data_24;
  reg                 io_in_r_bypass_regNext_13_2_load_store_24;
  reg                 io_in_r_bypass_regNext_13_2_df_is_ws_24;
  reg                 io_in_r_bypass_regNext_13_2_stall_24;
  reg        [15:0]   io_in_r_bypass_regNext_13_3_data_24;
  reg                 io_in_r_bypass_regNext_13_3_load_store_24;
  reg                 io_in_r_bypass_regNext_13_3_df_is_ws_24;
  reg                 io_in_r_bypass_regNext_13_3_stall_24;
  reg        [15:0]   io_in_r_bypass_regNext_14_0_data_24;
  reg                 io_in_r_bypass_regNext_14_0_load_store_24;
  reg                 io_in_r_bypass_regNext_14_0_df_is_ws_24;
  reg                 io_in_r_bypass_regNext_14_0_stall_24;
  reg        [15:0]   io_in_r_bypass_regNext_14_1_data_24;
  reg                 io_in_r_bypass_regNext_14_1_load_store_24;
  reg                 io_in_r_bypass_regNext_14_1_df_is_ws_24;
  reg                 io_in_r_bypass_regNext_14_1_stall_24;
  reg        [15:0]   io_in_r_bypass_regNext_14_2_data_24;
  reg                 io_in_r_bypass_regNext_14_2_load_store_24;
  reg                 io_in_r_bypass_regNext_14_2_df_is_ws_24;
  reg                 io_in_r_bypass_regNext_14_2_stall_24;
  reg        [15:0]   io_in_r_bypass_regNext_14_3_data_24;
  reg                 io_in_r_bypass_regNext_14_3_load_store_24;
  reg                 io_in_r_bypass_regNext_14_3_df_is_ws_24;
  reg                 io_in_r_bypass_regNext_14_3_stall_24;
  reg        [15:0]   io_in_r_bypass_regNext_15_0_data_24;
  reg                 io_in_r_bypass_regNext_15_0_load_store_24;
  reg                 io_in_r_bypass_regNext_15_0_df_is_ws_24;
  reg                 io_in_r_bypass_regNext_15_0_stall_24;
  reg        [15:0]   io_in_r_bypass_regNext_15_1_data_24;
  reg                 io_in_r_bypass_regNext_15_1_load_store_24;
  reg                 io_in_r_bypass_regNext_15_1_df_is_ws_24;
  reg                 io_in_r_bypass_regNext_15_1_stall_24;
  reg        [15:0]   io_in_r_bypass_regNext_15_2_data_24;
  reg                 io_in_r_bypass_regNext_15_2_load_store_24;
  reg                 io_in_r_bypass_regNext_15_2_df_is_ws_24;
  reg                 io_in_r_bypass_regNext_15_2_stall_24;
  reg        [15:0]   io_in_r_bypass_regNext_15_3_data_24;
  reg                 io_in_r_bypass_regNext_15_3_load_store_24;
  reg                 io_in_r_bypass_regNext_15_3_df_is_ws_24;
  reg                 io_in_r_bypass_regNext_15_3_stall_24;
  reg        [15:0]   io_in_r_bypass_regNext_16_0_data_24;
  reg                 io_in_r_bypass_regNext_16_0_load_store_24;
  reg                 io_in_r_bypass_regNext_16_0_df_is_ws_24;
  reg                 io_in_r_bypass_regNext_16_0_stall_24;
  reg        [15:0]   io_in_r_bypass_regNext_16_1_data_24;
  reg                 io_in_r_bypass_regNext_16_1_load_store_24;
  reg                 io_in_r_bypass_regNext_16_1_df_is_ws_24;
  reg                 io_in_r_bypass_regNext_16_1_stall_24;
  reg        [15:0]   io_in_r_bypass_regNext_16_2_data_24;
  reg                 io_in_r_bypass_regNext_16_2_load_store_24;
  reg                 io_in_r_bypass_regNext_16_2_df_is_ws_24;
  reg                 io_in_r_bypass_regNext_16_2_stall_24;
  reg        [15:0]   io_in_r_bypass_regNext_16_3_data_24;
  reg                 io_in_r_bypass_regNext_16_3_load_store_24;
  reg                 io_in_r_bypass_regNext_16_3_df_is_ws_24;
  reg                 io_in_r_bypass_regNext_16_3_stall_24;
  reg        [15:0]   io_in_r_bypass_regNext_17_0_data_24;
  reg                 io_in_r_bypass_regNext_17_0_load_store_24;
  reg                 io_in_r_bypass_regNext_17_0_df_is_ws_24;
  reg                 io_in_r_bypass_regNext_17_0_stall_24;
  reg        [15:0]   io_in_r_bypass_regNext_17_1_data_24;
  reg                 io_in_r_bypass_regNext_17_1_load_store_24;
  reg                 io_in_r_bypass_regNext_17_1_df_is_ws_24;
  reg                 io_in_r_bypass_regNext_17_1_stall_24;
  reg        [15:0]   io_in_r_bypass_regNext_17_2_data_24;
  reg                 io_in_r_bypass_regNext_17_2_load_store_24;
  reg                 io_in_r_bypass_regNext_17_2_df_is_ws_24;
  reg                 io_in_r_bypass_regNext_17_2_stall_24;
  reg        [15:0]   io_in_r_bypass_regNext_17_3_data_24;
  reg                 io_in_r_bypass_regNext_17_3_load_store_24;
  reg                 io_in_r_bypass_regNext_17_3_df_is_ws_24;
  reg                 io_in_r_bypass_regNext_17_3_stall_24;
  reg        [15:0]   io_in_r_bypass_regNext_18_0_data_24;
  reg                 io_in_r_bypass_regNext_18_0_load_store_24;
  reg                 io_in_r_bypass_regNext_18_0_df_is_ws_24;
  reg                 io_in_r_bypass_regNext_18_0_stall_24;
  reg        [15:0]   io_in_r_bypass_regNext_18_1_data_24;
  reg                 io_in_r_bypass_regNext_18_1_load_store_24;
  reg                 io_in_r_bypass_regNext_18_1_df_is_ws_24;
  reg                 io_in_r_bypass_regNext_18_1_stall_24;
  reg        [15:0]   io_in_r_bypass_regNext_18_2_data_24;
  reg                 io_in_r_bypass_regNext_18_2_load_store_24;
  reg                 io_in_r_bypass_regNext_18_2_df_is_ws_24;
  reg                 io_in_r_bypass_regNext_18_2_stall_24;
  reg        [15:0]   io_in_r_bypass_regNext_18_3_data_24;
  reg                 io_in_r_bypass_regNext_18_3_load_store_24;
  reg                 io_in_r_bypass_regNext_18_3_df_is_ws_24;
  reg                 io_in_r_bypass_regNext_18_3_stall_24;
  reg        [15:0]   io_in_r_bypass_regNext_19_0_data_24;
  reg                 io_in_r_bypass_regNext_19_0_load_store_24;
  reg                 io_in_r_bypass_regNext_19_0_df_is_ws_24;
  reg                 io_in_r_bypass_regNext_19_0_stall_24;
  reg        [15:0]   io_in_r_bypass_regNext_19_1_data_24;
  reg                 io_in_r_bypass_regNext_19_1_load_store_24;
  reg                 io_in_r_bypass_regNext_19_1_df_is_ws_24;
  reg                 io_in_r_bypass_regNext_19_1_stall_24;
  reg        [15:0]   io_in_r_bypass_regNext_19_2_data_24;
  reg                 io_in_r_bypass_regNext_19_2_load_store_24;
  reg                 io_in_r_bypass_regNext_19_2_df_is_ws_24;
  reg                 io_in_r_bypass_regNext_19_2_stall_24;
  reg        [15:0]   io_in_r_bypass_regNext_19_3_data_24;
  reg                 io_in_r_bypass_regNext_19_3_load_store_24;
  reg                 io_in_r_bypass_regNext_19_3_df_is_ws_24;
  reg                 io_in_r_bypass_regNext_19_3_stall_24;
  reg        [15:0]   io_in_r_bypass_regNext_20_0_data_24;
  reg                 io_in_r_bypass_regNext_20_0_load_store_24;
  reg                 io_in_r_bypass_regNext_20_0_df_is_ws_24;
  reg                 io_in_r_bypass_regNext_20_0_stall_24;
  reg        [15:0]   io_in_r_bypass_regNext_20_1_data_24;
  reg                 io_in_r_bypass_regNext_20_1_load_store_24;
  reg                 io_in_r_bypass_regNext_20_1_df_is_ws_24;
  reg                 io_in_r_bypass_regNext_20_1_stall_24;
  reg        [15:0]   io_in_r_bypass_regNext_20_2_data_24;
  reg                 io_in_r_bypass_regNext_20_2_load_store_24;
  reg                 io_in_r_bypass_regNext_20_2_df_is_ws_24;
  reg                 io_in_r_bypass_regNext_20_2_stall_24;
  reg        [15:0]   io_in_r_bypass_regNext_20_3_data_24;
  reg                 io_in_r_bypass_regNext_20_3_load_store_24;
  reg                 io_in_r_bypass_regNext_20_3_df_is_ws_24;
  reg                 io_in_r_bypass_regNext_20_3_stall_24;
  reg        [15:0]   io_in_r_bypass_regNext_21_0_data_24;
  reg                 io_in_r_bypass_regNext_21_0_load_store_24;
  reg                 io_in_r_bypass_regNext_21_0_df_is_ws_24;
  reg                 io_in_r_bypass_regNext_21_0_stall_24;
  reg        [15:0]   io_in_r_bypass_regNext_21_1_data_24;
  reg                 io_in_r_bypass_regNext_21_1_load_store_24;
  reg                 io_in_r_bypass_regNext_21_1_df_is_ws_24;
  reg                 io_in_r_bypass_regNext_21_1_stall_24;
  reg        [15:0]   io_in_r_bypass_regNext_21_2_data_24;
  reg                 io_in_r_bypass_regNext_21_2_load_store_24;
  reg                 io_in_r_bypass_regNext_21_2_df_is_ws_24;
  reg                 io_in_r_bypass_regNext_21_2_stall_24;
  reg        [15:0]   io_in_r_bypass_regNext_21_3_data_24;
  reg                 io_in_r_bypass_regNext_21_3_load_store_24;
  reg                 io_in_r_bypass_regNext_21_3_df_is_ws_24;
  reg                 io_in_r_bypass_regNext_21_3_stall_24;
  reg        [15:0]   io_in_r_bypass_regNext_22_0_data_24;
  reg                 io_in_r_bypass_regNext_22_0_load_store_24;
  reg                 io_in_r_bypass_regNext_22_0_df_is_ws_24;
  reg                 io_in_r_bypass_regNext_22_0_stall_24;
  reg        [15:0]   io_in_r_bypass_regNext_22_1_data_24;
  reg                 io_in_r_bypass_regNext_22_1_load_store_24;
  reg                 io_in_r_bypass_regNext_22_1_df_is_ws_24;
  reg                 io_in_r_bypass_regNext_22_1_stall_24;
  reg        [15:0]   io_in_r_bypass_regNext_22_2_data_24;
  reg                 io_in_r_bypass_regNext_22_2_load_store_24;
  reg                 io_in_r_bypass_regNext_22_2_df_is_ws_24;
  reg                 io_in_r_bypass_regNext_22_2_stall_24;
  reg        [15:0]   io_in_r_bypass_regNext_22_3_data_24;
  reg                 io_in_r_bypass_regNext_22_3_load_store_24;
  reg                 io_in_r_bypass_regNext_22_3_df_is_ws_24;
  reg                 io_in_r_bypass_regNext_22_3_stall_24;
  reg        [15:0]   io_in_r_bypass_regNext_23_0_data_24;
  reg                 io_in_r_bypass_regNext_23_0_load_store_24;
  reg                 io_in_r_bypass_regNext_23_0_df_is_ws_24;
  reg                 io_in_r_bypass_regNext_23_0_stall_24;
  reg        [15:0]   io_in_r_bypass_regNext_23_1_data_24;
  reg                 io_in_r_bypass_regNext_23_1_load_store_24;
  reg                 io_in_r_bypass_regNext_23_1_df_is_ws_24;
  reg                 io_in_r_bypass_regNext_23_1_stall_24;
  reg        [15:0]   io_in_r_bypass_regNext_23_2_data_24;
  reg                 io_in_r_bypass_regNext_23_2_load_store_24;
  reg                 io_in_r_bypass_regNext_23_2_df_is_ws_24;
  reg                 io_in_r_bypass_regNext_23_2_stall_24;
  reg        [15:0]   io_in_r_bypass_regNext_23_3_data_24;
  reg                 io_in_r_bypass_regNext_23_3_load_store_24;
  reg                 io_in_r_bypass_regNext_23_3_df_is_ws_24;
  reg                 io_in_r_bypass_regNext_23_3_stall_24;
  reg        [15:0]   io_in_r_bypass_regNext_24_0_data_24;
  reg                 io_in_r_bypass_regNext_24_0_load_store_24;
  reg                 io_in_r_bypass_regNext_24_0_df_is_ws_24;
  reg                 io_in_r_bypass_regNext_24_0_stall_24;
  reg        [15:0]   io_in_r_bypass_regNext_24_1_data_24;
  reg                 io_in_r_bypass_regNext_24_1_load_store_24;
  reg                 io_in_r_bypass_regNext_24_1_df_is_ws_24;
  reg                 io_in_r_bypass_regNext_24_1_stall_24;
  reg        [15:0]   io_in_r_bypass_regNext_24_2_data_24;
  reg                 io_in_r_bypass_regNext_24_2_load_store_24;
  reg                 io_in_r_bypass_regNext_24_2_df_is_ws_24;
  reg                 io_in_r_bypass_regNext_24_2_stall_24;
  reg        [15:0]   io_in_r_bypass_regNext_24_3_data_24;
  reg                 io_in_r_bypass_regNext_24_3_load_store_24;
  reg                 io_in_r_bypass_regNext_24_3_df_is_ws_24;
  reg                 io_in_r_bypass_regNext_24_3_stall_24;
  reg        [15:0]   io_in_r_bypass_regNext_25_0_data_24;
  reg                 io_in_r_bypass_regNext_25_0_load_store_24;
  reg                 io_in_r_bypass_regNext_25_0_df_is_ws_24;
  reg                 io_in_r_bypass_regNext_25_0_stall_24;
  reg        [15:0]   io_in_r_bypass_regNext_25_1_data_24;
  reg                 io_in_r_bypass_regNext_25_1_load_store_24;
  reg                 io_in_r_bypass_regNext_25_1_df_is_ws_24;
  reg                 io_in_r_bypass_regNext_25_1_stall_24;
  reg        [15:0]   io_in_r_bypass_regNext_25_2_data_24;
  reg                 io_in_r_bypass_regNext_25_2_load_store_24;
  reg                 io_in_r_bypass_regNext_25_2_df_is_ws_24;
  reg                 io_in_r_bypass_regNext_25_2_stall_24;
  reg        [15:0]   io_in_r_bypass_regNext_25_3_data_24;
  reg                 io_in_r_bypass_regNext_25_3_load_store_24;
  reg                 io_in_r_bypass_regNext_25_3_df_is_ws_24;
  reg                 io_in_r_bypass_regNext_25_3_stall_24;
  reg        [15:0]   io_in_r_bypass_regNext_26_0_data_24;
  reg                 io_in_r_bypass_regNext_26_0_load_store_24;
  reg                 io_in_r_bypass_regNext_26_0_df_is_ws_24;
  reg                 io_in_r_bypass_regNext_26_0_stall_24;
  reg        [15:0]   io_in_r_bypass_regNext_26_1_data_24;
  reg                 io_in_r_bypass_regNext_26_1_load_store_24;
  reg                 io_in_r_bypass_regNext_26_1_df_is_ws_24;
  reg                 io_in_r_bypass_regNext_26_1_stall_24;
  reg        [15:0]   io_in_r_bypass_regNext_26_2_data_24;
  reg                 io_in_r_bypass_regNext_26_2_load_store_24;
  reg                 io_in_r_bypass_regNext_26_2_df_is_ws_24;
  reg                 io_in_r_bypass_regNext_26_2_stall_24;
  reg        [15:0]   io_in_r_bypass_regNext_26_3_data_24;
  reg                 io_in_r_bypass_regNext_26_3_load_store_24;
  reg                 io_in_r_bypass_regNext_26_3_df_is_ws_24;
  reg                 io_in_r_bypass_regNext_26_3_stall_24;
  reg        [15:0]   io_in_r_bypass_regNext_27_0_data_24;
  reg                 io_in_r_bypass_regNext_27_0_load_store_24;
  reg                 io_in_r_bypass_regNext_27_0_df_is_ws_24;
  reg                 io_in_r_bypass_regNext_27_0_stall_24;
  reg        [15:0]   io_in_r_bypass_regNext_27_1_data_24;
  reg                 io_in_r_bypass_regNext_27_1_load_store_24;
  reg                 io_in_r_bypass_regNext_27_1_df_is_ws_24;
  reg                 io_in_r_bypass_regNext_27_1_stall_24;
  reg        [15:0]   io_in_r_bypass_regNext_27_2_data_24;
  reg                 io_in_r_bypass_regNext_27_2_load_store_24;
  reg                 io_in_r_bypass_regNext_27_2_df_is_ws_24;
  reg                 io_in_r_bypass_regNext_27_2_stall_24;
  reg        [15:0]   io_in_r_bypass_regNext_27_3_data_24;
  reg                 io_in_r_bypass_regNext_27_3_load_store_24;
  reg                 io_in_r_bypass_regNext_27_3_df_is_ws_24;
  reg                 io_in_r_bypass_regNext_27_3_stall_24;
  reg        [15:0]   io_in_r_bypass_regNext_28_0_data_24;
  reg                 io_in_r_bypass_regNext_28_0_load_store_24;
  reg                 io_in_r_bypass_regNext_28_0_df_is_ws_24;
  reg                 io_in_r_bypass_regNext_28_0_stall_24;
  reg        [15:0]   io_in_r_bypass_regNext_28_1_data_24;
  reg                 io_in_r_bypass_regNext_28_1_load_store_24;
  reg                 io_in_r_bypass_regNext_28_1_df_is_ws_24;
  reg                 io_in_r_bypass_regNext_28_1_stall_24;
  reg        [15:0]   io_in_r_bypass_regNext_28_2_data_24;
  reg                 io_in_r_bypass_regNext_28_2_load_store_24;
  reg                 io_in_r_bypass_regNext_28_2_df_is_ws_24;
  reg                 io_in_r_bypass_regNext_28_2_stall_24;
  reg        [15:0]   io_in_r_bypass_regNext_28_3_data_24;
  reg                 io_in_r_bypass_regNext_28_3_load_store_24;
  reg                 io_in_r_bypass_regNext_28_3_df_is_ws_24;
  reg                 io_in_r_bypass_regNext_28_3_stall_24;
  reg        [15:0]   io_in_r_bypass_regNext_29_0_data_24;
  reg                 io_in_r_bypass_regNext_29_0_load_store_24;
  reg                 io_in_r_bypass_regNext_29_0_df_is_ws_24;
  reg                 io_in_r_bypass_regNext_29_0_stall_24;
  reg        [15:0]   io_in_r_bypass_regNext_29_1_data_24;
  reg                 io_in_r_bypass_regNext_29_1_load_store_24;
  reg                 io_in_r_bypass_regNext_29_1_df_is_ws_24;
  reg                 io_in_r_bypass_regNext_29_1_stall_24;
  reg        [15:0]   io_in_r_bypass_regNext_29_2_data_24;
  reg                 io_in_r_bypass_regNext_29_2_load_store_24;
  reg                 io_in_r_bypass_regNext_29_2_df_is_ws_24;
  reg                 io_in_r_bypass_regNext_29_2_stall_24;
  reg        [15:0]   io_in_r_bypass_regNext_29_3_data_24;
  reg                 io_in_r_bypass_regNext_29_3_load_store_24;
  reg                 io_in_r_bypass_regNext_29_3_df_is_ws_24;
  reg                 io_in_r_bypass_regNext_29_3_stall_24;
  reg        [15:0]   io_in_r_bypass_regNext_30_0_data_24;
  reg                 io_in_r_bypass_regNext_30_0_load_store_24;
  reg                 io_in_r_bypass_regNext_30_0_df_is_ws_24;
  reg                 io_in_r_bypass_regNext_30_0_stall_24;
  reg        [15:0]   io_in_r_bypass_regNext_30_1_data_24;
  reg                 io_in_r_bypass_regNext_30_1_load_store_24;
  reg                 io_in_r_bypass_regNext_30_1_df_is_ws_24;
  reg                 io_in_r_bypass_regNext_30_1_stall_24;
  reg        [15:0]   io_in_r_bypass_regNext_30_2_data_24;
  reg                 io_in_r_bypass_regNext_30_2_load_store_24;
  reg                 io_in_r_bypass_regNext_30_2_df_is_ws_24;
  reg                 io_in_r_bypass_regNext_30_2_stall_24;
  reg        [15:0]   io_in_r_bypass_regNext_30_3_data_24;
  reg                 io_in_r_bypass_regNext_30_3_load_store_24;
  reg                 io_in_r_bypass_regNext_30_3_df_is_ws_24;
  reg                 io_in_r_bypass_regNext_30_3_stall_24;
  reg        [15:0]   io_in_r_bypass_regNext_31_0_data_24;
  reg                 io_in_r_bypass_regNext_31_0_load_store_24;
  reg                 io_in_r_bypass_regNext_31_0_df_is_ws_24;
  reg                 io_in_r_bypass_regNext_31_0_stall_24;
  reg        [15:0]   io_in_r_bypass_regNext_31_1_data_24;
  reg                 io_in_r_bypass_regNext_31_1_load_store_24;
  reg                 io_in_r_bypass_regNext_31_1_df_is_ws_24;
  reg                 io_in_r_bypass_regNext_31_1_stall_24;
  reg        [15:0]   io_in_r_bypass_regNext_31_2_data_24;
  reg                 io_in_r_bypass_regNext_31_2_load_store_24;
  reg                 io_in_r_bypass_regNext_31_2_df_is_ws_24;
  reg                 io_in_r_bypass_regNext_31_2_stall_24;
  reg        [15:0]   io_in_r_bypass_regNext_31_3_data_24;
  reg                 io_in_r_bypass_regNext_31_3_load_store_24;
  reg                 io_in_r_bypass_regNext_31_3_df_is_ws_24;
  reg                 io_in_r_bypass_regNext_31_3_stall_24;
  reg        [15:0]   io_in_r_bypass_regNext_0_0_data_25;
  reg                 io_in_r_bypass_regNext_0_0_load_store_25;
  reg                 io_in_r_bypass_regNext_0_0_df_is_ws_25;
  reg                 io_in_r_bypass_regNext_0_0_stall_25;
  reg        [15:0]   io_in_r_bypass_regNext_0_1_data_25;
  reg                 io_in_r_bypass_regNext_0_1_load_store_25;
  reg                 io_in_r_bypass_regNext_0_1_df_is_ws_25;
  reg                 io_in_r_bypass_regNext_0_1_stall_25;
  reg        [15:0]   io_in_r_bypass_regNext_0_2_data_25;
  reg                 io_in_r_bypass_regNext_0_2_load_store_25;
  reg                 io_in_r_bypass_regNext_0_2_df_is_ws_25;
  reg                 io_in_r_bypass_regNext_0_2_stall_25;
  reg        [15:0]   io_in_r_bypass_regNext_0_3_data_25;
  reg                 io_in_r_bypass_regNext_0_3_load_store_25;
  reg                 io_in_r_bypass_regNext_0_3_df_is_ws_25;
  reg                 io_in_r_bypass_regNext_0_3_stall_25;
  reg        [15:0]   io_in_r_bypass_regNext_1_0_data_25;
  reg                 io_in_r_bypass_regNext_1_0_load_store_25;
  reg                 io_in_r_bypass_regNext_1_0_df_is_ws_25;
  reg                 io_in_r_bypass_regNext_1_0_stall_25;
  reg        [15:0]   io_in_r_bypass_regNext_1_1_data_25;
  reg                 io_in_r_bypass_regNext_1_1_load_store_25;
  reg                 io_in_r_bypass_regNext_1_1_df_is_ws_25;
  reg                 io_in_r_bypass_regNext_1_1_stall_25;
  reg        [15:0]   io_in_r_bypass_regNext_1_2_data_25;
  reg                 io_in_r_bypass_regNext_1_2_load_store_25;
  reg                 io_in_r_bypass_regNext_1_2_df_is_ws_25;
  reg                 io_in_r_bypass_regNext_1_2_stall_25;
  reg        [15:0]   io_in_r_bypass_regNext_1_3_data_25;
  reg                 io_in_r_bypass_regNext_1_3_load_store_25;
  reg                 io_in_r_bypass_regNext_1_3_df_is_ws_25;
  reg                 io_in_r_bypass_regNext_1_3_stall_25;
  reg        [15:0]   io_in_r_bypass_regNext_2_0_data_25;
  reg                 io_in_r_bypass_regNext_2_0_load_store_25;
  reg                 io_in_r_bypass_regNext_2_0_df_is_ws_25;
  reg                 io_in_r_bypass_regNext_2_0_stall_25;
  reg        [15:0]   io_in_r_bypass_regNext_2_1_data_25;
  reg                 io_in_r_bypass_regNext_2_1_load_store_25;
  reg                 io_in_r_bypass_regNext_2_1_df_is_ws_25;
  reg                 io_in_r_bypass_regNext_2_1_stall_25;
  reg        [15:0]   io_in_r_bypass_regNext_2_2_data_25;
  reg                 io_in_r_bypass_regNext_2_2_load_store_25;
  reg                 io_in_r_bypass_regNext_2_2_df_is_ws_25;
  reg                 io_in_r_bypass_regNext_2_2_stall_25;
  reg        [15:0]   io_in_r_bypass_regNext_2_3_data_25;
  reg                 io_in_r_bypass_regNext_2_3_load_store_25;
  reg                 io_in_r_bypass_regNext_2_3_df_is_ws_25;
  reg                 io_in_r_bypass_regNext_2_3_stall_25;
  reg        [15:0]   io_in_r_bypass_regNext_3_0_data_25;
  reg                 io_in_r_bypass_regNext_3_0_load_store_25;
  reg                 io_in_r_bypass_regNext_3_0_df_is_ws_25;
  reg                 io_in_r_bypass_regNext_3_0_stall_25;
  reg        [15:0]   io_in_r_bypass_regNext_3_1_data_25;
  reg                 io_in_r_bypass_regNext_3_1_load_store_25;
  reg                 io_in_r_bypass_regNext_3_1_df_is_ws_25;
  reg                 io_in_r_bypass_regNext_3_1_stall_25;
  reg        [15:0]   io_in_r_bypass_regNext_3_2_data_25;
  reg                 io_in_r_bypass_regNext_3_2_load_store_25;
  reg                 io_in_r_bypass_regNext_3_2_df_is_ws_25;
  reg                 io_in_r_bypass_regNext_3_2_stall_25;
  reg        [15:0]   io_in_r_bypass_regNext_3_3_data_25;
  reg                 io_in_r_bypass_regNext_3_3_load_store_25;
  reg                 io_in_r_bypass_regNext_3_3_df_is_ws_25;
  reg                 io_in_r_bypass_regNext_3_3_stall_25;
  reg        [15:0]   io_in_r_bypass_regNext_4_0_data_25;
  reg                 io_in_r_bypass_regNext_4_0_load_store_25;
  reg                 io_in_r_bypass_regNext_4_0_df_is_ws_25;
  reg                 io_in_r_bypass_regNext_4_0_stall_25;
  reg        [15:0]   io_in_r_bypass_regNext_4_1_data_25;
  reg                 io_in_r_bypass_regNext_4_1_load_store_25;
  reg                 io_in_r_bypass_regNext_4_1_df_is_ws_25;
  reg                 io_in_r_bypass_regNext_4_1_stall_25;
  reg        [15:0]   io_in_r_bypass_regNext_4_2_data_25;
  reg                 io_in_r_bypass_regNext_4_2_load_store_25;
  reg                 io_in_r_bypass_regNext_4_2_df_is_ws_25;
  reg                 io_in_r_bypass_regNext_4_2_stall_25;
  reg        [15:0]   io_in_r_bypass_regNext_4_3_data_25;
  reg                 io_in_r_bypass_regNext_4_3_load_store_25;
  reg                 io_in_r_bypass_regNext_4_3_df_is_ws_25;
  reg                 io_in_r_bypass_regNext_4_3_stall_25;
  reg        [15:0]   io_in_r_bypass_regNext_5_0_data_25;
  reg                 io_in_r_bypass_regNext_5_0_load_store_25;
  reg                 io_in_r_bypass_regNext_5_0_df_is_ws_25;
  reg                 io_in_r_bypass_regNext_5_0_stall_25;
  reg        [15:0]   io_in_r_bypass_regNext_5_1_data_25;
  reg                 io_in_r_bypass_regNext_5_1_load_store_25;
  reg                 io_in_r_bypass_regNext_5_1_df_is_ws_25;
  reg                 io_in_r_bypass_regNext_5_1_stall_25;
  reg        [15:0]   io_in_r_bypass_regNext_5_2_data_25;
  reg                 io_in_r_bypass_regNext_5_2_load_store_25;
  reg                 io_in_r_bypass_regNext_5_2_df_is_ws_25;
  reg                 io_in_r_bypass_regNext_5_2_stall_25;
  reg        [15:0]   io_in_r_bypass_regNext_5_3_data_25;
  reg                 io_in_r_bypass_regNext_5_3_load_store_25;
  reg                 io_in_r_bypass_regNext_5_3_df_is_ws_25;
  reg                 io_in_r_bypass_regNext_5_3_stall_25;
  reg        [15:0]   io_in_r_bypass_regNext_6_0_data_25;
  reg                 io_in_r_bypass_regNext_6_0_load_store_25;
  reg                 io_in_r_bypass_regNext_6_0_df_is_ws_25;
  reg                 io_in_r_bypass_regNext_6_0_stall_25;
  reg        [15:0]   io_in_r_bypass_regNext_6_1_data_25;
  reg                 io_in_r_bypass_regNext_6_1_load_store_25;
  reg                 io_in_r_bypass_regNext_6_1_df_is_ws_25;
  reg                 io_in_r_bypass_regNext_6_1_stall_25;
  reg        [15:0]   io_in_r_bypass_regNext_6_2_data_25;
  reg                 io_in_r_bypass_regNext_6_2_load_store_25;
  reg                 io_in_r_bypass_regNext_6_2_df_is_ws_25;
  reg                 io_in_r_bypass_regNext_6_2_stall_25;
  reg        [15:0]   io_in_r_bypass_regNext_6_3_data_25;
  reg                 io_in_r_bypass_regNext_6_3_load_store_25;
  reg                 io_in_r_bypass_regNext_6_3_df_is_ws_25;
  reg                 io_in_r_bypass_regNext_6_3_stall_25;
  reg        [15:0]   io_in_r_bypass_regNext_7_0_data_25;
  reg                 io_in_r_bypass_regNext_7_0_load_store_25;
  reg                 io_in_r_bypass_regNext_7_0_df_is_ws_25;
  reg                 io_in_r_bypass_regNext_7_0_stall_25;
  reg        [15:0]   io_in_r_bypass_regNext_7_1_data_25;
  reg                 io_in_r_bypass_regNext_7_1_load_store_25;
  reg                 io_in_r_bypass_regNext_7_1_df_is_ws_25;
  reg                 io_in_r_bypass_regNext_7_1_stall_25;
  reg        [15:0]   io_in_r_bypass_regNext_7_2_data_25;
  reg                 io_in_r_bypass_regNext_7_2_load_store_25;
  reg                 io_in_r_bypass_regNext_7_2_df_is_ws_25;
  reg                 io_in_r_bypass_regNext_7_2_stall_25;
  reg        [15:0]   io_in_r_bypass_regNext_7_3_data_25;
  reg                 io_in_r_bypass_regNext_7_3_load_store_25;
  reg                 io_in_r_bypass_regNext_7_3_df_is_ws_25;
  reg                 io_in_r_bypass_regNext_7_3_stall_25;
  reg        [15:0]   io_in_r_bypass_regNext_8_0_data_25;
  reg                 io_in_r_bypass_regNext_8_0_load_store_25;
  reg                 io_in_r_bypass_regNext_8_0_df_is_ws_25;
  reg                 io_in_r_bypass_regNext_8_0_stall_25;
  reg        [15:0]   io_in_r_bypass_regNext_8_1_data_25;
  reg                 io_in_r_bypass_regNext_8_1_load_store_25;
  reg                 io_in_r_bypass_regNext_8_1_df_is_ws_25;
  reg                 io_in_r_bypass_regNext_8_1_stall_25;
  reg        [15:0]   io_in_r_bypass_regNext_8_2_data_25;
  reg                 io_in_r_bypass_regNext_8_2_load_store_25;
  reg                 io_in_r_bypass_regNext_8_2_df_is_ws_25;
  reg                 io_in_r_bypass_regNext_8_2_stall_25;
  reg        [15:0]   io_in_r_bypass_regNext_8_3_data_25;
  reg                 io_in_r_bypass_regNext_8_3_load_store_25;
  reg                 io_in_r_bypass_regNext_8_3_df_is_ws_25;
  reg                 io_in_r_bypass_regNext_8_3_stall_25;
  reg        [15:0]   io_in_r_bypass_regNext_9_0_data_25;
  reg                 io_in_r_bypass_regNext_9_0_load_store_25;
  reg                 io_in_r_bypass_regNext_9_0_df_is_ws_25;
  reg                 io_in_r_bypass_regNext_9_0_stall_25;
  reg        [15:0]   io_in_r_bypass_regNext_9_1_data_25;
  reg                 io_in_r_bypass_regNext_9_1_load_store_25;
  reg                 io_in_r_bypass_regNext_9_1_df_is_ws_25;
  reg                 io_in_r_bypass_regNext_9_1_stall_25;
  reg        [15:0]   io_in_r_bypass_regNext_9_2_data_25;
  reg                 io_in_r_bypass_regNext_9_2_load_store_25;
  reg                 io_in_r_bypass_regNext_9_2_df_is_ws_25;
  reg                 io_in_r_bypass_regNext_9_2_stall_25;
  reg        [15:0]   io_in_r_bypass_regNext_9_3_data_25;
  reg                 io_in_r_bypass_regNext_9_3_load_store_25;
  reg                 io_in_r_bypass_regNext_9_3_df_is_ws_25;
  reg                 io_in_r_bypass_regNext_9_3_stall_25;
  reg        [15:0]   io_in_r_bypass_regNext_10_0_data_25;
  reg                 io_in_r_bypass_regNext_10_0_load_store_25;
  reg                 io_in_r_bypass_regNext_10_0_df_is_ws_25;
  reg                 io_in_r_bypass_regNext_10_0_stall_25;
  reg        [15:0]   io_in_r_bypass_regNext_10_1_data_25;
  reg                 io_in_r_bypass_regNext_10_1_load_store_25;
  reg                 io_in_r_bypass_regNext_10_1_df_is_ws_25;
  reg                 io_in_r_bypass_regNext_10_1_stall_25;
  reg        [15:0]   io_in_r_bypass_regNext_10_2_data_25;
  reg                 io_in_r_bypass_regNext_10_2_load_store_25;
  reg                 io_in_r_bypass_regNext_10_2_df_is_ws_25;
  reg                 io_in_r_bypass_regNext_10_2_stall_25;
  reg        [15:0]   io_in_r_bypass_regNext_10_3_data_25;
  reg                 io_in_r_bypass_regNext_10_3_load_store_25;
  reg                 io_in_r_bypass_regNext_10_3_df_is_ws_25;
  reg                 io_in_r_bypass_regNext_10_3_stall_25;
  reg        [15:0]   io_in_r_bypass_regNext_11_0_data_25;
  reg                 io_in_r_bypass_regNext_11_0_load_store_25;
  reg                 io_in_r_bypass_regNext_11_0_df_is_ws_25;
  reg                 io_in_r_bypass_regNext_11_0_stall_25;
  reg        [15:0]   io_in_r_bypass_regNext_11_1_data_25;
  reg                 io_in_r_bypass_regNext_11_1_load_store_25;
  reg                 io_in_r_bypass_regNext_11_1_df_is_ws_25;
  reg                 io_in_r_bypass_regNext_11_1_stall_25;
  reg        [15:0]   io_in_r_bypass_regNext_11_2_data_25;
  reg                 io_in_r_bypass_regNext_11_2_load_store_25;
  reg                 io_in_r_bypass_regNext_11_2_df_is_ws_25;
  reg                 io_in_r_bypass_regNext_11_2_stall_25;
  reg        [15:0]   io_in_r_bypass_regNext_11_3_data_25;
  reg                 io_in_r_bypass_regNext_11_3_load_store_25;
  reg                 io_in_r_bypass_regNext_11_3_df_is_ws_25;
  reg                 io_in_r_bypass_regNext_11_3_stall_25;
  reg        [15:0]   io_in_r_bypass_regNext_12_0_data_25;
  reg                 io_in_r_bypass_regNext_12_0_load_store_25;
  reg                 io_in_r_bypass_regNext_12_0_df_is_ws_25;
  reg                 io_in_r_bypass_regNext_12_0_stall_25;
  reg        [15:0]   io_in_r_bypass_regNext_12_1_data_25;
  reg                 io_in_r_bypass_regNext_12_1_load_store_25;
  reg                 io_in_r_bypass_regNext_12_1_df_is_ws_25;
  reg                 io_in_r_bypass_regNext_12_1_stall_25;
  reg        [15:0]   io_in_r_bypass_regNext_12_2_data_25;
  reg                 io_in_r_bypass_regNext_12_2_load_store_25;
  reg                 io_in_r_bypass_regNext_12_2_df_is_ws_25;
  reg                 io_in_r_bypass_regNext_12_2_stall_25;
  reg        [15:0]   io_in_r_bypass_regNext_12_3_data_25;
  reg                 io_in_r_bypass_regNext_12_3_load_store_25;
  reg                 io_in_r_bypass_regNext_12_3_df_is_ws_25;
  reg                 io_in_r_bypass_regNext_12_3_stall_25;
  reg        [15:0]   io_in_r_bypass_regNext_13_0_data_25;
  reg                 io_in_r_bypass_regNext_13_0_load_store_25;
  reg                 io_in_r_bypass_regNext_13_0_df_is_ws_25;
  reg                 io_in_r_bypass_regNext_13_0_stall_25;
  reg        [15:0]   io_in_r_bypass_regNext_13_1_data_25;
  reg                 io_in_r_bypass_regNext_13_1_load_store_25;
  reg                 io_in_r_bypass_regNext_13_1_df_is_ws_25;
  reg                 io_in_r_bypass_regNext_13_1_stall_25;
  reg        [15:0]   io_in_r_bypass_regNext_13_2_data_25;
  reg                 io_in_r_bypass_regNext_13_2_load_store_25;
  reg                 io_in_r_bypass_regNext_13_2_df_is_ws_25;
  reg                 io_in_r_bypass_regNext_13_2_stall_25;
  reg        [15:0]   io_in_r_bypass_regNext_13_3_data_25;
  reg                 io_in_r_bypass_regNext_13_3_load_store_25;
  reg                 io_in_r_bypass_regNext_13_3_df_is_ws_25;
  reg                 io_in_r_bypass_regNext_13_3_stall_25;
  reg        [15:0]   io_in_r_bypass_regNext_14_0_data_25;
  reg                 io_in_r_bypass_regNext_14_0_load_store_25;
  reg                 io_in_r_bypass_regNext_14_0_df_is_ws_25;
  reg                 io_in_r_bypass_regNext_14_0_stall_25;
  reg        [15:0]   io_in_r_bypass_regNext_14_1_data_25;
  reg                 io_in_r_bypass_regNext_14_1_load_store_25;
  reg                 io_in_r_bypass_regNext_14_1_df_is_ws_25;
  reg                 io_in_r_bypass_regNext_14_1_stall_25;
  reg        [15:0]   io_in_r_bypass_regNext_14_2_data_25;
  reg                 io_in_r_bypass_regNext_14_2_load_store_25;
  reg                 io_in_r_bypass_regNext_14_2_df_is_ws_25;
  reg                 io_in_r_bypass_regNext_14_2_stall_25;
  reg        [15:0]   io_in_r_bypass_regNext_14_3_data_25;
  reg                 io_in_r_bypass_regNext_14_3_load_store_25;
  reg                 io_in_r_bypass_regNext_14_3_df_is_ws_25;
  reg                 io_in_r_bypass_regNext_14_3_stall_25;
  reg        [15:0]   io_in_r_bypass_regNext_15_0_data_25;
  reg                 io_in_r_bypass_regNext_15_0_load_store_25;
  reg                 io_in_r_bypass_regNext_15_0_df_is_ws_25;
  reg                 io_in_r_bypass_regNext_15_0_stall_25;
  reg        [15:0]   io_in_r_bypass_regNext_15_1_data_25;
  reg                 io_in_r_bypass_regNext_15_1_load_store_25;
  reg                 io_in_r_bypass_regNext_15_1_df_is_ws_25;
  reg                 io_in_r_bypass_regNext_15_1_stall_25;
  reg        [15:0]   io_in_r_bypass_regNext_15_2_data_25;
  reg                 io_in_r_bypass_regNext_15_2_load_store_25;
  reg                 io_in_r_bypass_regNext_15_2_df_is_ws_25;
  reg                 io_in_r_bypass_regNext_15_2_stall_25;
  reg        [15:0]   io_in_r_bypass_regNext_15_3_data_25;
  reg                 io_in_r_bypass_regNext_15_3_load_store_25;
  reg                 io_in_r_bypass_regNext_15_3_df_is_ws_25;
  reg                 io_in_r_bypass_regNext_15_3_stall_25;
  reg        [15:0]   io_in_r_bypass_regNext_16_0_data_25;
  reg                 io_in_r_bypass_regNext_16_0_load_store_25;
  reg                 io_in_r_bypass_regNext_16_0_df_is_ws_25;
  reg                 io_in_r_bypass_regNext_16_0_stall_25;
  reg        [15:0]   io_in_r_bypass_regNext_16_1_data_25;
  reg                 io_in_r_bypass_regNext_16_1_load_store_25;
  reg                 io_in_r_bypass_regNext_16_1_df_is_ws_25;
  reg                 io_in_r_bypass_regNext_16_1_stall_25;
  reg        [15:0]   io_in_r_bypass_regNext_16_2_data_25;
  reg                 io_in_r_bypass_regNext_16_2_load_store_25;
  reg                 io_in_r_bypass_regNext_16_2_df_is_ws_25;
  reg                 io_in_r_bypass_regNext_16_2_stall_25;
  reg        [15:0]   io_in_r_bypass_regNext_16_3_data_25;
  reg                 io_in_r_bypass_regNext_16_3_load_store_25;
  reg                 io_in_r_bypass_regNext_16_3_df_is_ws_25;
  reg                 io_in_r_bypass_regNext_16_3_stall_25;
  reg        [15:0]   io_in_r_bypass_regNext_17_0_data_25;
  reg                 io_in_r_bypass_regNext_17_0_load_store_25;
  reg                 io_in_r_bypass_regNext_17_0_df_is_ws_25;
  reg                 io_in_r_bypass_regNext_17_0_stall_25;
  reg        [15:0]   io_in_r_bypass_regNext_17_1_data_25;
  reg                 io_in_r_bypass_regNext_17_1_load_store_25;
  reg                 io_in_r_bypass_regNext_17_1_df_is_ws_25;
  reg                 io_in_r_bypass_regNext_17_1_stall_25;
  reg        [15:0]   io_in_r_bypass_regNext_17_2_data_25;
  reg                 io_in_r_bypass_regNext_17_2_load_store_25;
  reg                 io_in_r_bypass_regNext_17_2_df_is_ws_25;
  reg                 io_in_r_bypass_regNext_17_2_stall_25;
  reg        [15:0]   io_in_r_bypass_regNext_17_3_data_25;
  reg                 io_in_r_bypass_regNext_17_3_load_store_25;
  reg                 io_in_r_bypass_regNext_17_3_df_is_ws_25;
  reg                 io_in_r_bypass_regNext_17_3_stall_25;
  reg        [15:0]   io_in_r_bypass_regNext_18_0_data_25;
  reg                 io_in_r_bypass_regNext_18_0_load_store_25;
  reg                 io_in_r_bypass_regNext_18_0_df_is_ws_25;
  reg                 io_in_r_bypass_regNext_18_0_stall_25;
  reg        [15:0]   io_in_r_bypass_regNext_18_1_data_25;
  reg                 io_in_r_bypass_regNext_18_1_load_store_25;
  reg                 io_in_r_bypass_regNext_18_1_df_is_ws_25;
  reg                 io_in_r_bypass_regNext_18_1_stall_25;
  reg        [15:0]   io_in_r_bypass_regNext_18_2_data_25;
  reg                 io_in_r_bypass_regNext_18_2_load_store_25;
  reg                 io_in_r_bypass_regNext_18_2_df_is_ws_25;
  reg                 io_in_r_bypass_regNext_18_2_stall_25;
  reg        [15:0]   io_in_r_bypass_regNext_18_3_data_25;
  reg                 io_in_r_bypass_regNext_18_3_load_store_25;
  reg                 io_in_r_bypass_regNext_18_3_df_is_ws_25;
  reg                 io_in_r_bypass_regNext_18_3_stall_25;
  reg        [15:0]   io_in_r_bypass_regNext_19_0_data_25;
  reg                 io_in_r_bypass_regNext_19_0_load_store_25;
  reg                 io_in_r_bypass_regNext_19_0_df_is_ws_25;
  reg                 io_in_r_bypass_regNext_19_0_stall_25;
  reg        [15:0]   io_in_r_bypass_regNext_19_1_data_25;
  reg                 io_in_r_bypass_regNext_19_1_load_store_25;
  reg                 io_in_r_bypass_regNext_19_1_df_is_ws_25;
  reg                 io_in_r_bypass_regNext_19_1_stall_25;
  reg        [15:0]   io_in_r_bypass_regNext_19_2_data_25;
  reg                 io_in_r_bypass_regNext_19_2_load_store_25;
  reg                 io_in_r_bypass_regNext_19_2_df_is_ws_25;
  reg                 io_in_r_bypass_regNext_19_2_stall_25;
  reg        [15:0]   io_in_r_bypass_regNext_19_3_data_25;
  reg                 io_in_r_bypass_regNext_19_3_load_store_25;
  reg                 io_in_r_bypass_regNext_19_3_df_is_ws_25;
  reg                 io_in_r_bypass_regNext_19_3_stall_25;
  reg        [15:0]   io_in_r_bypass_regNext_20_0_data_25;
  reg                 io_in_r_bypass_regNext_20_0_load_store_25;
  reg                 io_in_r_bypass_regNext_20_0_df_is_ws_25;
  reg                 io_in_r_bypass_regNext_20_0_stall_25;
  reg        [15:0]   io_in_r_bypass_regNext_20_1_data_25;
  reg                 io_in_r_bypass_regNext_20_1_load_store_25;
  reg                 io_in_r_bypass_regNext_20_1_df_is_ws_25;
  reg                 io_in_r_bypass_regNext_20_1_stall_25;
  reg        [15:0]   io_in_r_bypass_regNext_20_2_data_25;
  reg                 io_in_r_bypass_regNext_20_2_load_store_25;
  reg                 io_in_r_bypass_regNext_20_2_df_is_ws_25;
  reg                 io_in_r_bypass_regNext_20_2_stall_25;
  reg        [15:0]   io_in_r_bypass_regNext_20_3_data_25;
  reg                 io_in_r_bypass_regNext_20_3_load_store_25;
  reg                 io_in_r_bypass_regNext_20_3_df_is_ws_25;
  reg                 io_in_r_bypass_regNext_20_3_stall_25;
  reg        [15:0]   io_in_r_bypass_regNext_21_0_data_25;
  reg                 io_in_r_bypass_regNext_21_0_load_store_25;
  reg                 io_in_r_bypass_regNext_21_0_df_is_ws_25;
  reg                 io_in_r_bypass_regNext_21_0_stall_25;
  reg        [15:0]   io_in_r_bypass_regNext_21_1_data_25;
  reg                 io_in_r_bypass_regNext_21_1_load_store_25;
  reg                 io_in_r_bypass_regNext_21_1_df_is_ws_25;
  reg                 io_in_r_bypass_regNext_21_1_stall_25;
  reg        [15:0]   io_in_r_bypass_regNext_21_2_data_25;
  reg                 io_in_r_bypass_regNext_21_2_load_store_25;
  reg                 io_in_r_bypass_regNext_21_2_df_is_ws_25;
  reg                 io_in_r_bypass_regNext_21_2_stall_25;
  reg        [15:0]   io_in_r_bypass_regNext_21_3_data_25;
  reg                 io_in_r_bypass_regNext_21_3_load_store_25;
  reg                 io_in_r_bypass_regNext_21_3_df_is_ws_25;
  reg                 io_in_r_bypass_regNext_21_3_stall_25;
  reg        [15:0]   io_in_r_bypass_regNext_22_0_data_25;
  reg                 io_in_r_bypass_regNext_22_0_load_store_25;
  reg                 io_in_r_bypass_regNext_22_0_df_is_ws_25;
  reg                 io_in_r_bypass_regNext_22_0_stall_25;
  reg        [15:0]   io_in_r_bypass_regNext_22_1_data_25;
  reg                 io_in_r_bypass_regNext_22_1_load_store_25;
  reg                 io_in_r_bypass_regNext_22_1_df_is_ws_25;
  reg                 io_in_r_bypass_regNext_22_1_stall_25;
  reg        [15:0]   io_in_r_bypass_regNext_22_2_data_25;
  reg                 io_in_r_bypass_regNext_22_2_load_store_25;
  reg                 io_in_r_bypass_regNext_22_2_df_is_ws_25;
  reg                 io_in_r_bypass_regNext_22_2_stall_25;
  reg        [15:0]   io_in_r_bypass_regNext_22_3_data_25;
  reg                 io_in_r_bypass_regNext_22_3_load_store_25;
  reg                 io_in_r_bypass_regNext_22_3_df_is_ws_25;
  reg                 io_in_r_bypass_regNext_22_3_stall_25;
  reg        [15:0]   io_in_r_bypass_regNext_23_0_data_25;
  reg                 io_in_r_bypass_regNext_23_0_load_store_25;
  reg                 io_in_r_bypass_regNext_23_0_df_is_ws_25;
  reg                 io_in_r_bypass_regNext_23_0_stall_25;
  reg        [15:0]   io_in_r_bypass_regNext_23_1_data_25;
  reg                 io_in_r_bypass_regNext_23_1_load_store_25;
  reg                 io_in_r_bypass_regNext_23_1_df_is_ws_25;
  reg                 io_in_r_bypass_regNext_23_1_stall_25;
  reg        [15:0]   io_in_r_bypass_regNext_23_2_data_25;
  reg                 io_in_r_bypass_regNext_23_2_load_store_25;
  reg                 io_in_r_bypass_regNext_23_2_df_is_ws_25;
  reg                 io_in_r_bypass_regNext_23_2_stall_25;
  reg        [15:0]   io_in_r_bypass_regNext_23_3_data_25;
  reg                 io_in_r_bypass_regNext_23_3_load_store_25;
  reg                 io_in_r_bypass_regNext_23_3_df_is_ws_25;
  reg                 io_in_r_bypass_regNext_23_3_stall_25;
  reg        [15:0]   io_in_r_bypass_regNext_24_0_data_25;
  reg                 io_in_r_bypass_regNext_24_0_load_store_25;
  reg                 io_in_r_bypass_regNext_24_0_df_is_ws_25;
  reg                 io_in_r_bypass_regNext_24_0_stall_25;
  reg        [15:0]   io_in_r_bypass_regNext_24_1_data_25;
  reg                 io_in_r_bypass_regNext_24_1_load_store_25;
  reg                 io_in_r_bypass_regNext_24_1_df_is_ws_25;
  reg                 io_in_r_bypass_regNext_24_1_stall_25;
  reg        [15:0]   io_in_r_bypass_regNext_24_2_data_25;
  reg                 io_in_r_bypass_regNext_24_2_load_store_25;
  reg                 io_in_r_bypass_regNext_24_2_df_is_ws_25;
  reg                 io_in_r_bypass_regNext_24_2_stall_25;
  reg        [15:0]   io_in_r_bypass_regNext_24_3_data_25;
  reg                 io_in_r_bypass_regNext_24_3_load_store_25;
  reg                 io_in_r_bypass_regNext_24_3_df_is_ws_25;
  reg                 io_in_r_bypass_regNext_24_3_stall_25;
  reg        [15:0]   io_in_r_bypass_regNext_25_0_data_25;
  reg                 io_in_r_bypass_regNext_25_0_load_store_25;
  reg                 io_in_r_bypass_regNext_25_0_df_is_ws_25;
  reg                 io_in_r_bypass_regNext_25_0_stall_25;
  reg        [15:0]   io_in_r_bypass_regNext_25_1_data_25;
  reg                 io_in_r_bypass_regNext_25_1_load_store_25;
  reg                 io_in_r_bypass_regNext_25_1_df_is_ws_25;
  reg                 io_in_r_bypass_regNext_25_1_stall_25;
  reg        [15:0]   io_in_r_bypass_regNext_25_2_data_25;
  reg                 io_in_r_bypass_regNext_25_2_load_store_25;
  reg                 io_in_r_bypass_regNext_25_2_df_is_ws_25;
  reg                 io_in_r_bypass_regNext_25_2_stall_25;
  reg        [15:0]   io_in_r_bypass_regNext_25_3_data_25;
  reg                 io_in_r_bypass_regNext_25_3_load_store_25;
  reg                 io_in_r_bypass_regNext_25_3_df_is_ws_25;
  reg                 io_in_r_bypass_regNext_25_3_stall_25;
  reg        [15:0]   io_in_r_bypass_regNext_26_0_data_25;
  reg                 io_in_r_bypass_regNext_26_0_load_store_25;
  reg                 io_in_r_bypass_regNext_26_0_df_is_ws_25;
  reg                 io_in_r_bypass_regNext_26_0_stall_25;
  reg        [15:0]   io_in_r_bypass_regNext_26_1_data_25;
  reg                 io_in_r_bypass_regNext_26_1_load_store_25;
  reg                 io_in_r_bypass_regNext_26_1_df_is_ws_25;
  reg                 io_in_r_bypass_regNext_26_1_stall_25;
  reg        [15:0]   io_in_r_bypass_regNext_26_2_data_25;
  reg                 io_in_r_bypass_regNext_26_2_load_store_25;
  reg                 io_in_r_bypass_regNext_26_2_df_is_ws_25;
  reg                 io_in_r_bypass_regNext_26_2_stall_25;
  reg        [15:0]   io_in_r_bypass_regNext_26_3_data_25;
  reg                 io_in_r_bypass_regNext_26_3_load_store_25;
  reg                 io_in_r_bypass_regNext_26_3_df_is_ws_25;
  reg                 io_in_r_bypass_regNext_26_3_stall_25;
  reg        [15:0]   io_in_r_bypass_regNext_27_0_data_25;
  reg                 io_in_r_bypass_regNext_27_0_load_store_25;
  reg                 io_in_r_bypass_regNext_27_0_df_is_ws_25;
  reg                 io_in_r_bypass_regNext_27_0_stall_25;
  reg        [15:0]   io_in_r_bypass_regNext_27_1_data_25;
  reg                 io_in_r_bypass_regNext_27_1_load_store_25;
  reg                 io_in_r_bypass_regNext_27_1_df_is_ws_25;
  reg                 io_in_r_bypass_regNext_27_1_stall_25;
  reg        [15:0]   io_in_r_bypass_regNext_27_2_data_25;
  reg                 io_in_r_bypass_regNext_27_2_load_store_25;
  reg                 io_in_r_bypass_regNext_27_2_df_is_ws_25;
  reg                 io_in_r_bypass_regNext_27_2_stall_25;
  reg        [15:0]   io_in_r_bypass_regNext_27_3_data_25;
  reg                 io_in_r_bypass_regNext_27_3_load_store_25;
  reg                 io_in_r_bypass_regNext_27_3_df_is_ws_25;
  reg                 io_in_r_bypass_regNext_27_3_stall_25;
  reg        [15:0]   io_in_r_bypass_regNext_28_0_data_25;
  reg                 io_in_r_bypass_regNext_28_0_load_store_25;
  reg                 io_in_r_bypass_regNext_28_0_df_is_ws_25;
  reg                 io_in_r_bypass_regNext_28_0_stall_25;
  reg        [15:0]   io_in_r_bypass_regNext_28_1_data_25;
  reg                 io_in_r_bypass_regNext_28_1_load_store_25;
  reg                 io_in_r_bypass_regNext_28_1_df_is_ws_25;
  reg                 io_in_r_bypass_regNext_28_1_stall_25;
  reg        [15:0]   io_in_r_bypass_regNext_28_2_data_25;
  reg                 io_in_r_bypass_regNext_28_2_load_store_25;
  reg                 io_in_r_bypass_regNext_28_2_df_is_ws_25;
  reg                 io_in_r_bypass_regNext_28_2_stall_25;
  reg        [15:0]   io_in_r_bypass_regNext_28_3_data_25;
  reg                 io_in_r_bypass_regNext_28_3_load_store_25;
  reg                 io_in_r_bypass_regNext_28_3_df_is_ws_25;
  reg                 io_in_r_bypass_regNext_28_3_stall_25;
  reg        [15:0]   io_in_r_bypass_regNext_29_0_data_25;
  reg                 io_in_r_bypass_regNext_29_0_load_store_25;
  reg                 io_in_r_bypass_regNext_29_0_df_is_ws_25;
  reg                 io_in_r_bypass_regNext_29_0_stall_25;
  reg        [15:0]   io_in_r_bypass_regNext_29_1_data_25;
  reg                 io_in_r_bypass_regNext_29_1_load_store_25;
  reg                 io_in_r_bypass_regNext_29_1_df_is_ws_25;
  reg                 io_in_r_bypass_regNext_29_1_stall_25;
  reg        [15:0]   io_in_r_bypass_regNext_29_2_data_25;
  reg                 io_in_r_bypass_regNext_29_2_load_store_25;
  reg                 io_in_r_bypass_regNext_29_2_df_is_ws_25;
  reg                 io_in_r_bypass_regNext_29_2_stall_25;
  reg        [15:0]   io_in_r_bypass_regNext_29_3_data_25;
  reg                 io_in_r_bypass_regNext_29_3_load_store_25;
  reg                 io_in_r_bypass_regNext_29_3_df_is_ws_25;
  reg                 io_in_r_bypass_regNext_29_3_stall_25;
  reg        [15:0]   io_in_r_bypass_regNext_30_0_data_25;
  reg                 io_in_r_bypass_regNext_30_0_load_store_25;
  reg                 io_in_r_bypass_regNext_30_0_df_is_ws_25;
  reg                 io_in_r_bypass_regNext_30_0_stall_25;
  reg        [15:0]   io_in_r_bypass_regNext_30_1_data_25;
  reg                 io_in_r_bypass_regNext_30_1_load_store_25;
  reg                 io_in_r_bypass_regNext_30_1_df_is_ws_25;
  reg                 io_in_r_bypass_regNext_30_1_stall_25;
  reg        [15:0]   io_in_r_bypass_regNext_30_2_data_25;
  reg                 io_in_r_bypass_regNext_30_2_load_store_25;
  reg                 io_in_r_bypass_regNext_30_2_df_is_ws_25;
  reg                 io_in_r_bypass_regNext_30_2_stall_25;
  reg        [15:0]   io_in_r_bypass_regNext_30_3_data_25;
  reg                 io_in_r_bypass_regNext_30_3_load_store_25;
  reg                 io_in_r_bypass_regNext_30_3_df_is_ws_25;
  reg                 io_in_r_bypass_regNext_30_3_stall_25;
  reg        [15:0]   io_in_r_bypass_regNext_31_0_data_25;
  reg                 io_in_r_bypass_regNext_31_0_load_store_25;
  reg                 io_in_r_bypass_regNext_31_0_df_is_ws_25;
  reg                 io_in_r_bypass_regNext_31_0_stall_25;
  reg        [15:0]   io_in_r_bypass_regNext_31_1_data_25;
  reg                 io_in_r_bypass_regNext_31_1_load_store_25;
  reg                 io_in_r_bypass_regNext_31_1_df_is_ws_25;
  reg                 io_in_r_bypass_regNext_31_1_stall_25;
  reg        [15:0]   io_in_r_bypass_regNext_31_2_data_25;
  reg                 io_in_r_bypass_regNext_31_2_load_store_25;
  reg                 io_in_r_bypass_regNext_31_2_df_is_ws_25;
  reg                 io_in_r_bypass_regNext_31_2_stall_25;
  reg        [15:0]   io_in_r_bypass_regNext_31_3_data_25;
  reg                 io_in_r_bypass_regNext_31_3_load_store_25;
  reg                 io_in_r_bypass_regNext_31_3_df_is_ws_25;
  reg                 io_in_r_bypass_regNext_31_3_stall_25;
  reg        [15:0]   io_in_r_bypass_regNext_0_0_data_26;
  reg                 io_in_r_bypass_regNext_0_0_load_store_26;
  reg                 io_in_r_bypass_regNext_0_0_df_is_ws_26;
  reg                 io_in_r_bypass_regNext_0_0_stall_26;
  reg        [15:0]   io_in_r_bypass_regNext_0_1_data_26;
  reg                 io_in_r_bypass_regNext_0_1_load_store_26;
  reg                 io_in_r_bypass_regNext_0_1_df_is_ws_26;
  reg                 io_in_r_bypass_regNext_0_1_stall_26;
  reg        [15:0]   io_in_r_bypass_regNext_0_2_data_26;
  reg                 io_in_r_bypass_regNext_0_2_load_store_26;
  reg                 io_in_r_bypass_regNext_0_2_df_is_ws_26;
  reg                 io_in_r_bypass_regNext_0_2_stall_26;
  reg        [15:0]   io_in_r_bypass_regNext_0_3_data_26;
  reg                 io_in_r_bypass_regNext_0_3_load_store_26;
  reg                 io_in_r_bypass_regNext_0_3_df_is_ws_26;
  reg                 io_in_r_bypass_regNext_0_3_stall_26;
  reg        [15:0]   io_in_r_bypass_regNext_1_0_data_26;
  reg                 io_in_r_bypass_regNext_1_0_load_store_26;
  reg                 io_in_r_bypass_regNext_1_0_df_is_ws_26;
  reg                 io_in_r_bypass_regNext_1_0_stall_26;
  reg        [15:0]   io_in_r_bypass_regNext_1_1_data_26;
  reg                 io_in_r_bypass_regNext_1_1_load_store_26;
  reg                 io_in_r_bypass_regNext_1_1_df_is_ws_26;
  reg                 io_in_r_bypass_regNext_1_1_stall_26;
  reg        [15:0]   io_in_r_bypass_regNext_1_2_data_26;
  reg                 io_in_r_bypass_regNext_1_2_load_store_26;
  reg                 io_in_r_bypass_regNext_1_2_df_is_ws_26;
  reg                 io_in_r_bypass_regNext_1_2_stall_26;
  reg        [15:0]   io_in_r_bypass_regNext_1_3_data_26;
  reg                 io_in_r_bypass_regNext_1_3_load_store_26;
  reg                 io_in_r_bypass_regNext_1_3_df_is_ws_26;
  reg                 io_in_r_bypass_regNext_1_3_stall_26;
  reg        [15:0]   io_in_r_bypass_regNext_2_0_data_26;
  reg                 io_in_r_bypass_regNext_2_0_load_store_26;
  reg                 io_in_r_bypass_regNext_2_0_df_is_ws_26;
  reg                 io_in_r_bypass_regNext_2_0_stall_26;
  reg        [15:0]   io_in_r_bypass_regNext_2_1_data_26;
  reg                 io_in_r_bypass_regNext_2_1_load_store_26;
  reg                 io_in_r_bypass_regNext_2_1_df_is_ws_26;
  reg                 io_in_r_bypass_regNext_2_1_stall_26;
  reg        [15:0]   io_in_r_bypass_regNext_2_2_data_26;
  reg                 io_in_r_bypass_regNext_2_2_load_store_26;
  reg                 io_in_r_bypass_regNext_2_2_df_is_ws_26;
  reg                 io_in_r_bypass_regNext_2_2_stall_26;
  reg        [15:0]   io_in_r_bypass_regNext_2_3_data_26;
  reg                 io_in_r_bypass_regNext_2_3_load_store_26;
  reg                 io_in_r_bypass_regNext_2_3_df_is_ws_26;
  reg                 io_in_r_bypass_regNext_2_3_stall_26;
  reg        [15:0]   io_in_r_bypass_regNext_3_0_data_26;
  reg                 io_in_r_bypass_regNext_3_0_load_store_26;
  reg                 io_in_r_bypass_regNext_3_0_df_is_ws_26;
  reg                 io_in_r_bypass_regNext_3_0_stall_26;
  reg        [15:0]   io_in_r_bypass_regNext_3_1_data_26;
  reg                 io_in_r_bypass_regNext_3_1_load_store_26;
  reg                 io_in_r_bypass_regNext_3_1_df_is_ws_26;
  reg                 io_in_r_bypass_regNext_3_1_stall_26;
  reg        [15:0]   io_in_r_bypass_regNext_3_2_data_26;
  reg                 io_in_r_bypass_regNext_3_2_load_store_26;
  reg                 io_in_r_bypass_regNext_3_2_df_is_ws_26;
  reg                 io_in_r_bypass_regNext_3_2_stall_26;
  reg        [15:0]   io_in_r_bypass_regNext_3_3_data_26;
  reg                 io_in_r_bypass_regNext_3_3_load_store_26;
  reg                 io_in_r_bypass_regNext_3_3_df_is_ws_26;
  reg                 io_in_r_bypass_regNext_3_3_stall_26;
  reg        [15:0]   io_in_r_bypass_regNext_4_0_data_26;
  reg                 io_in_r_bypass_regNext_4_0_load_store_26;
  reg                 io_in_r_bypass_regNext_4_0_df_is_ws_26;
  reg                 io_in_r_bypass_regNext_4_0_stall_26;
  reg        [15:0]   io_in_r_bypass_regNext_4_1_data_26;
  reg                 io_in_r_bypass_regNext_4_1_load_store_26;
  reg                 io_in_r_bypass_regNext_4_1_df_is_ws_26;
  reg                 io_in_r_bypass_regNext_4_1_stall_26;
  reg        [15:0]   io_in_r_bypass_regNext_4_2_data_26;
  reg                 io_in_r_bypass_regNext_4_2_load_store_26;
  reg                 io_in_r_bypass_regNext_4_2_df_is_ws_26;
  reg                 io_in_r_bypass_regNext_4_2_stall_26;
  reg        [15:0]   io_in_r_bypass_regNext_4_3_data_26;
  reg                 io_in_r_bypass_regNext_4_3_load_store_26;
  reg                 io_in_r_bypass_regNext_4_3_df_is_ws_26;
  reg                 io_in_r_bypass_regNext_4_3_stall_26;
  reg        [15:0]   io_in_r_bypass_regNext_5_0_data_26;
  reg                 io_in_r_bypass_regNext_5_0_load_store_26;
  reg                 io_in_r_bypass_regNext_5_0_df_is_ws_26;
  reg                 io_in_r_bypass_regNext_5_0_stall_26;
  reg        [15:0]   io_in_r_bypass_regNext_5_1_data_26;
  reg                 io_in_r_bypass_regNext_5_1_load_store_26;
  reg                 io_in_r_bypass_regNext_5_1_df_is_ws_26;
  reg                 io_in_r_bypass_regNext_5_1_stall_26;
  reg        [15:0]   io_in_r_bypass_regNext_5_2_data_26;
  reg                 io_in_r_bypass_regNext_5_2_load_store_26;
  reg                 io_in_r_bypass_regNext_5_2_df_is_ws_26;
  reg                 io_in_r_bypass_regNext_5_2_stall_26;
  reg        [15:0]   io_in_r_bypass_regNext_5_3_data_26;
  reg                 io_in_r_bypass_regNext_5_3_load_store_26;
  reg                 io_in_r_bypass_regNext_5_3_df_is_ws_26;
  reg                 io_in_r_bypass_regNext_5_3_stall_26;
  reg        [15:0]   io_in_r_bypass_regNext_6_0_data_26;
  reg                 io_in_r_bypass_regNext_6_0_load_store_26;
  reg                 io_in_r_bypass_regNext_6_0_df_is_ws_26;
  reg                 io_in_r_bypass_regNext_6_0_stall_26;
  reg        [15:0]   io_in_r_bypass_regNext_6_1_data_26;
  reg                 io_in_r_bypass_regNext_6_1_load_store_26;
  reg                 io_in_r_bypass_regNext_6_1_df_is_ws_26;
  reg                 io_in_r_bypass_regNext_6_1_stall_26;
  reg        [15:0]   io_in_r_bypass_regNext_6_2_data_26;
  reg                 io_in_r_bypass_regNext_6_2_load_store_26;
  reg                 io_in_r_bypass_regNext_6_2_df_is_ws_26;
  reg                 io_in_r_bypass_regNext_6_2_stall_26;
  reg        [15:0]   io_in_r_bypass_regNext_6_3_data_26;
  reg                 io_in_r_bypass_regNext_6_3_load_store_26;
  reg                 io_in_r_bypass_regNext_6_3_df_is_ws_26;
  reg                 io_in_r_bypass_regNext_6_3_stall_26;
  reg        [15:0]   io_in_r_bypass_regNext_7_0_data_26;
  reg                 io_in_r_bypass_regNext_7_0_load_store_26;
  reg                 io_in_r_bypass_regNext_7_0_df_is_ws_26;
  reg                 io_in_r_bypass_regNext_7_0_stall_26;
  reg        [15:0]   io_in_r_bypass_regNext_7_1_data_26;
  reg                 io_in_r_bypass_regNext_7_1_load_store_26;
  reg                 io_in_r_bypass_regNext_7_1_df_is_ws_26;
  reg                 io_in_r_bypass_regNext_7_1_stall_26;
  reg        [15:0]   io_in_r_bypass_regNext_7_2_data_26;
  reg                 io_in_r_bypass_regNext_7_2_load_store_26;
  reg                 io_in_r_bypass_regNext_7_2_df_is_ws_26;
  reg                 io_in_r_bypass_regNext_7_2_stall_26;
  reg        [15:0]   io_in_r_bypass_regNext_7_3_data_26;
  reg                 io_in_r_bypass_regNext_7_3_load_store_26;
  reg                 io_in_r_bypass_regNext_7_3_df_is_ws_26;
  reg                 io_in_r_bypass_regNext_7_3_stall_26;
  reg        [15:0]   io_in_r_bypass_regNext_8_0_data_26;
  reg                 io_in_r_bypass_regNext_8_0_load_store_26;
  reg                 io_in_r_bypass_regNext_8_0_df_is_ws_26;
  reg                 io_in_r_bypass_regNext_8_0_stall_26;
  reg        [15:0]   io_in_r_bypass_regNext_8_1_data_26;
  reg                 io_in_r_bypass_regNext_8_1_load_store_26;
  reg                 io_in_r_bypass_regNext_8_1_df_is_ws_26;
  reg                 io_in_r_bypass_regNext_8_1_stall_26;
  reg        [15:0]   io_in_r_bypass_regNext_8_2_data_26;
  reg                 io_in_r_bypass_regNext_8_2_load_store_26;
  reg                 io_in_r_bypass_regNext_8_2_df_is_ws_26;
  reg                 io_in_r_bypass_regNext_8_2_stall_26;
  reg        [15:0]   io_in_r_bypass_regNext_8_3_data_26;
  reg                 io_in_r_bypass_regNext_8_3_load_store_26;
  reg                 io_in_r_bypass_regNext_8_3_df_is_ws_26;
  reg                 io_in_r_bypass_regNext_8_3_stall_26;
  reg        [15:0]   io_in_r_bypass_regNext_9_0_data_26;
  reg                 io_in_r_bypass_regNext_9_0_load_store_26;
  reg                 io_in_r_bypass_regNext_9_0_df_is_ws_26;
  reg                 io_in_r_bypass_regNext_9_0_stall_26;
  reg        [15:0]   io_in_r_bypass_regNext_9_1_data_26;
  reg                 io_in_r_bypass_regNext_9_1_load_store_26;
  reg                 io_in_r_bypass_regNext_9_1_df_is_ws_26;
  reg                 io_in_r_bypass_regNext_9_1_stall_26;
  reg        [15:0]   io_in_r_bypass_regNext_9_2_data_26;
  reg                 io_in_r_bypass_regNext_9_2_load_store_26;
  reg                 io_in_r_bypass_regNext_9_2_df_is_ws_26;
  reg                 io_in_r_bypass_regNext_9_2_stall_26;
  reg        [15:0]   io_in_r_bypass_regNext_9_3_data_26;
  reg                 io_in_r_bypass_regNext_9_3_load_store_26;
  reg                 io_in_r_bypass_regNext_9_3_df_is_ws_26;
  reg                 io_in_r_bypass_regNext_9_3_stall_26;
  reg        [15:0]   io_in_r_bypass_regNext_10_0_data_26;
  reg                 io_in_r_bypass_regNext_10_0_load_store_26;
  reg                 io_in_r_bypass_regNext_10_0_df_is_ws_26;
  reg                 io_in_r_bypass_regNext_10_0_stall_26;
  reg        [15:0]   io_in_r_bypass_regNext_10_1_data_26;
  reg                 io_in_r_bypass_regNext_10_1_load_store_26;
  reg                 io_in_r_bypass_regNext_10_1_df_is_ws_26;
  reg                 io_in_r_bypass_regNext_10_1_stall_26;
  reg        [15:0]   io_in_r_bypass_regNext_10_2_data_26;
  reg                 io_in_r_bypass_regNext_10_2_load_store_26;
  reg                 io_in_r_bypass_regNext_10_2_df_is_ws_26;
  reg                 io_in_r_bypass_regNext_10_2_stall_26;
  reg        [15:0]   io_in_r_bypass_regNext_10_3_data_26;
  reg                 io_in_r_bypass_regNext_10_3_load_store_26;
  reg                 io_in_r_bypass_regNext_10_3_df_is_ws_26;
  reg                 io_in_r_bypass_regNext_10_3_stall_26;
  reg        [15:0]   io_in_r_bypass_regNext_11_0_data_26;
  reg                 io_in_r_bypass_regNext_11_0_load_store_26;
  reg                 io_in_r_bypass_regNext_11_0_df_is_ws_26;
  reg                 io_in_r_bypass_regNext_11_0_stall_26;
  reg        [15:0]   io_in_r_bypass_regNext_11_1_data_26;
  reg                 io_in_r_bypass_regNext_11_1_load_store_26;
  reg                 io_in_r_bypass_regNext_11_1_df_is_ws_26;
  reg                 io_in_r_bypass_regNext_11_1_stall_26;
  reg        [15:0]   io_in_r_bypass_regNext_11_2_data_26;
  reg                 io_in_r_bypass_regNext_11_2_load_store_26;
  reg                 io_in_r_bypass_regNext_11_2_df_is_ws_26;
  reg                 io_in_r_bypass_regNext_11_2_stall_26;
  reg        [15:0]   io_in_r_bypass_regNext_11_3_data_26;
  reg                 io_in_r_bypass_regNext_11_3_load_store_26;
  reg                 io_in_r_bypass_regNext_11_3_df_is_ws_26;
  reg                 io_in_r_bypass_regNext_11_3_stall_26;
  reg        [15:0]   io_in_r_bypass_regNext_12_0_data_26;
  reg                 io_in_r_bypass_regNext_12_0_load_store_26;
  reg                 io_in_r_bypass_regNext_12_0_df_is_ws_26;
  reg                 io_in_r_bypass_regNext_12_0_stall_26;
  reg        [15:0]   io_in_r_bypass_regNext_12_1_data_26;
  reg                 io_in_r_bypass_regNext_12_1_load_store_26;
  reg                 io_in_r_bypass_regNext_12_1_df_is_ws_26;
  reg                 io_in_r_bypass_regNext_12_1_stall_26;
  reg        [15:0]   io_in_r_bypass_regNext_12_2_data_26;
  reg                 io_in_r_bypass_regNext_12_2_load_store_26;
  reg                 io_in_r_bypass_regNext_12_2_df_is_ws_26;
  reg                 io_in_r_bypass_regNext_12_2_stall_26;
  reg        [15:0]   io_in_r_bypass_regNext_12_3_data_26;
  reg                 io_in_r_bypass_regNext_12_3_load_store_26;
  reg                 io_in_r_bypass_regNext_12_3_df_is_ws_26;
  reg                 io_in_r_bypass_regNext_12_3_stall_26;
  reg        [15:0]   io_in_r_bypass_regNext_13_0_data_26;
  reg                 io_in_r_bypass_regNext_13_0_load_store_26;
  reg                 io_in_r_bypass_regNext_13_0_df_is_ws_26;
  reg                 io_in_r_bypass_regNext_13_0_stall_26;
  reg        [15:0]   io_in_r_bypass_regNext_13_1_data_26;
  reg                 io_in_r_bypass_regNext_13_1_load_store_26;
  reg                 io_in_r_bypass_regNext_13_1_df_is_ws_26;
  reg                 io_in_r_bypass_regNext_13_1_stall_26;
  reg        [15:0]   io_in_r_bypass_regNext_13_2_data_26;
  reg                 io_in_r_bypass_regNext_13_2_load_store_26;
  reg                 io_in_r_bypass_regNext_13_2_df_is_ws_26;
  reg                 io_in_r_bypass_regNext_13_2_stall_26;
  reg        [15:0]   io_in_r_bypass_regNext_13_3_data_26;
  reg                 io_in_r_bypass_regNext_13_3_load_store_26;
  reg                 io_in_r_bypass_regNext_13_3_df_is_ws_26;
  reg                 io_in_r_bypass_regNext_13_3_stall_26;
  reg        [15:0]   io_in_r_bypass_regNext_14_0_data_26;
  reg                 io_in_r_bypass_regNext_14_0_load_store_26;
  reg                 io_in_r_bypass_regNext_14_0_df_is_ws_26;
  reg                 io_in_r_bypass_regNext_14_0_stall_26;
  reg        [15:0]   io_in_r_bypass_regNext_14_1_data_26;
  reg                 io_in_r_bypass_regNext_14_1_load_store_26;
  reg                 io_in_r_bypass_regNext_14_1_df_is_ws_26;
  reg                 io_in_r_bypass_regNext_14_1_stall_26;
  reg        [15:0]   io_in_r_bypass_regNext_14_2_data_26;
  reg                 io_in_r_bypass_regNext_14_2_load_store_26;
  reg                 io_in_r_bypass_regNext_14_2_df_is_ws_26;
  reg                 io_in_r_bypass_regNext_14_2_stall_26;
  reg        [15:0]   io_in_r_bypass_regNext_14_3_data_26;
  reg                 io_in_r_bypass_regNext_14_3_load_store_26;
  reg                 io_in_r_bypass_regNext_14_3_df_is_ws_26;
  reg                 io_in_r_bypass_regNext_14_3_stall_26;
  reg        [15:0]   io_in_r_bypass_regNext_15_0_data_26;
  reg                 io_in_r_bypass_regNext_15_0_load_store_26;
  reg                 io_in_r_bypass_regNext_15_0_df_is_ws_26;
  reg                 io_in_r_bypass_regNext_15_0_stall_26;
  reg        [15:0]   io_in_r_bypass_regNext_15_1_data_26;
  reg                 io_in_r_bypass_regNext_15_1_load_store_26;
  reg                 io_in_r_bypass_regNext_15_1_df_is_ws_26;
  reg                 io_in_r_bypass_regNext_15_1_stall_26;
  reg        [15:0]   io_in_r_bypass_regNext_15_2_data_26;
  reg                 io_in_r_bypass_regNext_15_2_load_store_26;
  reg                 io_in_r_bypass_regNext_15_2_df_is_ws_26;
  reg                 io_in_r_bypass_regNext_15_2_stall_26;
  reg        [15:0]   io_in_r_bypass_regNext_15_3_data_26;
  reg                 io_in_r_bypass_regNext_15_3_load_store_26;
  reg                 io_in_r_bypass_regNext_15_3_df_is_ws_26;
  reg                 io_in_r_bypass_regNext_15_3_stall_26;
  reg        [15:0]   io_in_r_bypass_regNext_16_0_data_26;
  reg                 io_in_r_bypass_regNext_16_0_load_store_26;
  reg                 io_in_r_bypass_regNext_16_0_df_is_ws_26;
  reg                 io_in_r_bypass_regNext_16_0_stall_26;
  reg        [15:0]   io_in_r_bypass_regNext_16_1_data_26;
  reg                 io_in_r_bypass_regNext_16_1_load_store_26;
  reg                 io_in_r_bypass_regNext_16_1_df_is_ws_26;
  reg                 io_in_r_bypass_regNext_16_1_stall_26;
  reg        [15:0]   io_in_r_bypass_regNext_16_2_data_26;
  reg                 io_in_r_bypass_regNext_16_2_load_store_26;
  reg                 io_in_r_bypass_regNext_16_2_df_is_ws_26;
  reg                 io_in_r_bypass_regNext_16_2_stall_26;
  reg        [15:0]   io_in_r_bypass_regNext_16_3_data_26;
  reg                 io_in_r_bypass_regNext_16_3_load_store_26;
  reg                 io_in_r_bypass_regNext_16_3_df_is_ws_26;
  reg                 io_in_r_bypass_regNext_16_3_stall_26;
  reg        [15:0]   io_in_r_bypass_regNext_17_0_data_26;
  reg                 io_in_r_bypass_regNext_17_0_load_store_26;
  reg                 io_in_r_bypass_regNext_17_0_df_is_ws_26;
  reg                 io_in_r_bypass_regNext_17_0_stall_26;
  reg        [15:0]   io_in_r_bypass_regNext_17_1_data_26;
  reg                 io_in_r_bypass_regNext_17_1_load_store_26;
  reg                 io_in_r_bypass_regNext_17_1_df_is_ws_26;
  reg                 io_in_r_bypass_regNext_17_1_stall_26;
  reg        [15:0]   io_in_r_bypass_regNext_17_2_data_26;
  reg                 io_in_r_bypass_regNext_17_2_load_store_26;
  reg                 io_in_r_bypass_regNext_17_2_df_is_ws_26;
  reg                 io_in_r_bypass_regNext_17_2_stall_26;
  reg        [15:0]   io_in_r_bypass_regNext_17_3_data_26;
  reg                 io_in_r_bypass_regNext_17_3_load_store_26;
  reg                 io_in_r_bypass_regNext_17_3_df_is_ws_26;
  reg                 io_in_r_bypass_regNext_17_3_stall_26;
  reg        [15:0]   io_in_r_bypass_regNext_18_0_data_26;
  reg                 io_in_r_bypass_regNext_18_0_load_store_26;
  reg                 io_in_r_bypass_regNext_18_0_df_is_ws_26;
  reg                 io_in_r_bypass_regNext_18_0_stall_26;
  reg        [15:0]   io_in_r_bypass_regNext_18_1_data_26;
  reg                 io_in_r_bypass_regNext_18_1_load_store_26;
  reg                 io_in_r_bypass_regNext_18_1_df_is_ws_26;
  reg                 io_in_r_bypass_regNext_18_1_stall_26;
  reg        [15:0]   io_in_r_bypass_regNext_18_2_data_26;
  reg                 io_in_r_bypass_regNext_18_2_load_store_26;
  reg                 io_in_r_bypass_regNext_18_2_df_is_ws_26;
  reg                 io_in_r_bypass_regNext_18_2_stall_26;
  reg        [15:0]   io_in_r_bypass_regNext_18_3_data_26;
  reg                 io_in_r_bypass_regNext_18_3_load_store_26;
  reg                 io_in_r_bypass_regNext_18_3_df_is_ws_26;
  reg                 io_in_r_bypass_regNext_18_3_stall_26;
  reg        [15:0]   io_in_r_bypass_regNext_19_0_data_26;
  reg                 io_in_r_bypass_regNext_19_0_load_store_26;
  reg                 io_in_r_bypass_regNext_19_0_df_is_ws_26;
  reg                 io_in_r_bypass_regNext_19_0_stall_26;
  reg        [15:0]   io_in_r_bypass_regNext_19_1_data_26;
  reg                 io_in_r_bypass_regNext_19_1_load_store_26;
  reg                 io_in_r_bypass_regNext_19_1_df_is_ws_26;
  reg                 io_in_r_bypass_regNext_19_1_stall_26;
  reg        [15:0]   io_in_r_bypass_regNext_19_2_data_26;
  reg                 io_in_r_bypass_regNext_19_2_load_store_26;
  reg                 io_in_r_bypass_regNext_19_2_df_is_ws_26;
  reg                 io_in_r_bypass_regNext_19_2_stall_26;
  reg        [15:0]   io_in_r_bypass_regNext_19_3_data_26;
  reg                 io_in_r_bypass_regNext_19_3_load_store_26;
  reg                 io_in_r_bypass_regNext_19_3_df_is_ws_26;
  reg                 io_in_r_bypass_regNext_19_3_stall_26;
  reg        [15:0]   io_in_r_bypass_regNext_20_0_data_26;
  reg                 io_in_r_bypass_regNext_20_0_load_store_26;
  reg                 io_in_r_bypass_regNext_20_0_df_is_ws_26;
  reg                 io_in_r_bypass_regNext_20_0_stall_26;
  reg        [15:0]   io_in_r_bypass_regNext_20_1_data_26;
  reg                 io_in_r_bypass_regNext_20_1_load_store_26;
  reg                 io_in_r_bypass_regNext_20_1_df_is_ws_26;
  reg                 io_in_r_bypass_regNext_20_1_stall_26;
  reg        [15:0]   io_in_r_bypass_regNext_20_2_data_26;
  reg                 io_in_r_bypass_regNext_20_2_load_store_26;
  reg                 io_in_r_bypass_regNext_20_2_df_is_ws_26;
  reg                 io_in_r_bypass_regNext_20_2_stall_26;
  reg        [15:0]   io_in_r_bypass_regNext_20_3_data_26;
  reg                 io_in_r_bypass_regNext_20_3_load_store_26;
  reg                 io_in_r_bypass_regNext_20_3_df_is_ws_26;
  reg                 io_in_r_bypass_regNext_20_3_stall_26;
  reg        [15:0]   io_in_r_bypass_regNext_21_0_data_26;
  reg                 io_in_r_bypass_regNext_21_0_load_store_26;
  reg                 io_in_r_bypass_regNext_21_0_df_is_ws_26;
  reg                 io_in_r_bypass_regNext_21_0_stall_26;
  reg        [15:0]   io_in_r_bypass_regNext_21_1_data_26;
  reg                 io_in_r_bypass_regNext_21_1_load_store_26;
  reg                 io_in_r_bypass_regNext_21_1_df_is_ws_26;
  reg                 io_in_r_bypass_regNext_21_1_stall_26;
  reg        [15:0]   io_in_r_bypass_regNext_21_2_data_26;
  reg                 io_in_r_bypass_regNext_21_2_load_store_26;
  reg                 io_in_r_bypass_regNext_21_2_df_is_ws_26;
  reg                 io_in_r_bypass_regNext_21_2_stall_26;
  reg        [15:0]   io_in_r_bypass_regNext_21_3_data_26;
  reg                 io_in_r_bypass_regNext_21_3_load_store_26;
  reg                 io_in_r_bypass_regNext_21_3_df_is_ws_26;
  reg                 io_in_r_bypass_regNext_21_3_stall_26;
  reg        [15:0]   io_in_r_bypass_regNext_22_0_data_26;
  reg                 io_in_r_bypass_regNext_22_0_load_store_26;
  reg                 io_in_r_bypass_regNext_22_0_df_is_ws_26;
  reg                 io_in_r_bypass_regNext_22_0_stall_26;
  reg        [15:0]   io_in_r_bypass_regNext_22_1_data_26;
  reg                 io_in_r_bypass_regNext_22_1_load_store_26;
  reg                 io_in_r_bypass_regNext_22_1_df_is_ws_26;
  reg                 io_in_r_bypass_regNext_22_1_stall_26;
  reg        [15:0]   io_in_r_bypass_regNext_22_2_data_26;
  reg                 io_in_r_bypass_regNext_22_2_load_store_26;
  reg                 io_in_r_bypass_regNext_22_2_df_is_ws_26;
  reg                 io_in_r_bypass_regNext_22_2_stall_26;
  reg        [15:0]   io_in_r_bypass_regNext_22_3_data_26;
  reg                 io_in_r_bypass_regNext_22_3_load_store_26;
  reg                 io_in_r_bypass_regNext_22_3_df_is_ws_26;
  reg                 io_in_r_bypass_regNext_22_3_stall_26;
  reg        [15:0]   io_in_r_bypass_regNext_23_0_data_26;
  reg                 io_in_r_bypass_regNext_23_0_load_store_26;
  reg                 io_in_r_bypass_regNext_23_0_df_is_ws_26;
  reg                 io_in_r_bypass_regNext_23_0_stall_26;
  reg        [15:0]   io_in_r_bypass_regNext_23_1_data_26;
  reg                 io_in_r_bypass_regNext_23_1_load_store_26;
  reg                 io_in_r_bypass_regNext_23_1_df_is_ws_26;
  reg                 io_in_r_bypass_regNext_23_1_stall_26;
  reg        [15:0]   io_in_r_bypass_regNext_23_2_data_26;
  reg                 io_in_r_bypass_regNext_23_2_load_store_26;
  reg                 io_in_r_bypass_regNext_23_2_df_is_ws_26;
  reg                 io_in_r_bypass_regNext_23_2_stall_26;
  reg        [15:0]   io_in_r_bypass_regNext_23_3_data_26;
  reg                 io_in_r_bypass_regNext_23_3_load_store_26;
  reg                 io_in_r_bypass_regNext_23_3_df_is_ws_26;
  reg                 io_in_r_bypass_regNext_23_3_stall_26;
  reg        [15:0]   io_in_r_bypass_regNext_24_0_data_26;
  reg                 io_in_r_bypass_regNext_24_0_load_store_26;
  reg                 io_in_r_bypass_regNext_24_0_df_is_ws_26;
  reg                 io_in_r_bypass_regNext_24_0_stall_26;
  reg        [15:0]   io_in_r_bypass_regNext_24_1_data_26;
  reg                 io_in_r_bypass_regNext_24_1_load_store_26;
  reg                 io_in_r_bypass_regNext_24_1_df_is_ws_26;
  reg                 io_in_r_bypass_regNext_24_1_stall_26;
  reg        [15:0]   io_in_r_bypass_regNext_24_2_data_26;
  reg                 io_in_r_bypass_regNext_24_2_load_store_26;
  reg                 io_in_r_bypass_regNext_24_2_df_is_ws_26;
  reg                 io_in_r_bypass_regNext_24_2_stall_26;
  reg        [15:0]   io_in_r_bypass_regNext_24_3_data_26;
  reg                 io_in_r_bypass_regNext_24_3_load_store_26;
  reg                 io_in_r_bypass_regNext_24_3_df_is_ws_26;
  reg                 io_in_r_bypass_regNext_24_3_stall_26;
  reg        [15:0]   io_in_r_bypass_regNext_25_0_data_26;
  reg                 io_in_r_bypass_regNext_25_0_load_store_26;
  reg                 io_in_r_bypass_regNext_25_0_df_is_ws_26;
  reg                 io_in_r_bypass_regNext_25_0_stall_26;
  reg        [15:0]   io_in_r_bypass_regNext_25_1_data_26;
  reg                 io_in_r_bypass_regNext_25_1_load_store_26;
  reg                 io_in_r_bypass_regNext_25_1_df_is_ws_26;
  reg                 io_in_r_bypass_regNext_25_1_stall_26;
  reg        [15:0]   io_in_r_bypass_regNext_25_2_data_26;
  reg                 io_in_r_bypass_regNext_25_2_load_store_26;
  reg                 io_in_r_bypass_regNext_25_2_df_is_ws_26;
  reg                 io_in_r_bypass_regNext_25_2_stall_26;
  reg        [15:0]   io_in_r_bypass_regNext_25_3_data_26;
  reg                 io_in_r_bypass_regNext_25_3_load_store_26;
  reg                 io_in_r_bypass_regNext_25_3_df_is_ws_26;
  reg                 io_in_r_bypass_regNext_25_3_stall_26;
  reg        [15:0]   io_in_r_bypass_regNext_26_0_data_26;
  reg                 io_in_r_bypass_regNext_26_0_load_store_26;
  reg                 io_in_r_bypass_regNext_26_0_df_is_ws_26;
  reg                 io_in_r_bypass_regNext_26_0_stall_26;
  reg        [15:0]   io_in_r_bypass_regNext_26_1_data_26;
  reg                 io_in_r_bypass_regNext_26_1_load_store_26;
  reg                 io_in_r_bypass_regNext_26_1_df_is_ws_26;
  reg                 io_in_r_bypass_regNext_26_1_stall_26;
  reg        [15:0]   io_in_r_bypass_regNext_26_2_data_26;
  reg                 io_in_r_bypass_regNext_26_2_load_store_26;
  reg                 io_in_r_bypass_regNext_26_2_df_is_ws_26;
  reg                 io_in_r_bypass_regNext_26_2_stall_26;
  reg        [15:0]   io_in_r_bypass_regNext_26_3_data_26;
  reg                 io_in_r_bypass_regNext_26_3_load_store_26;
  reg                 io_in_r_bypass_regNext_26_3_df_is_ws_26;
  reg                 io_in_r_bypass_regNext_26_3_stall_26;
  reg        [15:0]   io_in_r_bypass_regNext_27_0_data_26;
  reg                 io_in_r_bypass_regNext_27_0_load_store_26;
  reg                 io_in_r_bypass_regNext_27_0_df_is_ws_26;
  reg                 io_in_r_bypass_regNext_27_0_stall_26;
  reg        [15:0]   io_in_r_bypass_regNext_27_1_data_26;
  reg                 io_in_r_bypass_regNext_27_1_load_store_26;
  reg                 io_in_r_bypass_regNext_27_1_df_is_ws_26;
  reg                 io_in_r_bypass_regNext_27_1_stall_26;
  reg        [15:0]   io_in_r_bypass_regNext_27_2_data_26;
  reg                 io_in_r_bypass_regNext_27_2_load_store_26;
  reg                 io_in_r_bypass_regNext_27_2_df_is_ws_26;
  reg                 io_in_r_bypass_regNext_27_2_stall_26;
  reg        [15:0]   io_in_r_bypass_regNext_27_3_data_26;
  reg                 io_in_r_bypass_regNext_27_3_load_store_26;
  reg                 io_in_r_bypass_regNext_27_3_df_is_ws_26;
  reg                 io_in_r_bypass_regNext_27_3_stall_26;
  reg        [15:0]   io_in_r_bypass_regNext_28_0_data_26;
  reg                 io_in_r_bypass_regNext_28_0_load_store_26;
  reg                 io_in_r_bypass_regNext_28_0_df_is_ws_26;
  reg                 io_in_r_bypass_regNext_28_0_stall_26;
  reg        [15:0]   io_in_r_bypass_regNext_28_1_data_26;
  reg                 io_in_r_bypass_regNext_28_1_load_store_26;
  reg                 io_in_r_bypass_regNext_28_1_df_is_ws_26;
  reg                 io_in_r_bypass_regNext_28_1_stall_26;
  reg        [15:0]   io_in_r_bypass_regNext_28_2_data_26;
  reg                 io_in_r_bypass_regNext_28_2_load_store_26;
  reg                 io_in_r_bypass_regNext_28_2_df_is_ws_26;
  reg                 io_in_r_bypass_regNext_28_2_stall_26;
  reg        [15:0]   io_in_r_bypass_regNext_28_3_data_26;
  reg                 io_in_r_bypass_regNext_28_3_load_store_26;
  reg                 io_in_r_bypass_regNext_28_3_df_is_ws_26;
  reg                 io_in_r_bypass_regNext_28_3_stall_26;
  reg        [15:0]   io_in_r_bypass_regNext_29_0_data_26;
  reg                 io_in_r_bypass_regNext_29_0_load_store_26;
  reg                 io_in_r_bypass_regNext_29_0_df_is_ws_26;
  reg                 io_in_r_bypass_regNext_29_0_stall_26;
  reg        [15:0]   io_in_r_bypass_regNext_29_1_data_26;
  reg                 io_in_r_bypass_regNext_29_1_load_store_26;
  reg                 io_in_r_bypass_regNext_29_1_df_is_ws_26;
  reg                 io_in_r_bypass_regNext_29_1_stall_26;
  reg        [15:0]   io_in_r_bypass_regNext_29_2_data_26;
  reg                 io_in_r_bypass_regNext_29_2_load_store_26;
  reg                 io_in_r_bypass_regNext_29_2_df_is_ws_26;
  reg                 io_in_r_bypass_regNext_29_2_stall_26;
  reg        [15:0]   io_in_r_bypass_regNext_29_3_data_26;
  reg                 io_in_r_bypass_regNext_29_3_load_store_26;
  reg                 io_in_r_bypass_regNext_29_3_df_is_ws_26;
  reg                 io_in_r_bypass_regNext_29_3_stall_26;
  reg        [15:0]   io_in_r_bypass_regNext_30_0_data_26;
  reg                 io_in_r_bypass_regNext_30_0_load_store_26;
  reg                 io_in_r_bypass_regNext_30_0_df_is_ws_26;
  reg                 io_in_r_bypass_regNext_30_0_stall_26;
  reg        [15:0]   io_in_r_bypass_regNext_30_1_data_26;
  reg                 io_in_r_bypass_regNext_30_1_load_store_26;
  reg                 io_in_r_bypass_regNext_30_1_df_is_ws_26;
  reg                 io_in_r_bypass_regNext_30_1_stall_26;
  reg        [15:0]   io_in_r_bypass_regNext_30_2_data_26;
  reg                 io_in_r_bypass_regNext_30_2_load_store_26;
  reg                 io_in_r_bypass_regNext_30_2_df_is_ws_26;
  reg                 io_in_r_bypass_regNext_30_2_stall_26;
  reg        [15:0]   io_in_r_bypass_regNext_30_3_data_26;
  reg                 io_in_r_bypass_regNext_30_3_load_store_26;
  reg                 io_in_r_bypass_regNext_30_3_df_is_ws_26;
  reg                 io_in_r_bypass_regNext_30_3_stall_26;
  reg        [15:0]   io_in_r_bypass_regNext_31_0_data_26;
  reg                 io_in_r_bypass_regNext_31_0_load_store_26;
  reg                 io_in_r_bypass_regNext_31_0_df_is_ws_26;
  reg                 io_in_r_bypass_regNext_31_0_stall_26;
  reg        [15:0]   io_in_r_bypass_regNext_31_1_data_26;
  reg                 io_in_r_bypass_regNext_31_1_load_store_26;
  reg                 io_in_r_bypass_regNext_31_1_df_is_ws_26;
  reg                 io_in_r_bypass_regNext_31_1_stall_26;
  reg        [15:0]   io_in_r_bypass_regNext_31_2_data_26;
  reg                 io_in_r_bypass_regNext_31_2_load_store_26;
  reg                 io_in_r_bypass_regNext_31_2_df_is_ws_26;
  reg                 io_in_r_bypass_regNext_31_2_stall_26;
  reg        [15:0]   io_in_r_bypass_regNext_31_3_data_26;
  reg                 io_in_r_bypass_regNext_31_3_load_store_26;
  reg                 io_in_r_bypass_regNext_31_3_df_is_ws_26;
  reg                 io_in_r_bypass_regNext_31_3_stall_26;
  reg        [15:0]   io_in_r_bypass_regNext_0_0_data_27;
  reg                 io_in_r_bypass_regNext_0_0_load_store_27;
  reg                 io_in_r_bypass_regNext_0_0_df_is_ws_27;
  reg                 io_in_r_bypass_regNext_0_0_stall_27;
  reg        [15:0]   io_in_r_bypass_regNext_0_1_data_27;
  reg                 io_in_r_bypass_regNext_0_1_load_store_27;
  reg                 io_in_r_bypass_regNext_0_1_df_is_ws_27;
  reg                 io_in_r_bypass_regNext_0_1_stall_27;
  reg        [15:0]   io_in_r_bypass_regNext_0_2_data_27;
  reg                 io_in_r_bypass_regNext_0_2_load_store_27;
  reg                 io_in_r_bypass_regNext_0_2_df_is_ws_27;
  reg                 io_in_r_bypass_regNext_0_2_stall_27;
  reg        [15:0]   io_in_r_bypass_regNext_0_3_data_27;
  reg                 io_in_r_bypass_regNext_0_3_load_store_27;
  reg                 io_in_r_bypass_regNext_0_3_df_is_ws_27;
  reg                 io_in_r_bypass_regNext_0_3_stall_27;
  reg        [15:0]   io_in_r_bypass_regNext_1_0_data_27;
  reg                 io_in_r_bypass_regNext_1_0_load_store_27;
  reg                 io_in_r_bypass_regNext_1_0_df_is_ws_27;
  reg                 io_in_r_bypass_regNext_1_0_stall_27;
  reg        [15:0]   io_in_r_bypass_regNext_1_1_data_27;
  reg                 io_in_r_bypass_regNext_1_1_load_store_27;
  reg                 io_in_r_bypass_regNext_1_1_df_is_ws_27;
  reg                 io_in_r_bypass_regNext_1_1_stall_27;
  reg        [15:0]   io_in_r_bypass_regNext_1_2_data_27;
  reg                 io_in_r_bypass_regNext_1_2_load_store_27;
  reg                 io_in_r_bypass_regNext_1_2_df_is_ws_27;
  reg                 io_in_r_bypass_regNext_1_2_stall_27;
  reg        [15:0]   io_in_r_bypass_regNext_1_3_data_27;
  reg                 io_in_r_bypass_regNext_1_3_load_store_27;
  reg                 io_in_r_bypass_regNext_1_3_df_is_ws_27;
  reg                 io_in_r_bypass_regNext_1_3_stall_27;
  reg        [15:0]   io_in_r_bypass_regNext_2_0_data_27;
  reg                 io_in_r_bypass_regNext_2_0_load_store_27;
  reg                 io_in_r_bypass_regNext_2_0_df_is_ws_27;
  reg                 io_in_r_bypass_regNext_2_0_stall_27;
  reg        [15:0]   io_in_r_bypass_regNext_2_1_data_27;
  reg                 io_in_r_bypass_regNext_2_1_load_store_27;
  reg                 io_in_r_bypass_regNext_2_1_df_is_ws_27;
  reg                 io_in_r_bypass_regNext_2_1_stall_27;
  reg        [15:0]   io_in_r_bypass_regNext_2_2_data_27;
  reg                 io_in_r_bypass_regNext_2_2_load_store_27;
  reg                 io_in_r_bypass_regNext_2_2_df_is_ws_27;
  reg                 io_in_r_bypass_regNext_2_2_stall_27;
  reg        [15:0]   io_in_r_bypass_regNext_2_3_data_27;
  reg                 io_in_r_bypass_regNext_2_3_load_store_27;
  reg                 io_in_r_bypass_regNext_2_3_df_is_ws_27;
  reg                 io_in_r_bypass_regNext_2_3_stall_27;
  reg        [15:0]   io_in_r_bypass_regNext_3_0_data_27;
  reg                 io_in_r_bypass_regNext_3_0_load_store_27;
  reg                 io_in_r_bypass_regNext_3_0_df_is_ws_27;
  reg                 io_in_r_bypass_regNext_3_0_stall_27;
  reg        [15:0]   io_in_r_bypass_regNext_3_1_data_27;
  reg                 io_in_r_bypass_regNext_3_1_load_store_27;
  reg                 io_in_r_bypass_regNext_3_1_df_is_ws_27;
  reg                 io_in_r_bypass_regNext_3_1_stall_27;
  reg        [15:0]   io_in_r_bypass_regNext_3_2_data_27;
  reg                 io_in_r_bypass_regNext_3_2_load_store_27;
  reg                 io_in_r_bypass_regNext_3_2_df_is_ws_27;
  reg                 io_in_r_bypass_regNext_3_2_stall_27;
  reg        [15:0]   io_in_r_bypass_regNext_3_3_data_27;
  reg                 io_in_r_bypass_regNext_3_3_load_store_27;
  reg                 io_in_r_bypass_regNext_3_3_df_is_ws_27;
  reg                 io_in_r_bypass_regNext_3_3_stall_27;
  reg        [15:0]   io_in_r_bypass_regNext_4_0_data_27;
  reg                 io_in_r_bypass_regNext_4_0_load_store_27;
  reg                 io_in_r_bypass_regNext_4_0_df_is_ws_27;
  reg                 io_in_r_bypass_regNext_4_0_stall_27;
  reg        [15:0]   io_in_r_bypass_regNext_4_1_data_27;
  reg                 io_in_r_bypass_regNext_4_1_load_store_27;
  reg                 io_in_r_bypass_regNext_4_1_df_is_ws_27;
  reg                 io_in_r_bypass_regNext_4_1_stall_27;
  reg        [15:0]   io_in_r_bypass_regNext_4_2_data_27;
  reg                 io_in_r_bypass_regNext_4_2_load_store_27;
  reg                 io_in_r_bypass_regNext_4_2_df_is_ws_27;
  reg                 io_in_r_bypass_regNext_4_2_stall_27;
  reg        [15:0]   io_in_r_bypass_regNext_4_3_data_27;
  reg                 io_in_r_bypass_regNext_4_3_load_store_27;
  reg                 io_in_r_bypass_regNext_4_3_df_is_ws_27;
  reg                 io_in_r_bypass_regNext_4_3_stall_27;
  reg        [15:0]   io_in_r_bypass_regNext_5_0_data_27;
  reg                 io_in_r_bypass_regNext_5_0_load_store_27;
  reg                 io_in_r_bypass_regNext_5_0_df_is_ws_27;
  reg                 io_in_r_bypass_regNext_5_0_stall_27;
  reg        [15:0]   io_in_r_bypass_regNext_5_1_data_27;
  reg                 io_in_r_bypass_regNext_5_1_load_store_27;
  reg                 io_in_r_bypass_regNext_5_1_df_is_ws_27;
  reg                 io_in_r_bypass_regNext_5_1_stall_27;
  reg        [15:0]   io_in_r_bypass_regNext_5_2_data_27;
  reg                 io_in_r_bypass_regNext_5_2_load_store_27;
  reg                 io_in_r_bypass_regNext_5_2_df_is_ws_27;
  reg                 io_in_r_bypass_regNext_5_2_stall_27;
  reg        [15:0]   io_in_r_bypass_regNext_5_3_data_27;
  reg                 io_in_r_bypass_regNext_5_3_load_store_27;
  reg                 io_in_r_bypass_regNext_5_3_df_is_ws_27;
  reg                 io_in_r_bypass_regNext_5_3_stall_27;
  reg        [15:0]   io_in_r_bypass_regNext_6_0_data_27;
  reg                 io_in_r_bypass_regNext_6_0_load_store_27;
  reg                 io_in_r_bypass_regNext_6_0_df_is_ws_27;
  reg                 io_in_r_bypass_regNext_6_0_stall_27;
  reg        [15:0]   io_in_r_bypass_regNext_6_1_data_27;
  reg                 io_in_r_bypass_regNext_6_1_load_store_27;
  reg                 io_in_r_bypass_regNext_6_1_df_is_ws_27;
  reg                 io_in_r_bypass_regNext_6_1_stall_27;
  reg        [15:0]   io_in_r_bypass_regNext_6_2_data_27;
  reg                 io_in_r_bypass_regNext_6_2_load_store_27;
  reg                 io_in_r_bypass_regNext_6_2_df_is_ws_27;
  reg                 io_in_r_bypass_regNext_6_2_stall_27;
  reg        [15:0]   io_in_r_bypass_regNext_6_3_data_27;
  reg                 io_in_r_bypass_regNext_6_3_load_store_27;
  reg                 io_in_r_bypass_regNext_6_3_df_is_ws_27;
  reg                 io_in_r_bypass_regNext_6_3_stall_27;
  reg        [15:0]   io_in_r_bypass_regNext_7_0_data_27;
  reg                 io_in_r_bypass_regNext_7_0_load_store_27;
  reg                 io_in_r_bypass_regNext_7_0_df_is_ws_27;
  reg                 io_in_r_bypass_regNext_7_0_stall_27;
  reg        [15:0]   io_in_r_bypass_regNext_7_1_data_27;
  reg                 io_in_r_bypass_regNext_7_1_load_store_27;
  reg                 io_in_r_bypass_regNext_7_1_df_is_ws_27;
  reg                 io_in_r_bypass_regNext_7_1_stall_27;
  reg        [15:0]   io_in_r_bypass_regNext_7_2_data_27;
  reg                 io_in_r_bypass_regNext_7_2_load_store_27;
  reg                 io_in_r_bypass_regNext_7_2_df_is_ws_27;
  reg                 io_in_r_bypass_regNext_7_2_stall_27;
  reg        [15:0]   io_in_r_bypass_regNext_7_3_data_27;
  reg                 io_in_r_bypass_regNext_7_3_load_store_27;
  reg                 io_in_r_bypass_regNext_7_3_df_is_ws_27;
  reg                 io_in_r_bypass_regNext_7_3_stall_27;
  reg        [15:0]   io_in_r_bypass_regNext_8_0_data_27;
  reg                 io_in_r_bypass_regNext_8_0_load_store_27;
  reg                 io_in_r_bypass_regNext_8_0_df_is_ws_27;
  reg                 io_in_r_bypass_regNext_8_0_stall_27;
  reg        [15:0]   io_in_r_bypass_regNext_8_1_data_27;
  reg                 io_in_r_bypass_regNext_8_1_load_store_27;
  reg                 io_in_r_bypass_regNext_8_1_df_is_ws_27;
  reg                 io_in_r_bypass_regNext_8_1_stall_27;
  reg        [15:0]   io_in_r_bypass_regNext_8_2_data_27;
  reg                 io_in_r_bypass_regNext_8_2_load_store_27;
  reg                 io_in_r_bypass_regNext_8_2_df_is_ws_27;
  reg                 io_in_r_bypass_regNext_8_2_stall_27;
  reg        [15:0]   io_in_r_bypass_regNext_8_3_data_27;
  reg                 io_in_r_bypass_regNext_8_3_load_store_27;
  reg                 io_in_r_bypass_regNext_8_3_df_is_ws_27;
  reg                 io_in_r_bypass_regNext_8_3_stall_27;
  reg        [15:0]   io_in_r_bypass_regNext_9_0_data_27;
  reg                 io_in_r_bypass_regNext_9_0_load_store_27;
  reg                 io_in_r_bypass_regNext_9_0_df_is_ws_27;
  reg                 io_in_r_bypass_regNext_9_0_stall_27;
  reg        [15:0]   io_in_r_bypass_regNext_9_1_data_27;
  reg                 io_in_r_bypass_regNext_9_1_load_store_27;
  reg                 io_in_r_bypass_regNext_9_1_df_is_ws_27;
  reg                 io_in_r_bypass_regNext_9_1_stall_27;
  reg        [15:0]   io_in_r_bypass_regNext_9_2_data_27;
  reg                 io_in_r_bypass_regNext_9_2_load_store_27;
  reg                 io_in_r_bypass_regNext_9_2_df_is_ws_27;
  reg                 io_in_r_bypass_regNext_9_2_stall_27;
  reg        [15:0]   io_in_r_bypass_regNext_9_3_data_27;
  reg                 io_in_r_bypass_regNext_9_3_load_store_27;
  reg                 io_in_r_bypass_regNext_9_3_df_is_ws_27;
  reg                 io_in_r_bypass_regNext_9_3_stall_27;
  reg        [15:0]   io_in_r_bypass_regNext_10_0_data_27;
  reg                 io_in_r_bypass_regNext_10_0_load_store_27;
  reg                 io_in_r_bypass_regNext_10_0_df_is_ws_27;
  reg                 io_in_r_bypass_regNext_10_0_stall_27;
  reg        [15:0]   io_in_r_bypass_regNext_10_1_data_27;
  reg                 io_in_r_bypass_regNext_10_1_load_store_27;
  reg                 io_in_r_bypass_regNext_10_1_df_is_ws_27;
  reg                 io_in_r_bypass_regNext_10_1_stall_27;
  reg        [15:0]   io_in_r_bypass_regNext_10_2_data_27;
  reg                 io_in_r_bypass_regNext_10_2_load_store_27;
  reg                 io_in_r_bypass_regNext_10_2_df_is_ws_27;
  reg                 io_in_r_bypass_regNext_10_2_stall_27;
  reg        [15:0]   io_in_r_bypass_regNext_10_3_data_27;
  reg                 io_in_r_bypass_regNext_10_3_load_store_27;
  reg                 io_in_r_bypass_regNext_10_3_df_is_ws_27;
  reg                 io_in_r_bypass_regNext_10_3_stall_27;
  reg        [15:0]   io_in_r_bypass_regNext_11_0_data_27;
  reg                 io_in_r_bypass_regNext_11_0_load_store_27;
  reg                 io_in_r_bypass_regNext_11_0_df_is_ws_27;
  reg                 io_in_r_bypass_regNext_11_0_stall_27;
  reg        [15:0]   io_in_r_bypass_regNext_11_1_data_27;
  reg                 io_in_r_bypass_regNext_11_1_load_store_27;
  reg                 io_in_r_bypass_regNext_11_1_df_is_ws_27;
  reg                 io_in_r_bypass_regNext_11_1_stall_27;
  reg        [15:0]   io_in_r_bypass_regNext_11_2_data_27;
  reg                 io_in_r_bypass_regNext_11_2_load_store_27;
  reg                 io_in_r_bypass_regNext_11_2_df_is_ws_27;
  reg                 io_in_r_bypass_regNext_11_2_stall_27;
  reg        [15:0]   io_in_r_bypass_regNext_11_3_data_27;
  reg                 io_in_r_bypass_regNext_11_3_load_store_27;
  reg                 io_in_r_bypass_regNext_11_3_df_is_ws_27;
  reg                 io_in_r_bypass_regNext_11_3_stall_27;
  reg        [15:0]   io_in_r_bypass_regNext_12_0_data_27;
  reg                 io_in_r_bypass_regNext_12_0_load_store_27;
  reg                 io_in_r_bypass_regNext_12_0_df_is_ws_27;
  reg                 io_in_r_bypass_regNext_12_0_stall_27;
  reg        [15:0]   io_in_r_bypass_regNext_12_1_data_27;
  reg                 io_in_r_bypass_regNext_12_1_load_store_27;
  reg                 io_in_r_bypass_regNext_12_1_df_is_ws_27;
  reg                 io_in_r_bypass_regNext_12_1_stall_27;
  reg        [15:0]   io_in_r_bypass_regNext_12_2_data_27;
  reg                 io_in_r_bypass_regNext_12_2_load_store_27;
  reg                 io_in_r_bypass_regNext_12_2_df_is_ws_27;
  reg                 io_in_r_bypass_regNext_12_2_stall_27;
  reg        [15:0]   io_in_r_bypass_regNext_12_3_data_27;
  reg                 io_in_r_bypass_regNext_12_3_load_store_27;
  reg                 io_in_r_bypass_regNext_12_3_df_is_ws_27;
  reg                 io_in_r_bypass_regNext_12_3_stall_27;
  reg        [15:0]   io_in_r_bypass_regNext_13_0_data_27;
  reg                 io_in_r_bypass_regNext_13_0_load_store_27;
  reg                 io_in_r_bypass_regNext_13_0_df_is_ws_27;
  reg                 io_in_r_bypass_regNext_13_0_stall_27;
  reg        [15:0]   io_in_r_bypass_regNext_13_1_data_27;
  reg                 io_in_r_bypass_regNext_13_1_load_store_27;
  reg                 io_in_r_bypass_regNext_13_1_df_is_ws_27;
  reg                 io_in_r_bypass_regNext_13_1_stall_27;
  reg        [15:0]   io_in_r_bypass_regNext_13_2_data_27;
  reg                 io_in_r_bypass_regNext_13_2_load_store_27;
  reg                 io_in_r_bypass_regNext_13_2_df_is_ws_27;
  reg                 io_in_r_bypass_regNext_13_2_stall_27;
  reg        [15:0]   io_in_r_bypass_regNext_13_3_data_27;
  reg                 io_in_r_bypass_regNext_13_3_load_store_27;
  reg                 io_in_r_bypass_regNext_13_3_df_is_ws_27;
  reg                 io_in_r_bypass_regNext_13_3_stall_27;
  reg        [15:0]   io_in_r_bypass_regNext_14_0_data_27;
  reg                 io_in_r_bypass_regNext_14_0_load_store_27;
  reg                 io_in_r_bypass_regNext_14_0_df_is_ws_27;
  reg                 io_in_r_bypass_regNext_14_0_stall_27;
  reg        [15:0]   io_in_r_bypass_regNext_14_1_data_27;
  reg                 io_in_r_bypass_regNext_14_1_load_store_27;
  reg                 io_in_r_bypass_regNext_14_1_df_is_ws_27;
  reg                 io_in_r_bypass_regNext_14_1_stall_27;
  reg        [15:0]   io_in_r_bypass_regNext_14_2_data_27;
  reg                 io_in_r_bypass_regNext_14_2_load_store_27;
  reg                 io_in_r_bypass_regNext_14_2_df_is_ws_27;
  reg                 io_in_r_bypass_regNext_14_2_stall_27;
  reg        [15:0]   io_in_r_bypass_regNext_14_3_data_27;
  reg                 io_in_r_bypass_regNext_14_3_load_store_27;
  reg                 io_in_r_bypass_regNext_14_3_df_is_ws_27;
  reg                 io_in_r_bypass_regNext_14_3_stall_27;
  reg        [15:0]   io_in_r_bypass_regNext_15_0_data_27;
  reg                 io_in_r_bypass_regNext_15_0_load_store_27;
  reg                 io_in_r_bypass_regNext_15_0_df_is_ws_27;
  reg                 io_in_r_bypass_regNext_15_0_stall_27;
  reg        [15:0]   io_in_r_bypass_regNext_15_1_data_27;
  reg                 io_in_r_bypass_regNext_15_1_load_store_27;
  reg                 io_in_r_bypass_regNext_15_1_df_is_ws_27;
  reg                 io_in_r_bypass_regNext_15_1_stall_27;
  reg        [15:0]   io_in_r_bypass_regNext_15_2_data_27;
  reg                 io_in_r_bypass_regNext_15_2_load_store_27;
  reg                 io_in_r_bypass_regNext_15_2_df_is_ws_27;
  reg                 io_in_r_bypass_regNext_15_2_stall_27;
  reg        [15:0]   io_in_r_bypass_regNext_15_3_data_27;
  reg                 io_in_r_bypass_regNext_15_3_load_store_27;
  reg                 io_in_r_bypass_regNext_15_3_df_is_ws_27;
  reg                 io_in_r_bypass_regNext_15_3_stall_27;
  reg        [15:0]   io_in_r_bypass_regNext_16_0_data_27;
  reg                 io_in_r_bypass_regNext_16_0_load_store_27;
  reg                 io_in_r_bypass_regNext_16_0_df_is_ws_27;
  reg                 io_in_r_bypass_regNext_16_0_stall_27;
  reg        [15:0]   io_in_r_bypass_regNext_16_1_data_27;
  reg                 io_in_r_bypass_regNext_16_1_load_store_27;
  reg                 io_in_r_bypass_regNext_16_1_df_is_ws_27;
  reg                 io_in_r_bypass_regNext_16_1_stall_27;
  reg        [15:0]   io_in_r_bypass_regNext_16_2_data_27;
  reg                 io_in_r_bypass_regNext_16_2_load_store_27;
  reg                 io_in_r_bypass_regNext_16_2_df_is_ws_27;
  reg                 io_in_r_bypass_regNext_16_2_stall_27;
  reg        [15:0]   io_in_r_bypass_regNext_16_3_data_27;
  reg                 io_in_r_bypass_regNext_16_3_load_store_27;
  reg                 io_in_r_bypass_regNext_16_3_df_is_ws_27;
  reg                 io_in_r_bypass_regNext_16_3_stall_27;
  reg        [15:0]   io_in_r_bypass_regNext_17_0_data_27;
  reg                 io_in_r_bypass_regNext_17_0_load_store_27;
  reg                 io_in_r_bypass_regNext_17_0_df_is_ws_27;
  reg                 io_in_r_bypass_regNext_17_0_stall_27;
  reg        [15:0]   io_in_r_bypass_regNext_17_1_data_27;
  reg                 io_in_r_bypass_regNext_17_1_load_store_27;
  reg                 io_in_r_bypass_regNext_17_1_df_is_ws_27;
  reg                 io_in_r_bypass_regNext_17_1_stall_27;
  reg        [15:0]   io_in_r_bypass_regNext_17_2_data_27;
  reg                 io_in_r_bypass_regNext_17_2_load_store_27;
  reg                 io_in_r_bypass_regNext_17_2_df_is_ws_27;
  reg                 io_in_r_bypass_regNext_17_2_stall_27;
  reg        [15:0]   io_in_r_bypass_regNext_17_3_data_27;
  reg                 io_in_r_bypass_regNext_17_3_load_store_27;
  reg                 io_in_r_bypass_regNext_17_3_df_is_ws_27;
  reg                 io_in_r_bypass_regNext_17_3_stall_27;
  reg        [15:0]   io_in_r_bypass_regNext_18_0_data_27;
  reg                 io_in_r_bypass_regNext_18_0_load_store_27;
  reg                 io_in_r_bypass_regNext_18_0_df_is_ws_27;
  reg                 io_in_r_bypass_regNext_18_0_stall_27;
  reg        [15:0]   io_in_r_bypass_regNext_18_1_data_27;
  reg                 io_in_r_bypass_regNext_18_1_load_store_27;
  reg                 io_in_r_bypass_regNext_18_1_df_is_ws_27;
  reg                 io_in_r_bypass_regNext_18_1_stall_27;
  reg        [15:0]   io_in_r_bypass_regNext_18_2_data_27;
  reg                 io_in_r_bypass_regNext_18_2_load_store_27;
  reg                 io_in_r_bypass_regNext_18_2_df_is_ws_27;
  reg                 io_in_r_bypass_regNext_18_2_stall_27;
  reg        [15:0]   io_in_r_bypass_regNext_18_3_data_27;
  reg                 io_in_r_bypass_regNext_18_3_load_store_27;
  reg                 io_in_r_bypass_regNext_18_3_df_is_ws_27;
  reg                 io_in_r_bypass_regNext_18_3_stall_27;
  reg        [15:0]   io_in_r_bypass_regNext_19_0_data_27;
  reg                 io_in_r_bypass_regNext_19_0_load_store_27;
  reg                 io_in_r_bypass_regNext_19_0_df_is_ws_27;
  reg                 io_in_r_bypass_regNext_19_0_stall_27;
  reg        [15:0]   io_in_r_bypass_regNext_19_1_data_27;
  reg                 io_in_r_bypass_regNext_19_1_load_store_27;
  reg                 io_in_r_bypass_regNext_19_1_df_is_ws_27;
  reg                 io_in_r_bypass_regNext_19_1_stall_27;
  reg        [15:0]   io_in_r_bypass_regNext_19_2_data_27;
  reg                 io_in_r_bypass_regNext_19_2_load_store_27;
  reg                 io_in_r_bypass_regNext_19_2_df_is_ws_27;
  reg                 io_in_r_bypass_regNext_19_2_stall_27;
  reg        [15:0]   io_in_r_bypass_regNext_19_3_data_27;
  reg                 io_in_r_bypass_regNext_19_3_load_store_27;
  reg                 io_in_r_bypass_regNext_19_3_df_is_ws_27;
  reg                 io_in_r_bypass_regNext_19_3_stall_27;
  reg        [15:0]   io_in_r_bypass_regNext_20_0_data_27;
  reg                 io_in_r_bypass_regNext_20_0_load_store_27;
  reg                 io_in_r_bypass_regNext_20_0_df_is_ws_27;
  reg                 io_in_r_bypass_regNext_20_0_stall_27;
  reg        [15:0]   io_in_r_bypass_regNext_20_1_data_27;
  reg                 io_in_r_bypass_regNext_20_1_load_store_27;
  reg                 io_in_r_bypass_regNext_20_1_df_is_ws_27;
  reg                 io_in_r_bypass_regNext_20_1_stall_27;
  reg        [15:0]   io_in_r_bypass_regNext_20_2_data_27;
  reg                 io_in_r_bypass_regNext_20_2_load_store_27;
  reg                 io_in_r_bypass_regNext_20_2_df_is_ws_27;
  reg                 io_in_r_bypass_regNext_20_2_stall_27;
  reg        [15:0]   io_in_r_bypass_regNext_20_3_data_27;
  reg                 io_in_r_bypass_regNext_20_3_load_store_27;
  reg                 io_in_r_bypass_regNext_20_3_df_is_ws_27;
  reg                 io_in_r_bypass_regNext_20_3_stall_27;
  reg        [15:0]   io_in_r_bypass_regNext_21_0_data_27;
  reg                 io_in_r_bypass_regNext_21_0_load_store_27;
  reg                 io_in_r_bypass_regNext_21_0_df_is_ws_27;
  reg                 io_in_r_bypass_regNext_21_0_stall_27;
  reg        [15:0]   io_in_r_bypass_regNext_21_1_data_27;
  reg                 io_in_r_bypass_regNext_21_1_load_store_27;
  reg                 io_in_r_bypass_regNext_21_1_df_is_ws_27;
  reg                 io_in_r_bypass_regNext_21_1_stall_27;
  reg        [15:0]   io_in_r_bypass_regNext_21_2_data_27;
  reg                 io_in_r_bypass_regNext_21_2_load_store_27;
  reg                 io_in_r_bypass_regNext_21_2_df_is_ws_27;
  reg                 io_in_r_bypass_regNext_21_2_stall_27;
  reg        [15:0]   io_in_r_bypass_regNext_21_3_data_27;
  reg                 io_in_r_bypass_regNext_21_3_load_store_27;
  reg                 io_in_r_bypass_regNext_21_3_df_is_ws_27;
  reg                 io_in_r_bypass_regNext_21_3_stall_27;
  reg        [15:0]   io_in_r_bypass_regNext_22_0_data_27;
  reg                 io_in_r_bypass_regNext_22_0_load_store_27;
  reg                 io_in_r_bypass_regNext_22_0_df_is_ws_27;
  reg                 io_in_r_bypass_regNext_22_0_stall_27;
  reg        [15:0]   io_in_r_bypass_regNext_22_1_data_27;
  reg                 io_in_r_bypass_regNext_22_1_load_store_27;
  reg                 io_in_r_bypass_regNext_22_1_df_is_ws_27;
  reg                 io_in_r_bypass_regNext_22_1_stall_27;
  reg        [15:0]   io_in_r_bypass_regNext_22_2_data_27;
  reg                 io_in_r_bypass_regNext_22_2_load_store_27;
  reg                 io_in_r_bypass_regNext_22_2_df_is_ws_27;
  reg                 io_in_r_bypass_regNext_22_2_stall_27;
  reg        [15:0]   io_in_r_bypass_regNext_22_3_data_27;
  reg                 io_in_r_bypass_regNext_22_3_load_store_27;
  reg                 io_in_r_bypass_regNext_22_3_df_is_ws_27;
  reg                 io_in_r_bypass_regNext_22_3_stall_27;
  reg        [15:0]   io_in_r_bypass_regNext_23_0_data_27;
  reg                 io_in_r_bypass_regNext_23_0_load_store_27;
  reg                 io_in_r_bypass_regNext_23_0_df_is_ws_27;
  reg                 io_in_r_bypass_regNext_23_0_stall_27;
  reg        [15:0]   io_in_r_bypass_regNext_23_1_data_27;
  reg                 io_in_r_bypass_regNext_23_1_load_store_27;
  reg                 io_in_r_bypass_regNext_23_1_df_is_ws_27;
  reg                 io_in_r_bypass_regNext_23_1_stall_27;
  reg        [15:0]   io_in_r_bypass_regNext_23_2_data_27;
  reg                 io_in_r_bypass_regNext_23_2_load_store_27;
  reg                 io_in_r_bypass_regNext_23_2_df_is_ws_27;
  reg                 io_in_r_bypass_regNext_23_2_stall_27;
  reg        [15:0]   io_in_r_bypass_regNext_23_3_data_27;
  reg                 io_in_r_bypass_regNext_23_3_load_store_27;
  reg                 io_in_r_bypass_regNext_23_3_df_is_ws_27;
  reg                 io_in_r_bypass_regNext_23_3_stall_27;
  reg        [15:0]   io_in_r_bypass_regNext_24_0_data_27;
  reg                 io_in_r_bypass_regNext_24_0_load_store_27;
  reg                 io_in_r_bypass_regNext_24_0_df_is_ws_27;
  reg                 io_in_r_bypass_regNext_24_0_stall_27;
  reg        [15:0]   io_in_r_bypass_regNext_24_1_data_27;
  reg                 io_in_r_bypass_regNext_24_1_load_store_27;
  reg                 io_in_r_bypass_regNext_24_1_df_is_ws_27;
  reg                 io_in_r_bypass_regNext_24_1_stall_27;
  reg        [15:0]   io_in_r_bypass_regNext_24_2_data_27;
  reg                 io_in_r_bypass_regNext_24_2_load_store_27;
  reg                 io_in_r_bypass_regNext_24_2_df_is_ws_27;
  reg                 io_in_r_bypass_regNext_24_2_stall_27;
  reg        [15:0]   io_in_r_bypass_regNext_24_3_data_27;
  reg                 io_in_r_bypass_regNext_24_3_load_store_27;
  reg                 io_in_r_bypass_regNext_24_3_df_is_ws_27;
  reg                 io_in_r_bypass_regNext_24_3_stall_27;
  reg        [15:0]   io_in_r_bypass_regNext_25_0_data_27;
  reg                 io_in_r_bypass_regNext_25_0_load_store_27;
  reg                 io_in_r_bypass_regNext_25_0_df_is_ws_27;
  reg                 io_in_r_bypass_regNext_25_0_stall_27;
  reg        [15:0]   io_in_r_bypass_regNext_25_1_data_27;
  reg                 io_in_r_bypass_regNext_25_1_load_store_27;
  reg                 io_in_r_bypass_regNext_25_1_df_is_ws_27;
  reg                 io_in_r_bypass_regNext_25_1_stall_27;
  reg        [15:0]   io_in_r_bypass_regNext_25_2_data_27;
  reg                 io_in_r_bypass_regNext_25_2_load_store_27;
  reg                 io_in_r_bypass_regNext_25_2_df_is_ws_27;
  reg                 io_in_r_bypass_regNext_25_2_stall_27;
  reg        [15:0]   io_in_r_bypass_regNext_25_3_data_27;
  reg                 io_in_r_bypass_regNext_25_3_load_store_27;
  reg                 io_in_r_bypass_regNext_25_3_df_is_ws_27;
  reg                 io_in_r_bypass_regNext_25_3_stall_27;
  reg        [15:0]   io_in_r_bypass_regNext_26_0_data_27;
  reg                 io_in_r_bypass_regNext_26_0_load_store_27;
  reg                 io_in_r_bypass_regNext_26_0_df_is_ws_27;
  reg                 io_in_r_bypass_regNext_26_0_stall_27;
  reg        [15:0]   io_in_r_bypass_regNext_26_1_data_27;
  reg                 io_in_r_bypass_regNext_26_1_load_store_27;
  reg                 io_in_r_bypass_regNext_26_1_df_is_ws_27;
  reg                 io_in_r_bypass_regNext_26_1_stall_27;
  reg        [15:0]   io_in_r_bypass_regNext_26_2_data_27;
  reg                 io_in_r_bypass_regNext_26_2_load_store_27;
  reg                 io_in_r_bypass_regNext_26_2_df_is_ws_27;
  reg                 io_in_r_bypass_regNext_26_2_stall_27;
  reg        [15:0]   io_in_r_bypass_regNext_26_3_data_27;
  reg                 io_in_r_bypass_regNext_26_3_load_store_27;
  reg                 io_in_r_bypass_regNext_26_3_df_is_ws_27;
  reg                 io_in_r_bypass_regNext_26_3_stall_27;
  reg        [15:0]   io_in_r_bypass_regNext_27_0_data_27;
  reg                 io_in_r_bypass_regNext_27_0_load_store_27;
  reg                 io_in_r_bypass_regNext_27_0_df_is_ws_27;
  reg                 io_in_r_bypass_regNext_27_0_stall_27;
  reg        [15:0]   io_in_r_bypass_regNext_27_1_data_27;
  reg                 io_in_r_bypass_regNext_27_1_load_store_27;
  reg                 io_in_r_bypass_regNext_27_1_df_is_ws_27;
  reg                 io_in_r_bypass_regNext_27_1_stall_27;
  reg        [15:0]   io_in_r_bypass_regNext_27_2_data_27;
  reg                 io_in_r_bypass_regNext_27_2_load_store_27;
  reg                 io_in_r_bypass_regNext_27_2_df_is_ws_27;
  reg                 io_in_r_bypass_regNext_27_2_stall_27;
  reg        [15:0]   io_in_r_bypass_regNext_27_3_data_27;
  reg                 io_in_r_bypass_regNext_27_3_load_store_27;
  reg                 io_in_r_bypass_regNext_27_3_df_is_ws_27;
  reg                 io_in_r_bypass_regNext_27_3_stall_27;
  reg        [15:0]   io_in_r_bypass_regNext_28_0_data_27;
  reg                 io_in_r_bypass_regNext_28_0_load_store_27;
  reg                 io_in_r_bypass_regNext_28_0_df_is_ws_27;
  reg                 io_in_r_bypass_regNext_28_0_stall_27;
  reg        [15:0]   io_in_r_bypass_regNext_28_1_data_27;
  reg                 io_in_r_bypass_regNext_28_1_load_store_27;
  reg                 io_in_r_bypass_regNext_28_1_df_is_ws_27;
  reg                 io_in_r_bypass_regNext_28_1_stall_27;
  reg        [15:0]   io_in_r_bypass_regNext_28_2_data_27;
  reg                 io_in_r_bypass_regNext_28_2_load_store_27;
  reg                 io_in_r_bypass_regNext_28_2_df_is_ws_27;
  reg                 io_in_r_bypass_regNext_28_2_stall_27;
  reg        [15:0]   io_in_r_bypass_regNext_28_3_data_27;
  reg                 io_in_r_bypass_regNext_28_3_load_store_27;
  reg                 io_in_r_bypass_regNext_28_3_df_is_ws_27;
  reg                 io_in_r_bypass_regNext_28_3_stall_27;
  reg        [15:0]   io_in_r_bypass_regNext_29_0_data_27;
  reg                 io_in_r_bypass_regNext_29_0_load_store_27;
  reg                 io_in_r_bypass_regNext_29_0_df_is_ws_27;
  reg                 io_in_r_bypass_regNext_29_0_stall_27;
  reg        [15:0]   io_in_r_bypass_regNext_29_1_data_27;
  reg                 io_in_r_bypass_regNext_29_1_load_store_27;
  reg                 io_in_r_bypass_regNext_29_1_df_is_ws_27;
  reg                 io_in_r_bypass_regNext_29_1_stall_27;
  reg        [15:0]   io_in_r_bypass_regNext_29_2_data_27;
  reg                 io_in_r_bypass_regNext_29_2_load_store_27;
  reg                 io_in_r_bypass_regNext_29_2_df_is_ws_27;
  reg                 io_in_r_bypass_regNext_29_2_stall_27;
  reg        [15:0]   io_in_r_bypass_regNext_29_3_data_27;
  reg                 io_in_r_bypass_regNext_29_3_load_store_27;
  reg                 io_in_r_bypass_regNext_29_3_df_is_ws_27;
  reg                 io_in_r_bypass_regNext_29_3_stall_27;
  reg        [15:0]   io_in_r_bypass_regNext_30_0_data_27;
  reg                 io_in_r_bypass_regNext_30_0_load_store_27;
  reg                 io_in_r_bypass_regNext_30_0_df_is_ws_27;
  reg                 io_in_r_bypass_regNext_30_0_stall_27;
  reg        [15:0]   io_in_r_bypass_regNext_30_1_data_27;
  reg                 io_in_r_bypass_regNext_30_1_load_store_27;
  reg                 io_in_r_bypass_regNext_30_1_df_is_ws_27;
  reg                 io_in_r_bypass_regNext_30_1_stall_27;
  reg        [15:0]   io_in_r_bypass_regNext_30_2_data_27;
  reg                 io_in_r_bypass_regNext_30_2_load_store_27;
  reg                 io_in_r_bypass_regNext_30_2_df_is_ws_27;
  reg                 io_in_r_bypass_regNext_30_2_stall_27;
  reg        [15:0]   io_in_r_bypass_regNext_30_3_data_27;
  reg                 io_in_r_bypass_regNext_30_3_load_store_27;
  reg                 io_in_r_bypass_regNext_30_3_df_is_ws_27;
  reg                 io_in_r_bypass_regNext_30_3_stall_27;
  reg        [15:0]   io_in_r_bypass_regNext_31_0_data_27;
  reg                 io_in_r_bypass_regNext_31_0_load_store_27;
  reg                 io_in_r_bypass_regNext_31_0_df_is_ws_27;
  reg                 io_in_r_bypass_regNext_31_0_stall_27;
  reg        [15:0]   io_in_r_bypass_regNext_31_1_data_27;
  reg                 io_in_r_bypass_regNext_31_1_load_store_27;
  reg                 io_in_r_bypass_regNext_31_1_df_is_ws_27;
  reg                 io_in_r_bypass_regNext_31_1_stall_27;
  reg        [15:0]   io_in_r_bypass_regNext_31_2_data_27;
  reg                 io_in_r_bypass_regNext_31_2_load_store_27;
  reg                 io_in_r_bypass_regNext_31_2_df_is_ws_27;
  reg                 io_in_r_bypass_regNext_31_2_stall_27;
  reg        [15:0]   io_in_r_bypass_regNext_31_3_data_27;
  reg                 io_in_r_bypass_regNext_31_3_load_store_27;
  reg                 io_in_r_bypass_regNext_31_3_df_is_ws_27;
  reg                 io_in_r_bypass_regNext_31_3_stall_27;
  reg        [15:0]   io_in_r_bypass_regNext_0_0_data_28;
  reg                 io_in_r_bypass_regNext_0_0_load_store_28;
  reg                 io_in_r_bypass_regNext_0_0_df_is_ws_28;
  reg                 io_in_r_bypass_regNext_0_0_stall_28;
  reg        [15:0]   io_in_r_bypass_regNext_0_1_data_28;
  reg                 io_in_r_bypass_regNext_0_1_load_store_28;
  reg                 io_in_r_bypass_regNext_0_1_df_is_ws_28;
  reg                 io_in_r_bypass_regNext_0_1_stall_28;
  reg        [15:0]   io_in_r_bypass_regNext_0_2_data_28;
  reg                 io_in_r_bypass_regNext_0_2_load_store_28;
  reg                 io_in_r_bypass_regNext_0_2_df_is_ws_28;
  reg                 io_in_r_bypass_regNext_0_2_stall_28;
  reg        [15:0]   io_in_r_bypass_regNext_0_3_data_28;
  reg                 io_in_r_bypass_regNext_0_3_load_store_28;
  reg                 io_in_r_bypass_regNext_0_3_df_is_ws_28;
  reg                 io_in_r_bypass_regNext_0_3_stall_28;
  reg        [15:0]   io_in_r_bypass_regNext_1_0_data_28;
  reg                 io_in_r_bypass_regNext_1_0_load_store_28;
  reg                 io_in_r_bypass_regNext_1_0_df_is_ws_28;
  reg                 io_in_r_bypass_regNext_1_0_stall_28;
  reg        [15:0]   io_in_r_bypass_regNext_1_1_data_28;
  reg                 io_in_r_bypass_regNext_1_1_load_store_28;
  reg                 io_in_r_bypass_regNext_1_1_df_is_ws_28;
  reg                 io_in_r_bypass_regNext_1_1_stall_28;
  reg        [15:0]   io_in_r_bypass_regNext_1_2_data_28;
  reg                 io_in_r_bypass_regNext_1_2_load_store_28;
  reg                 io_in_r_bypass_regNext_1_2_df_is_ws_28;
  reg                 io_in_r_bypass_regNext_1_2_stall_28;
  reg        [15:0]   io_in_r_bypass_regNext_1_3_data_28;
  reg                 io_in_r_bypass_regNext_1_3_load_store_28;
  reg                 io_in_r_bypass_regNext_1_3_df_is_ws_28;
  reg                 io_in_r_bypass_regNext_1_3_stall_28;
  reg        [15:0]   io_in_r_bypass_regNext_2_0_data_28;
  reg                 io_in_r_bypass_regNext_2_0_load_store_28;
  reg                 io_in_r_bypass_regNext_2_0_df_is_ws_28;
  reg                 io_in_r_bypass_regNext_2_0_stall_28;
  reg        [15:0]   io_in_r_bypass_regNext_2_1_data_28;
  reg                 io_in_r_bypass_regNext_2_1_load_store_28;
  reg                 io_in_r_bypass_regNext_2_1_df_is_ws_28;
  reg                 io_in_r_bypass_regNext_2_1_stall_28;
  reg        [15:0]   io_in_r_bypass_regNext_2_2_data_28;
  reg                 io_in_r_bypass_regNext_2_2_load_store_28;
  reg                 io_in_r_bypass_regNext_2_2_df_is_ws_28;
  reg                 io_in_r_bypass_regNext_2_2_stall_28;
  reg        [15:0]   io_in_r_bypass_regNext_2_3_data_28;
  reg                 io_in_r_bypass_regNext_2_3_load_store_28;
  reg                 io_in_r_bypass_regNext_2_3_df_is_ws_28;
  reg                 io_in_r_bypass_regNext_2_3_stall_28;
  reg        [15:0]   io_in_r_bypass_regNext_3_0_data_28;
  reg                 io_in_r_bypass_regNext_3_0_load_store_28;
  reg                 io_in_r_bypass_regNext_3_0_df_is_ws_28;
  reg                 io_in_r_bypass_regNext_3_0_stall_28;
  reg        [15:0]   io_in_r_bypass_regNext_3_1_data_28;
  reg                 io_in_r_bypass_regNext_3_1_load_store_28;
  reg                 io_in_r_bypass_regNext_3_1_df_is_ws_28;
  reg                 io_in_r_bypass_regNext_3_1_stall_28;
  reg        [15:0]   io_in_r_bypass_regNext_3_2_data_28;
  reg                 io_in_r_bypass_regNext_3_2_load_store_28;
  reg                 io_in_r_bypass_regNext_3_2_df_is_ws_28;
  reg                 io_in_r_bypass_regNext_3_2_stall_28;
  reg        [15:0]   io_in_r_bypass_regNext_3_3_data_28;
  reg                 io_in_r_bypass_regNext_3_3_load_store_28;
  reg                 io_in_r_bypass_regNext_3_3_df_is_ws_28;
  reg                 io_in_r_bypass_regNext_3_3_stall_28;
  reg        [15:0]   io_in_r_bypass_regNext_4_0_data_28;
  reg                 io_in_r_bypass_regNext_4_0_load_store_28;
  reg                 io_in_r_bypass_regNext_4_0_df_is_ws_28;
  reg                 io_in_r_bypass_regNext_4_0_stall_28;
  reg        [15:0]   io_in_r_bypass_regNext_4_1_data_28;
  reg                 io_in_r_bypass_regNext_4_1_load_store_28;
  reg                 io_in_r_bypass_regNext_4_1_df_is_ws_28;
  reg                 io_in_r_bypass_regNext_4_1_stall_28;
  reg        [15:0]   io_in_r_bypass_regNext_4_2_data_28;
  reg                 io_in_r_bypass_regNext_4_2_load_store_28;
  reg                 io_in_r_bypass_regNext_4_2_df_is_ws_28;
  reg                 io_in_r_bypass_regNext_4_2_stall_28;
  reg        [15:0]   io_in_r_bypass_regNext_4_3_data_28;
  reg                 io_in_r_bypass_regNext_4_3_load_store_28;
  reg                 io_in_r_bypass_regNext_4_3_df_is_ws_28;
  reg                 io_in_r_bypass_regNext_4_3_stall_28;
  reg        [15:0]   io_in_r_bypass_regNext_5_0_data_28;
  reg                 io_in_r_bypass_regNext_5_0_load_store_28;
  reg                 io_in_r_bypass_regNext_5_0_df_is_ws_28;
  reg                 io_in_r_bypass_regNext_5_0_stall_28;
  reg        [15:0]   io_in_r_bypass_regNext_5_1_data_28;
  reg                 io_in_r_bypass_regNext_5_1_load_store_28;
  reg                 io_in_r_bypass_regNext_5_1_df_is_ws_28;
  reg                 io_in_r_bypass_regNext_5_1_stall_28;
  reg        [15:0]   io_in_r_bypass_regNext_5_2_data_28;
  reg                 io_in_r_bypass_regNext_5_2_load_store_28;
  reg                 io_in_r_bypass_regNext_5_2_df_is_ws_28;
  reg                 io_in_r_bypass_regNext_5_2_stall_28;
  reg        [15:0]   io_in_r_bypass_regNext_5_3_data_28;
  reg                 io_in_r_bypass_regNext_5_3_load_store_28;
  reg                 io_in_r_bypass_regNext_5_3_df_is_ws_28;
  reg                 io_in_r_bypass_regNext_5_3_stall_28;
  reg        [15:0]   io_in_r_bypass_regNext_6_0_data_28;
  reg                 io_in_r_bypass_regNext_6_0_load_store_28;
  reg                 io_in_r_bypass_regNext_6_0_df_is_ws_28;
  reg                 io_in_r_bypass_regNext_6_0_stall_28;
  reg        [15:0]   io_in_r_bypass_regNext_6_1_data_28;
  reg                 io_in_r_bypass_regNext_6_1_load_store_28;
  reg                 io_in_r_bypass_regNext_6_1_df_is_ws_28;
  reg                 io_in_r_bypass_regNext_6_1_stall_28;
  reg        [15:0]   io_in_r_bypass_regNext_6_2_data_28;
  reg                 io_in_r_bypass_regNext_6_2_load_store_28;
  reg                 io_in_r_bypass_regNext_6_2_df_is_ws_28;
  reg                 io_in_r_bypass_regNext_6_2_stall_28;
  reg        [15:0]   io_in_r_bypass_regNext_6_3_data_28;
  reg                 io_in_r_bypass_regNext_6_3_load_store_28;
  reg                 io_in_r_bypass_regNext_6_3_df_is_ws_28;
  reg                 io_in_r_bypass_regNext_6_3_stall_28;
  reg        [15:0]   io_in_r_bypass_regNext_7_0_data_28;
  reg                 io_in_r_bypass_regNext_7_0_load_store_28;
  reg                 io_in_r_bypass_regNext_7_0_df_is_ws_28;
  reg                 io_in_r_bypass_regNext_7_0_stall_28;
  reg        [15:0]   io_in_r_bypass_regNext_7_1_data_28;
  reg                 io_in_r_bypass_regNext_7_1_load_store_28;
  reg                 io_in_r_bypass_regNext_7_1_df_is_ws_28;
  reg                 io_in_r_bypass_regNext_7_1_stall_28;
  reg        [15:0]   io_in_r_bypass_regNext_7_2_data_28;
  reg                 io_in_r_bypass_regNext_7_2_load_store_28;
  reg                 io_in_r_bypass_regNext_7_2_df_is_ws_28;
  reg                 io_in_r_bypass_regNext_7_2_stall_28;
  reg        [15:0]   io_in_r_bypass_regNext_7_3_data_28;
  reg                 io_in_r_bypass_regNext_7_3_load_store_28;
  reg                 io_in_r_bypass_regNext_7_3_df_is_ws_28;
  reg                 io_in_r_bypass_regNext_7_3_stall_28;
  reg        [15:0]   io_in_r_bypass_regNext_8_0_data_28;
  reg                 io_in_r_bypass_regNext_8_0_load_store_28;
  reg                 io_in_r_bypass_regNext_8_0_df_is_ws_28;
  reg                 io_in_r_bypass_regNext_8_0_stall_28;
  reg        [15:0]   io_in_r_bypass_regNext_8_1_data_28;
  reg                 io_in_r_bypass_regNext_8_1_load_store_28;
  reg                 io_in_r_bypass_regNext_8_1_df_is_ws_28;
  reg                 io_in_r_bypass_regNext_8_1_stall_28;
  reg        [15:0]   io_in_r_bypass_regNext_8_2_data_28;
  reg                 io_in_r_bypass_regNext_8_2_load_store_28;
  reg                 io_in_r_bypass_regNext_8_2_df_is_ws_28;
  reg                 io_in_r_bypass_regNext_8_2_stall_28;
  reg        [15:0]   io_in_r_bypass_regNext_8_3_data_28;
  reg                 io_in_r_bypass_regNext_8_3_load_store_28;
  reg                 io_in_r_bypass_regNext_8_3_df_is_ws_28;
  reg                 io_in_r_bypass_regNext_8_3_stall_28;
  reg        [15:0]   io_in_r_bypass_regNext_9_0_data_28;
  reg                 io_in_r_bypass_regNext_9_0_load_store_28;
  reg                 io_in_r_bypass_regNext_9_0_df_is_ws_28;
  reg                 io_in_r_bypass_regNext_9_0_stall_28;
  reg        [15:0]   io_in_r_bypass_regNext_9_1_data_28;
  reg                 io_in_r_bypass_regNext_9_1_load_store_28;
  reg                 io_in_r_bypass_regNext_9_1_df_is_ws_28;
  reg                 io_in_r_bypass_regNext_9_1_stall_28;
  reg        [15:0]   io_in_r_bypass_regNext_9_2_data_28;
  reg                 io_in_r_bypass_regNext_9_2_load_store_28;
  reg                 io_in_r_bypass_regNext_9_2_df_is_ws_28;
  reg                 io_in_r_bypass_regNext_9_2_stall_28;
  reg        [15:0]   io_in_r_bypass_regNext_9_3_data_28;
  reg                 io_in_r_bypass_regNext_9_3_load_store_28;
  reg                 io_in_r_bypass_regNext_9_3_df_is_ws_28;
  reg                 io_in_r_bypass_regNext_9_3_stall_28;
  reg        [15:0]   io_in_r_bypass_regNext_10_0_data_28;
  reg                 io_in_r_bypass_regNext_10_0_load_store_28;
  reg                 io_in_r_bypass_regNext_10_0_df_is_ws_28;
  reg                 io_in_r_bypass_regNext_10_0_stall_28;
  reg        [15:0]   io_in_r_bypass_regNext_10_1_data_28;
  reg                 io_in_r_bypass_regNext_10_1_load_store_28;
  reg                 io_in_r_bypass_regNext_10_1_df_is_ws_28;
  reg                 io_in_r_bypass_regNext_10_1_stall_28;
  reg        [15:0]   io_in_r_bypass_regNext_10_2_data_28;
  reg                 io_in_r_bypass_regNext_10_2_load_store_28;
  reg                 io_in_r_bypass_regNext_10_2_df_is_ws_28;
  reg                 io_in_r_bypass_regNext_10_2_stall_28;
  reg        [15:0]   io_in_r_bypass_regNext_10_3_data_28;
  reg                 io_in_r_bypass_regNext_10_3_load_store_28;
  reg                 io_in_r_bypass_regNext_10_3_df_is_ws_28;
  reg                 io_in_r_bypass_regNext_10_3_stall_28;
  reg        [15:0]   io_in_r_bypass_regNext_11_0_data_28;
  reg                 io_in_r_bypass_regNext_11_0_load_store_28;
  reg                 io_in_r_bypass_regNext_11_0_df_is_ws_28;
  reg                 io_in_r_bypass_regNext_11_0_stall_28;
  reg        [15:0]   io_in_r_bypass_regNext_11_1_data_28;
  reg                 io_in_r_bypass_regNext_11_1_load_store_28;
  reg                 io_in_r_bypass_regNext_11_1_df_is_ws_28;
  reg                 io_in_r_bypass_regNext_11_1_stall_28;
  reg        [15:0]   io_in_r_bypass_regNext_11_2_data_28;
  reg                 io_in_r_bypass_regNext_11_2_load_store_28;
  reg                 io_in_r_bypass_regNext_11_2_df_is_ws_28;
  reg                 io_in_r_bypass_regNext_11_2_stall_28;
  reg        [15:0]   io_in_r_bypass_regNext_11_3_data_28;
  reg                 io_in_r_bypass_regNext_11_3_load_store_28;
  reg                 io_in_r_bypass_regNext_11_3_df_is_ws_28;
  reg                 io_in_r_bypass_regNext_11_3_stall_28;
  reg        [15:0]   io_in_r_bypass_regNext_12_0_data_28;
  reg                 io_in_r_bypass_regNext_12_0_load_store_28;
  reg                 io_in_r_bypass_regNext_12_0_df_is_ws_28;
  reg                 io_in_r_bypass_regNext_12_0_stall_28;
  reg        [15:0]   io_in_r_bypass_regNext_12_1_data_28;
  reg                 io_in_r_bypass_regNext_12_1_load_store_28;
  reg                 io_in_r_bypass_regNext_12_1_df_is_ws_28;
  reg                 io_in_r_bypass_regNext_12_1_stall_28;
  reg        [15:0]   io_in_r_bypass_regNext_12_2_data_28;
  reg                 io_in_r_bypass_regNext_12_2_load_store_28;
  reg                 io_in_r_bypass_regNext_12_2_df_is_ws_28;
  reg                 io_in_r_bypass_regNext_12_2_stall_28;
  reg        [15:0]   io_in_r_bypass_regNext_12_3_data_28;
  reg                 io_in_r_bypass_regNext_12_3_load_store_28;
  reg                 io_in_r_bypass_regNext_12_3_df_is_ws_28;
  reg                 io_in_r_bypass_regNext_12_3_stall_28;
  reg        [15:0]   io_in_r_bypass_regNext_13_0_data_28;
  reg                 io_in_r_bypass_regNext_13_0_load_store_28;
  reg                 io_in_r_bypass_regNext_13_0_df_is_ws_28;
  reg                 io_in_r_bypass_regNext_13_0_stall_28;
  reg        [15:0]   io_in_r_bypass_regNext_13_1_data_28;
  reg                 io_in_r_bypass_regNext_13_1_load_store_28;
  reg                 io_in_r_bypass_regNext_13_1_df_is_ws_28;
  reg                 io_in_r_bypass_regNext_13_1_stall_28;
  reg        [15:0]   io_in_r_bypass_regNext_13_2_data_28;
  reg                 io_in_r_bypass_regNext_13_2_load_store_28;
  reg                 io_in_r_bypass_regNext_13_2_df_is_ws_28;
  reg                 io_in_r_bypass_regNext_13_2_stall_28;
  reg        [15:0]   io_in_r_bypass_regNext_13_3_data_28;
  reg                 io_in_r_bypass_regNext_13_3_load_store_28;
  reg                 io_in_r_bypass_regNext_13_3_df_is_ws_28;
  reg                 io_in_r_bypass_regNext_13_3_stall_28;
  reg        [15:0]   io_in_r_bypass_regNext_14_0_data_28;
  reg                 io_in_r_bypass_regNext_14_0_load_store_28;
  reg                 io_in_r_bypass_regNext_14_0_df_is_ws_28;
  reg                 io_in_r_bypass_regNext_14_0_stall_28;
  reg        [15:0]   io_in_r_bypass_regNext_14_1_data_28;
  reg                 io_in_r_bypass_regNext_14_1_load_store_28;
  reg                 io_in_r_bypass_regNext_14_1_df_is_ws_28;
  reg                 io_in_r_bypass_regNext_14_1_stall_28;
  reg        [15:0]   io_in_r_bypass_regNext_14_2_data_28;
  reg                 io_in_r_bypass_regNext_14_2_load_store_28;
  reg                 io_in_r_bypass_regNext_14_2_df_is_ws_28;
  reg                 io_in_r_bypass_regNext_14_2_stall_28;
  reg        [15:0]   io_in_r_bypass_regNext_14_3_data_28;
  reg                 io_in_r_bypass_regNext_14_3_load_store_28;
  reg                 io_in_r_bypass_regNext_14_3_df_is_ws_28;
  reg                 io_in_r_bypass_regNext_14_3_stall_28;
  reg        [15:0]   io_in_r_bypass_regNext_15_0_data_28;
  reg                 io_in_r_bypass_regNext_15_0_load_store_28;
  reg                 io_in_r_bypass_regNext_15_0_df_is_ws_28;
  reg                 io_in_r_bypass_regNext_15_0_stall_28;
  reg        [15:0]   io_in_r_bypass_regNext_15_1_data_28;
  reg                 io_in_r_bypass_regNext_15_1_load_store_28;
  reg                 io_in_r_bypass_regNext_15_1_df_is_ws_28;
  reg                 io_in_r_bypass_regNext_15_1_stall_28;
  reg        [15:0]   io_in_r_bypass_regNext_15_2_data_28;
  reg                 io_in_r_bypass_regNext_15_2_load_store_28;
  reg                 io_in_r_bypass_regNext_15_2_df_is_ws_28;
  reg                 io_in_r_bypass_regNext_15_2_stall_28;
  reg        [15:0]   io_in_r_bypass_regNext_15_3_data_28;
  reg                 io_in_r_bypass_regNext_15_3_load_store_28;
  reg                 io_in_r_bypass_regNext_15_3_df_is_ws_28;
  reg                 io_in_r_bypass_regNext_15_3_stall_28;
  reg        [15:0]   io_in_r_bypass_regNext_16_0_data_28;
  reg                 io_in_r_bypass_regNext_16_0_load_store_28;
  reg                 io_in_r_bypass_regNext_16_0_df_is_ws_28;
  reg                 io_in_r_bypass_regNext_16_0_stall_28;
  reg        [15:0]   io_in_r_bypass_regNext_16_1_data_28;
  reg                 io_in_r_bypass_regNext_16_1_load_store_28;
  reg                 io_in_r_bypass_regNext_16_1_df_is_ws_28;
  reg                 io_in_r_bypass_regNext_16_1_stall_28;
  reg        [15:0]   io_in_r_bypass_regNext_16_2_data_28;
  reg                 io_in_r_bypass_regNext_16_2_load_store_28;
  reg                 io_in_r_bypass_regNext_16_2_df_is_ws_28;
  reg                 io_in_r_bypass_regNext_16_2_stall_28;
  reg        [15:0]   io_in_r_bypass_regNext_16_3_data_28;
  reg                 io_in_r_bypass_regNext_16_3_load_store_28;
  reg                 io_in_r_bypass_regNext_16_3_df_is_ws_28;
  reg                 io_in_r_bypass_regNext_16_3_stall_28;
  reg        [15:0]   io_in_r_bypass_regNext_17_0_data_28;
  reg                 io_in_r_bypass_regNext_17_0_load_store_28;
  reg                 io_in_r_bypass_regNext_17_0_df_is_ws_28;
  reg                 io_in_r_bypass_regNext_17_0_stall_28;
  reg        [15:0]   io_in_r_bypass_regNext_17_1_data_28;
  reg                 io_in_r_bypass_regNext_17_1_load_store_28;
  reg                 io_in_r_bypass_regNext_17_1_df_is_ws_28;
  reg                 io_in_r_bypass_regNext_17_1_stall_28;
  reg        [15:0]   io_in_r_bypass_regNext_17_2_data_28;
  reg                 io_in_r_bypass_regNext_17_2_load_store_28;
  reg                 io_in_r_bypass_regNext_17_2_df_is_ws_28;
  reg                 io_in_r_bypass_regNext_17_2_stall_28;
  reg        [15:0]   io_in_r_bypass_regNext_17_3_data_28;
  reg                 io_in_r_bypass_regNext_17_3_load_store_28;
  reg                 io_in_r_bypass_regNext_17_3_df_is_ws_28;
  reg                 io_in_r_bypass_regNext_17_3_stall_28;
  reg        [15:0]   io_in_r_bypass_regNext_18_0_data_28;
  reg                 io_in_r_bypass_regNext_18_0_load_store_28;
  reg                 io_in_r_bypass_regNext_18_0_df_is_ws_28;
  reg                 io_in_r_bypass_regNext_18_0_stall_28;
  reg        [15:0]   io_in_r_bypass_regNext_18_1_data_28;
  reg                 io_in_r_bypass_regNext_18_1_load_store_28;
  reg                 io_in_r_bypass_regNext_18_1_df_is_ws_28;
  reg                 io_in_r_bypass_regNext_18_1_stall_28;
  reg        [15:0]   io_in_r_bypass_regNext_18_2_data_28;
  reg                 io_in_r_bypass_regNext_18_2_load_store_28;
  reg                 io_in_r_bypass_regNext_18_2_df_is_ws_28;
  reg                 io_in_r_bypass_regNext_18_2_stall_28;
  reg        [15:0]   io_in_r_bypass_regNext_18_3_data_28;
  reg                 io_in_r_bypass_regNext_18_3_load_store_28;
  reg                 io_in_r_bypass_regNext_18_3_df_is_ws_28;
  reg                 io_in_r_bypass_regNext_18_3_stall_28;
  reg        [15:0]   io_in_r_bypass_regNext_19_0_data_28;
  reg                 io_in_r_bypass_regNext_19_0_load_store_28;
  reg                 io_in_r_bypass_regNext_19_0_df_is_ws_28;
  reg                 io_in_r_bypass_regNext_19_0_stall_28;
  reg        [15:0]   io_in_r_bypass_regNext_19_1_data_28;
  reg                 io_in_r_bypass_regNext_19_1_load_store_28;
  reg                 io_in_r_bypass_regNext_19_1_df_is_ws_28;
  reg                 io_in_r_bypass_regNext_19_1_stall_28;
  reg        [15:0]   io_in_r_bypass_regNext_19_2_data_28;
  reg                 io_in_r_bypass_regNext_19_2_load_store_28;
  reg                 io_in_r_bypass_regNext_19_2_df_is_ws_28;
  reg                 io_in_r_bypass_regNext_19_2_stall_28;
  reg        [15:0]   io_in_r_bypass_regNext_19_3_data_28;
  reg                 io_in_r_bypass_regNext_19_3_load_store_28;
  reg                 io_in_r_bypass_regNext_19_3_df_is_ws_28;
  reg                 io_in_r_bypass_regNext_19_3_stall_28;
  reg        [15:0]   io_in_r_bypass_regNext_20_0_data_28;
  reg                 io_in_r_bypass_regNext_20_0_load_store_28;
  reg                 io_in_r_bypass_regNext_20_0_df_is_ws_28;
  reg                 io_in_r_bypass_regNext_20_0_stall_28;
  reg        [15:0]   io_in_r_bypass_regNext_20_1_data_28;
  reg                 io_in_r_bypass_regNext_20_1_load_store_28;
  reg                 io_in_r_bypass_regNext_20_1_df_is_ws_28;
  reg                 io_in_r_bypass_regNext_20_1_stall_28;
  reg        [15:0]   io_in_r_bypass_regNext_20_2_data_28;
  reg                 io_in_r_bypass_regNext_20_2_load_store_28;
  reg                 io_in_r_bypass_regNext_20_2_df_is_ws_28;
  reg                 io_in_r_bypass_regNext_20_2_stall_28;
  reg        [15:0]   io_in_r_bypass_regNext_20_3_data_28;
  reg                 io_in_r_bypass_regNext_20_3_load_store_28;
  reg                 io_in_r_bypass_regNext_20_3_df_is_ws_28;
  reg                 io_in_r_bypass_regNext_20_3_stall_28;
  reg        [15:0]   io_in_r_bypass_regNext_21_0_data_28;
  reg                 io_in_r_bypass_regNext_21_0_load_store_28;
  reg                 io_in_r_bypass_regNext_21_0_df_is_ws_28;
  reg                 io_in_r_bypass_regNext_21_0_stall_28;
  reg        [15:0]   io_in_r_bypass_regNext_21_1_data_28;
  reg                 io_in_r_bypass_regNext_21_1_load_store_28;
  reg                 io_in_r_bypass_regNext_21_1_df_is_ws_28;
  reg                 io_in_r_bypass_regNext_21_1_stall_28;
  reg        [15:0]   io_in_r_bypass_regNext_21_2_data_28;
  reg                 io_in_r_bypass_regNext_21_2_load_store_28;
  reg                 io_in_r_bypass_regNext_21_2_df_is_ws_28;
  reg                 io_in_r_bypass_regNext_21_2_stall_28;
  reg        [15:0]   io_in_r_bypass_regNext_21_3_data_28;
  reg                 io_in_r_bypass_regNext_21_3_load_store_28;
  reg                 io_in_r_bypass_regNext_21_3_df_is_ws_28;
  reg                 io_in_r_bypass_regNext_21_3_stall_28;
  reg        [15:0]   io_in_r_bypass_regNext_22_0_data_28;
  reg                 io_in_r_bypass_regNext_22_0_load_store_28;
  reg                 io_in_r_bypass_regNext_22_0_df_is_ws_28;
  reg                 io_in_r_bypass_regNext_22_0_stall_28;
  reg        [15:0]   io_in_r_bypass_regNext_22_1_data_28;
  reg                 io_in_r_bypass_regNext_22_1_load_store_28;
  reg                 io_in_r_bypass_regNext_22_1_df_is_ws_28;
  reg                 io_in_r_bypass_regNext_22_1_stall_28;
  reg        [15:0]   io_in_r_bypass_regNext_22_2_data_28;
  reg                 io_in_r_bypass_regNext_22_2_load_store_28;
  reg                 io_in_r_bypass_regNext_22_2_df_is_ws_28;
  reg                 io_in_r_bypass_regNext_22_2_stall_28;
  reg        [15:0]   io_in_r_bypass_regNext_22_3_data_28;
  reg                 io_in_r_bypass_regNext_22_3_load_store_28;
  reg                 io_in_r_bypass_regNext_22_3_df_is_ws_28;
  reg                 io_in_r_bypass_regNext_22_3_stall_28;
  reg        [15:0]   io_in_r_bypass_regNext_23_0_data_28;
  reg                 io_in_r_bypass_regNext_23_0_load_store_28;
  reg                 io_in_r_bypass_regNext_23_0_df_is_ws_28;
  reg                 io_in_r_bypass_regNext_23_0_stall_28;
  reg        [15:0]   io_in_r_bypass_regNext_23_1_data_28;
  reg                 io_in_r_bypass_regNext_23_1_load_store_28;
  reg                 io_in_r_bypass_regNext_23_1_df_is_ws_28;
  reg                 io_in_r_bypass_regNext_23_1_stall_28;
  reg        [15:0]   io_in_r_bypass_regNext_23_2_data_28;
  reg                 io_in_r_bypass_regNext_23_2_load_store_28;
  reg                 io_in_r_bypass_regNext_23_2_df_is_ws_28;
  reg                 io_in_r_bypass_regNext_23_2_stall_28;
  reg        [15:0]   io_in_r_bypass_regNext_23_3_data_28;
  reg                 io_in_r_bypass_regNext_23_3_load_store_28;
  reg                 io_in_r_bypass_regNext_23_3_df_is_ws_28;
  reg                 io_in_r_bypass_regNext_23_3_stall_28;
  reg        [15:0]   io_in_r_bypass_regNext_24_0_data_28;
  reg                 io_in_r_bypass_regNext_24_0_load_store_28;
  reg                 io_in_r_bypass_regNext_24_0_df_is_ws_28;
  reg                 io_in_r_bypass_regNext_24_0_stall_28;
  reg        [15:0]   io_in_r_bypass_regNext_24_1_data_28;
  reg                 io_in_r_bypass_regNext_24_1_load_store_28;
  reg                 io_in_r_bypass_regNext_24_1_df_is_ws_28;
  reg                 io_in_r_bypass_regNext_24_1_stall_28;
  reg        [15:0]   io_in_r_bypass_regNext_24_2_data_28;
  reg                 io_in_r_bypass_regNext_24_2_load_store_28;
  reg                 io_in_r_bypass_regNext_24_2_df_is_ws_28;
  reg                 io_in_r_bypass_regNext_24_2_stall_28;
  reg        [15:0]   io_in_r_bypass_regNext_24_3_data_28;
  reg                 io_in_r_bypass_regNext_24_3_load_store_28;
  reg                 io_in_r_bypass_regNext_24_3_df_is_ws_28;
  reg                 io_in_r_bypass_regNext_24_3_stall_28;
  reg        [15:0]   io_in_r_bypass_regNext_25_0_data_28;
  reg                 io_in_r_bypass_regNext_25_0_load_store_28;
  reg                 io_in_r_bypass_regNext_25_0_df_is_ws_28;
  reg                 io_in_r_bypass_regNext_25_0_stall_28;
  reg        [15:0]   io_in_r_bypass_regNext_25_1_data_28;
  reg                 io_in_r_bypass_regNext_25_1_load_store_28;
  reg                 io_in_r_bypass_regNext_25_1_df_is_ws_28;
  reg                 io_in_r_bypass_regNext_25_1_stall_28;
  reg        [15:0]   io_in_r_bypass_regNext_25_2_data_28;
  reg                 io_in_r_bypass_regNext_25_2_load_store_28;
  reg                 io_in_r_bypass_regNext_25_2_df_is_ws_28;
  reg                 io_in_r_bypass_regNext_25_2_stall_28;
  reg        [15:0]   io_in_r_bypass_regNext_25_3_data_28;
  reg                 io_in_r_bypass_regNext_25_3_load_store_28;
  reg                 io_in_r_bypass_regNext_25_3_df_is_ws_28;
  reg                 io_in_r_bypass_regNext_25_3_stall_28;
  reg        [15:0]   io_in_r_bypass_regNext_26_0_data_28;
  reg                 io_in_r_bypass_regNext_26_0_load_store_28;
  reg                 io_in_r_bypass_regNext_26_0_df_is_ws_28;
  reg                 io_in_r_bypass_regNext_26_0_stall_28;
  reg        [15:0]   io_in_r_bypass_regNext_26_1_data_28;
  reg                 io_in_r_bypass_regNext_26_1_load_store_28;
  reg                 io_in_r_bypass_regNext_26_1_df_is_ws_28;
  reg                 io_in_r_bypass_regNext_26_1_stall_28;
  reg        [15:0]   io_in_r_bypass_regNext_26_2_data_28;
  reg                 io_in_r_bypass_regNext_26_2_load_store_28;
  reg                 io_in_r_bypass_regNext_26_2_df_is_ws_28;
  reg                 io_in_r_bypass_regNext_26_2_stall_28;
  reg        [15:0]   io_in_r_bypass_regNext_26_3_data_28;
  reg                 io_in_r_bypass_regNext_26_3_load_store_28;
  reg                 io_in_r_bypass_regNext_26_3_df_is_ws_28;
  reg                 io_in_r_bypass_regNext_26_3_stall_28;
  reg        [15:0]   io_in_r_bypass_regNext_27_0_data_28;
  reg                 io_in_r_bypass_regNext_27_0_load_store_28;
  reg                 io_in_r_bypass_regNext_27_0_df_is_ws_28;
  reg                 io_in_r_bypass_regNext_27_0_stall_28;
  reg        [15:0]   io_in_r_bypass_regNext_27_1_data_28;
  reg                 io_in_r_bypass_regNext_27_1_load_store_28;
  reg                 io_in_r_bypass_regNext_27_1_df_is_ws_28;
  reg                 io_in_r_bypass_regNext_27_1_stall_28;
  reg        [15:0]   io_in_r_bypass_regNext_27_2_data_28;
  reg                 io_in_r_bypass_regNext_27_2_load_store_28;
  reg                 io_in_r_bypass_regNext_27_2_df_is_ws_28;
  reg                 io_in_r_bypass_regNext_27_2_stall_28;
  reg        [15:0]   io_in_r_bypass_regNext_27_3_data_28;
  reg                 io_in_r_bypass_regNext_27_3_load_store_28;
  reg                 io_in_r_bypass_regNext_27_3_df_is_ws_28;
  reg                 io_in_r_bypass_regNext_27_3_stall_28;
  reg        [15:0]   io_in_r_bypass_regNext_28_0_data_28;
  reg                 io_in_r_bypass_regNext_28_0_load_store_28;
  reg                 io_in_r_bypass_regNext_28_0_df_is_ws_28;
  reg                 io_in_r_bypass_regNext_28_0_stall_28;
  reg        [15:0]   io_in_r_bypass_regNext_28_1_data_28;
  reg                 io_in_r_bypass_regNext_28_1_load_store_28;
  reg                 io_in_r_bypass_regNext_28_1_df_is_ws_28;
  reg                 io_in_r_bypass_regNext_28_1_stall_28;
  reg        [15:0]   io_in_r_bypass_regNext_28_2_data_28;
  reg                 io_in_r_bypass_regNext_28_2_load_store_28;
  reg                 io_in_r_bypass_regNext_28_2_df_is_ws_28;
  reg                 io_in_r_bypass_regNext_28_2_stall_28;
  reg        [15:0]   io_in_r_bypass_regNext_28_3_data_28;
  reg                 io_in_r_bypass_regNext_28_3_load_store_28;
  reg                 io_in_r_bypass_regNext_28_3_df_is_ws_28;
  reg                 io_in_r_bypass_regNext_28_3_stall_28;
  reg        [15:0]   io_in_r_bypass_regNext_29_0_data_28;
  reg                 io_in_r_bypass_regNext_29_0_load_store_28;
  reg                 io_in_r_bypass_regNext_29_0_df_is_ws_28;
  reg                 io_in_r_bypass_regNext_29_0_stall_28;
  reg        [15:0]   io_in_r_bypass_regNext_29_1_data_28;
  reg                 io_in_r_bypass_regNext_29_1_load_store_28;
  reg                 io_in_r_bypass_regNext_29_1_df_is_ws_28;
  reg                 io_in_r_bypass_regNext_29_1_stall_28;
  reg        [15:0]   io_in_r_bypass_regNext_29_2_data_28;
  reg                 io_in_r_bypass_regNext_29_2_load_store_28;
  reg                 io_in_r_bypass_regNext_29_2_df_is_ws_28;
  reg                 io_in_r_bypass_regNext_29_2_stall_28;
  reg        [15:0]   io_in_r_bypass_regNext_29_3_data_28;
  reg                 io_in_r_bypass_regNext_29_3_load_store_28;
  reg                 io_in_r_bypass_regNext_29_3_df_is_ws_28;
  reg                 io_in_r_bypass_regNext_29_3_stall_28;
  reg        [15:0]   io_in_r_bypass_regNext_30_0_data_28;
  reg                 io_in_r_bypass_regNext_30_0_load_store_28;
  reg                 io_in_r_bypass_regNext_30_0_df_is_ws_28;
  reg                 io_in_r_bypass_regNext_30_0_stall_28;
  reg        [15:0]   io_in_r_bypass_regNext_30_1_data_28;
  reg                 io_in_r_bypass_regNext_30_1_load_store_28;
  reg                 io_in_r_bypass_regNext_30_1_df_is_ws_28;
  reg                 io_in_r_bypass_regNext_30_1_stall_28;
  reg        [15:0]   io_in_r_bypass_regNext_30_2_data_28;
  reg                 io_in_r_bypass_regNext_30_2_load_store_28;
  reg                 io_in_r_bypass_regNext_30_2_df_is_ws_28;
  reg                 io_in_r_bypass_regNext_30_2_stall_28;
  reg        [15:0]   io_in_r_bypass_regNext_30_3_data_28;
  reg                 io_in_r_bypass_regNext_30_3_load_store_28;
  reg                 io_in_r_bypass_regNext_30_3_df_is_ws_28;
  reg                 io_in_r_bypass_regNext_30_3_stall_28;
  reg        [15:0]   io_in_r_bypass_regNext_31_0_data_28;
  reg                 io_in_r_bypass_regNext_31_0_load_store_28;
  reg                 io_in_r_bypass_regNext_31_0_df_is_ws_28;
  reg                 io_in_r_bypass_regNext_31_0_stall_28;
  reg        [15:0]   io_in_r_bypass_regNext_31_1_data_28;
  reg                 io_in_r_bypass_regNext_31_1_load_store_28;
  reg                 io_in_r_bypass_regNext_31_1_df_is_ws_28;
  reg                 io_in_r_bypass_regNext_31_1_stall_28;
  reg        [15:0]   io_in_r_bypass_regNext_31_2_data_28;
  reg                 io_in_r_bypass_regNext_31_2_load_store_28;
  reg                 io_in_r_bypass_regNext_31_2_df_is_ws_28;
  reg                 io_in_r_bypass_regNext_31_2_stall_28;
  reg        [15:0]   io_in_r_bypass_regNext_31_3_data_28;
  reg                 io_in_r_bypass_regNext_31_3_load_store_28;
  reg                 io_in_r_bypass_regNext_31_3_df_is_ws_28;
  reg                 io_in_r_bypass_regNext_31_3_stall_28;
  reg        [15:0]   io_in_r_bypass_regNext_0_0_data_29;
  reg                 io_in_r_bypass_regNext_0_0_load_store_29;
  reg                 io_in_r_bypass_regNext_0_0_df_is_ws_29;
  reg                 io_in_r_bypass_regNext_0_0_stall_29;
  reg        [15:0]   io_in_r_bypass_regNext_0_1_data_29;
  reg                 io_in_r_bypass_regNext_0_1_load_store_29;
  reg                 io_in_r_bypass_regNext_0_1_df_is_ws_29;
  reg                 io_in_r_bypass_regNext_0_1_stall_29;
  reg        [15:0]   io_in_r_bypass_regNext_0_2_data_29;
  reg                 io_in_r_bypass_regNext_0_2_load_store_29;
  reg                 io_in_r_bypass_regNext_0_2_df_is_ws_29;
  reg                 io_in_r_bypass_regNext_0_2_stall_29;
  reg        [15:0]   io_in_r_bypass_regNext_0_3_data_29;
  reg                 io_in_r_bypass_regNext_0_3_load_store_29;
  reg                 io_in_r_bypass_regNext_0_3_df_is_ws_29;
  reg                 io_in_r_bypass_regNext_0_3_stall_29;
  reg        [15:0]   io_in_r_bypass_regNext_1_0_data_29;
  reg                 io_in_r_bypass_regNext_1_0_load_store_29;
  reg                 io_in_r_bypass_regNext_1_0_df_is_ws_29;
  reg                 io_in_r_bypass_regNext_1_0_stall_29;
  reg        [15:0]   io_in_r_bypass_regNext_1_1_data_29;
  reg                 io_in_r_bypass_regNext_1_1_load_store_29;
  reg                 io_in_r_bypass_regNext_1_1_df_is_ws_29;
  reg                 io_in_r_bypass_regNext_1_1_stall_29;
  reg        [15:0]   io_in_r_bypass_regNext_1_2_data_29;
  reg                 io_in_r_bypass_regNext_1_2_load_store_29;
  reg                 io_in_r_bypass_regNext_1_2_df_is_ws_29;
  reg                 io_in_r_bypass_regNext_1_2_stall_29;
  reg        [15:0]   io_in_r_bypass_regNext_1_3_data_29;
  reg                 io_in_r_bypass_regNext_1_3_load_store_29;
  reg                 io_in_r_bypass_regNext_1_3_df_is_ws_29;
  reg                 io_in_r_bypass_regNext_1_3_stall_29;
  reg        [15:0]   io_in_r_bypass_regNext_2_0_data_29;
  reg                 io_in_r_bypass_regNext_2_0_load_store_29;
  reg                 io_in_r_bypass_regNext_2_0_df_is_ws_29;
  reg                 io_in_r_bypass_regNext_2_0_stall_29;
  reg        [15:0]   io_in_r_bypass_regNext_2_1_data_29;
  reg                 io_in_r_bypass_regNext_2_1_load_store_29;
  reg                 io_in_r_bypass_regNext_2_1_df_is_ws_29;
  reg                 io_in_r_bypass_regNext_2_1_stall_29;
  reg        [15:0]   io_in_r_bypass_regNext_2_2_data_29;
  reg                 io_in_r_bypass_regNext_2_2_load_store_29;
  reg                 io_in_r_bypass_regNext_2_2_df_is_ws_29;
  reg                 io_in_r_bypass_regNext_2_2_stall_29;
  reg        [15:0]   io_in_r_bypass_regNext_2_3_data_29;
  reg                 io_in_r_bypass_regNext_2_3_load_store_29;
  reg                 io_in_r_bypass_regNext_2_3_df_is_ws_29;
  reg                 io_in_r_bypass_regNext_2_3_stall_29;
  reg        [15:0]   io_in_r_bypass_regNext_3_0_data_29;
  reg                 io_in_r_bypass_regNext_3_0_load_store_29;
  reg                 io_in_r_bypass_regNext_3_0_df_is_ws_29;
  reg                 io_in_r_bypass_regNext_3_0_stall_29;
  reg        [15:0]   io_in_r_bypass_regNext_3_1_data_29;
  reg                 io_in_r_bypass_regNext_3_1_load_store_29;
  reg                 io_in_r_bypass_regNext_3_1_df_is_ws_29;
  reg                 io_in_r_bypass_regNext_3_1_stall_29;
  reg        [15:0]   io_in_r_bypass_regNext_3_2_data_29;
  reg                 io_in_r_bypass_regNext_3_2_load_store_29;
  reg                 io_in_r_bypass_regNext_3_2_df_is_ws_29;
  reg                 io_in_r_bypass_regNext_3_2_stall_29;
  reg        [15:0]   io_in_r_bypass_regNext_3_3_data_29;
  reg                 io_in_r_bypass_regNext_3_3_load_store_29;
  reg                 io_in_r_bypass_regNext_3_3_df_is_ws_29;
  reg                 io_in_r_bypass_regNext_3_3_stall_29;
  reg        [15:0]   io_in_r_bypass_regNext_4_0_data_29;
  reg                 io_in_r_bypass_regNext_4_0_load_store_29;
  reg                 io_in_r_bypass_regNext_4_0_df_is_ws_29;
  reg                 io_in_r_bypass_regNext_4_0_stall_29;
  reg        [15:0]   io_in_r_bypass_regNext_4_1_data_29;
  reg                 io_in_r_bypass_regNext_4_1_load_store_29;
  reg                 io_in_r_bypass_regNext_4_1_df_is_ws_29;
  reg                 io_in_r_bypass_regNext_4_1_stall_29;
  reg        [15:0]   io_in_r_bypass_regNext_4_2_data_29;
  reg                 io_in_r_bypass_regNext_4_2_load_store_29;
  reg                 io_in_r_bypass_regNext_4_2_df_is_ws_29;
  reg                 io_in_r_bypass_regNext_4_2_stall_29;
  reg        [15:0]   io_in_r_bypass_regNext_4_3_data_29;
  reg                 io_in_r_bypass_regNext_4_3_load_store_29;
  reg                 io_in_r_bypass_regNext_4_3_df_is_ws_29;
  reg                 io_in_r_bypass_regNext_4_3_stall_29;
  reg        [15:0]   io_in_r_bypass_regNext_5_0_data_29;
  reg                 io_in_r_bypass_regNext_5_0_load_store_29;
  reg                 io_in_r_bypass_regNext_5_0_df_is_ws_29;
  reg                 io_in_r_bypass_regNext_5_0_stall_29;
  reg        [15:0]   io_in_r_bypass_regNext_5_1_data_29;
  reg                 io_in_r_bypass_regNext_5_1_load_store_29;
  reg                 io_in_r_bypass_regNext_5_1_df_is_ws_29;
  reg                 io_in_r_bypass_regNext_5_1_stall_29;
  reg        [15:0]   io_in_r_bypass_regNext_5_2_data_29;
  reg                 io_in_r_bypass_regNext_5_2_load_store_29;
  reg                 io_in_r_bypass_regNext_5_2_df_is_ws_29;
  reg                 io_in_r_bypass_regNext_5_2_stall_29;
  reg        [15:0]   io_in_r_bypass_regNext_5_3_data_29;
  reg                 io_in_r_bypass_regNext_5_3_load_store_29;
  reg                 io_in_r_bypass_regNext_5_3_df_is_ws_29;
  reg                 io_in_r_bypass_regNext_5_3_stall_29;
  reg        [15:0]   io_in_r_bypass_regNext_6_0_data_29;
  reg                 io_in_r_bypass_regNext_6_0_load_store_29;
  reg                 io_in_r_bypass_regNext_6_0_df_is_ws_29;
  reg                 io_in_r_bypass_regNext_6_0_stall_29;
  reg        [15:0]   io_in_r_bypass_regNext_6_1_data_29;
  reg                 io_in_r_bypass_regNext_6_1_load_store_29;
  reg                 io_in_r_bypass_regNext_6_1_df_is_ws_29;
  reg                 io_in_r_bypass_regNext_6_1_stall_29;
  reg        [15:0]   io_in_r_bypass_regNext_6_2_data_29;
  reg                 io_in_r_bypass_regNext_6_2_load_store_29;
  reg                 io_in_r_bypass_regNext_6_2_df_is_ws_29;
  reg                 io_in_r_bypass_regNext_6_2_stall_29;
  reg        [15:0]   io_in_r_bypass_regNext_6_3_data_29;
  reg                 io_in_r_bypass_regNext_6_3_load_store_29;
  reg                 io_in_r_bypass_regNext_6_3_df_is_ws_29;
  reg                 io_in_r_bypass_regNext_6_3_stall_29;
  reg        [15:0]   io_in_r_bypass_regNext_7_0_data_29;
  reg                 io_in_r_bypass_regNext_7_0_load_store_29;
  reg                 io_in_r_bypass_regNext_7_0_df_is_ws_29;
  reg                 io_in_r_bypass_regNext_7_0_stall_29;
  reg        [15:0]   io_in_r_bypass_regNext_7_1_data_29;
  reg                 io_in_r_bypass_regNext_7_1_load_store_29;
  reg                 io_in_r_bypass_regNext_7_1_df_is_ws_29;
  reg                 io_in_r_bypass_regNext_7_1_stall_29;
  reg        [15:0]   io_in_r_bypass_regNext_7_2_data_29;
  reg                 io_in_r_bypass_regNext_7_2_load_store_29;
  reg                 io_in_r_bypass_regNext_7_2_df_is_ws_29;
  reg                 io_in_r_bypass_regNext_7_2_stall_29;
  reg        [15:0]   io_in_r_bypass_regNext_7_3_data_29;
  reg                 io_in_r_bypass_regNext_7_3_load_store_29;
  reg                 io_in_r_bypass_regNext_7_3_df_is_ws_29;
  reg                 io_in_r_bypass_regNext_7_3_stall_29;
  reg        [15:0]   io_in_r_bypass_regNext_8_0_data_29;
  reg                 io_in_r_bypass_regNext_8_0_load_store_29;
  reg                 io_in_r_bypass_regNext_8_0_df_is_ws_29;
  reg                 io_in_r_bypass_regNext_8_0_stall_29;
  reg        [15:0]   io_in_r_bypass_regNext_8_1_data_29;
  reg                 io_in_r_bypass_regNext_8_1_load_store_29;
  reg                 io_in_r_bypass_regNext_8_1_df_is_ws_29;
  reg                 io_in_r_bypass_regNext_8_1_stall_29;
  reg        [15:0]   io_in_r_bypass_regNext_8_2_data_29;
  reg                 io_in_r_bypass_regNext_8_2_load_store_29;
  reg                 io_in_r_bypass_regNext_8_2_df_is_ws_29;
  reg                 io_in_r_bypass_regNext_8_2_stall_29;
  reg        [15:0]   io_in_r_bypass_regNext_8_3_data_29;
  reg                 io_in_r_bypass_regNext_8_3_load_store_29;
  reg                 io_in_r_bypass_regNext_8_3_df_is_ws_29;
  reg                 io_in_r_bypass_regNext_8_3_stall_29;
  reg        [15:0]   io_in_r_bypass_regNext_9_0_data_29;
  reg                 io_in_r_bypass_regNext_9_0_load_store_29;
  reg                 io_in_r_bypass_regNext_9_0_df_is_ws_29;
  reg                 io_in_r_bypass_regNext_9_0_stall_29;
  reg        [15:0]   io_in_r_bypass_regNext_9_1_data_29;
  reg                 io_in_r_bypass_regNext_9_1_load_store_29;
  reg                 io_in_r_bypass_regNext_9_1_df_is_ws_29;
  reg                 io_in_r_bypass_regNext_9_1_stall_29;
  reg        [15:0]   io_in_r_bypass_regNext_9_2_data_29;
  reg                 io_in_r_bypass_regNext_9_2_load_store_29;
  reg                 io_in_r_bypass_regNext_9_2_df_is_ws_29;
  reg                 io_in_r_bypass_regNext_9_2_stall_29;
  reg        [15:0]   io_in_r_bypass_regNext_9_3_data_29;
  reg                 io_in_r_bypass_regNext_9_3_load_store_29;
  reg                 io_in_r_bypass_regNext_9_3_df_is_ws_29;
  reg                 io_in_r_bypass_regNext_9_3_stall_29;
  reg        [15:0]   io_in_r_bypass_regNext_10_0_data_29;
  reg                 io_in_r_bypass_regNext_10_0_load_store_29;
  reg                 io_in_r_bypass_regNext_10_0_df_is_ws_29;
  reg                 io_in_r_bypass_regNext_10_0_stall_29;
  reg        [15:0]   io_in_r_bypass_regNext_10_1_data_29;
  reg                 io_in_r_bypass_regNext_10_1_load_store_29;
  reg                 io_in_r_bypass_regNext_10_1_df_is_ws_29;
  reg                 io_in_r_bypass_regNext_10_1_stall_29;
  reg        [15:0]   io_in_r_bypass_regNext_10_2_data_29;
  reg                 io_in_r_bypass_regNext_10_2_load_store_29;
  reg                 io_in_r_bypass_regNext_10_2_df_is_ws_29;
  reg                 io_in_r_bypass_regNext_10_2_stall_29;
  reg        [15:0]   io_in_r_bypass_regNext_10_3_data_29;
  reg                 io_in_r_bypass_regNext_10_3_load_store_29;
  reg                 io_in_r_bypass_regNext_10_3_df_is_ws_29;
  reg                 io_in_r_bypass_regNext_10_3_stall_29;
  reg        [15:0]   io_in_r_bypass_regNext_11_0_data_29;
  reg                 io_in_r_bypass_regNext_11_0_load_store_29;
  reg                 io_in_r_bypass_regNext_11_0_df_is_ws_29;
  reg                 io_in_r_bypass_regNext_11_0_stall_29;
  reg        [15:0]   io_in_r_bypass_regNext_11_1_data_29;
  reg                 io_in_r_bypass_regNext_11_1_load_store_29;
  reg                 io_in_r_bypass_regNext_11_1_df_is_ws_29;
  reg                 io_in_r_bypass_regNext_11_1_stall_29;
  reg        [15:0]   io_in_r_bypass_regNext_11_2_data_29;
  reg                 io_in_r_bypass_regNext_11_2_load_store_29;
  reg                 io_in_r_bypass_regNext_11_2_df_is_ws_29;
  reg                 io_in_r_bypass_regNext_11_2_stall_29;
  reg        [15:0]   io_in_r_bypass_regNext_11_3_data_29;
  reg                 io_in_r_bypass_regNext_11_3_load_store_29;
  reg                 io_in_r_bypass_regNext_11_3_df_is_ws_29;
  reg                 io_in_r_bypass_regNext_11_3_stall_29;
  reg        [15:0]   io_in_r_bypass_regNext_12_0_data_29;
  reg                 io_in_r_bypass_regNext_12_0_load_store_29;
  reg                 io_in_r_bypass_regNext_12_0_df_is_ws_29;
  reg                 io_in_r_bypass_regNext_12_0_stall_29;
  reg        [15:0]   io_in_r_bypass_regNext_12_1_data_29;
  reg                 io_in_r_bypass_regNext_12_1_load_store_29;
  reg                 io_in_r_bypass_regNext_12_1_df_is_ws_29;
  reg                 io_in_r_bypass_regNext_12_1_stall_29;
  reg        [15:0]   io_in_r_bypass_regNext_12_2_data_29;
  reg                 io_in_r_bypass_regNext_12_2_load_store_29;
  reg                 io_in_r_bypass_regNext_12_2_df_is_ws_29;
  reg                 io_in_r_bypass_regNext_12_2_stall_29;
  reg        [15:0]   io_in_r_bypass_regNext_12_3_data_29;
  reg                 io_in_r_bypass_regNext_12_3_load_store_29;
  reg                 io_in_r_bypass_regNext_12_3_df_is_ws_29;
  reg                 io_in_r_bypass_regNext_12_3_stall_29;
  reg        [15:0]   io_in_r_bypass_regNext_13_0_data_29;
  reg                 io_in_r_bypass_regNext_13_0_load_store_29;
  reg                 io_in_r_bypass_regNext_13_0_df_is_ws_29;
  reg                 io_in_r_bypass_regNext_13_0_stall_29;
  reg        [15:0]   io_in_r_bypass_regNext_13_1_data_29;
  reg                 io_in_r_bypass_regNext_13_1_load_store_29;
  reg                 io_in_r_bypass_regNext_13_1_df_is_ws_29;
  reg                 io_in_r_bypass_regNext_13_1_stall_29;
  reg        [15:0]   io_in_r_bypass_regNext_13_2_data_29;
  reg                 io_in_r_bypass_regNext_13_2_load_store_29;
  reg                 io_in_r_bypass_regNext_13_2_df_is_ws_29;
  reg                 io_in_r_bypass_regNext_13_2_stall_29;
  reg        [15:0]   io_in_r_bypass_regNext_13_3_data_29;
  reg                 io_in_r_bypass_regNext_13_3_load_store_29;
  reg                 io_in_r_bypass_regNext_13_3_df_is_ws_29;
  reg                 io_in_r_bypass_regNext_13_3_stall_29;
  reg        [15:0]   io_in_r_bypass_regNext_14_0_data_29;
  reg                 io_in_r_bypass_regNext_14_0_load_store_29;
  reg                 io_in_r_bypass_regNext_14_0_df_is_ws_29;
  reg                 io_in_r_bypass_regNext_14_0_stall_29;
  reg        [15:0]   io_in_r_bypass_regNext_14_1_data_29;
  reg                 io_in_r_bypass_regNext_14_1_load_store_29;
  reg                 io_in_r_bypass_regNext_14_1_df_is_ws_29;
  reg                 io_in_r_bypass_regNext_14_1_stall_29;
  reg        [15:0]   io_in_r_bypass_regNext_14_2_data_29;
  reg                 io_in_r_bypass_regNext_14_2_load_store_29;
  reg                 io_in_r_bypass_regNext_14_2_df_is_ws_29;
  reg                 io_in_r_bypass_regNext_14_2_stall_29;
  reg        [15:0]   io_in_r_bypass_regNext_14_3_data_29;
  reg                 io_in_r_bypass_regNext_14_3_load_store_29;
  reg                 io_in_r_bypass_regNext_14_3_df_is_ws_29;
  reg                 io_in_r_bypass_regNext_14_3_stall_29;
  reg        [15:0]   io_in_r_bypass_regNext_15_0_data_29;
  reg                 io_in_r_bypass_regNext_15_0_load_store_29;
  reg                 io_in_r_bypass_regNext_15_0_df_is_ws_29;
  reg                 io_in_r_bypass_regNext_15_0_stall_29;
  reg        [15:0]   io_in_r_bypass_regNext_15_1_data_29;
  reg                 io_in_r_bypass_regNext_15_1_load_store_29;
  reg                 io_in_r_bypass_regNext_15_1_df_is_ws_29;
  reg                 io_in_r_bypass_regNext_15_1_stall_29;
  reg        [15:0]   io_in_r_bypass_regNext_15_2_data_29;
  reg                 io_in_r_bypass_regNext_15_2_load_store_29;
  reg                 io_in_r_bypass_regNext_15_2_df_is_ws_29;
  reg                 io_in_r_bypass_regNext_15_2_stall_29;
  reg        [15:0]   io_in_r_bypass_regNext_15_3_data_29;
  reg                 io_in_r_bypass_regNext_15_3_load_store_29;
  reg                 io_in_r_bypass_regNext_15_3_df_is_ws_29;
  reg                 io_in_r_bypass_regNext_15_3_stall_29;
  reg        [15:0]   io_in_r_bypass_regNext_16_0_data_29;
  reg                 io_in_r_bypass_regNext_16_0_load_store_29;
  reg                 io_in_r_bypass_regNext_16_0_df_is_ws_29;
  reg                 io_in_r_bypass_regNext_16_0_stall_29;
  reg        [15:0]   io_in_r_bypass_regNext_16_1_data_29;
  reg                 io_in_r_bypass_regNext_16_1_load_store_29;
  reg                 io_in_r_bypass_regNext_16_1_df_is_ws_29;
  reg                 io_in_r_bypass_regNext_16_1_stall_29;
  reg        [15:0]   io_in_r_bypass_regNext_16_2_data_29;
  reg                 io_in_r_bypass_regNext_16_2_load_store_29;
  reg                 io_in_r_bypass_regNext_16_2_df_is_ws_29;
  reg                 io_in_r_bypass_regNext_16_2_stall_29;
  reg        [15:0]   io_in_r_bypass_regNext_16_3_data_29;
  reg                 io_in_r_bypass_regNext_16_3_load_store_29;
  reg                 io_in_r_bypass_regNext_16_3_df_is_ws_29;
  reg                 io_in_r_bypass_regNext_16_3_stall_29;
  reg        [15:0]   io_in_r_bypass_regNext_17_0_data_29;
  reg                 io_in_r_bypass_regNext_17_0_load_store_29;
  reg                 io_in_r_bypass_regNext_17_0_df_is_ws_29;
  reg                 io_in_r_bypass_regNext_17_0_stall_29;
  reg        [15:0]   io_in_r_bypass_regNext_17_1_data_29;
  reg                 io_in_r_bypass_regNext_17_1_load_store_29;
  reg                 io_in_r_bypass_regNext_17_1_df_is_ws_29;
  reg                 io_in_r_bypass_regNext_17_1_stall_29;
  reg        [15:0]   io_in_r_bypass_regNext_17_2_data_29;
  reg                 io_in_r_bypass_regNext_17_2_load_store_29;
  reg                 io_in_r_bypass_regNext_17_2_df_is_ws_29;
  reg                 io_in_r_bypass_regNext_17_2_stall_29;
  reg        [15:0]   io_in_r_bypass_regNext_17_3_data_29;
  reg                 io_in_r_bypass_regNext_17_3_load_store_29;
  reg                 io_in_r_bypass_regNext_17_3_df_is_ws_29;
  reg                 io_in_r_bypass_regNext_17_3_stall_29;
  reg        [15:0]   io_in_r_bypass_regNext_18_0_data_29;
  reg                 io_in_r_bypass_regNext_18_0_load_store_29;
  reg                 io_in_r_bypass_regNext_18_0_df_is_ws_29;
  reg                 io_in_r_bypass_regNext_18_0_stall_29;
  reg        [15:0]   io_in_r_bypass_regNext_18_1_data_29;
  reg                 io_in_r_bypass_regNext_18_1_load_store_29;
  reg                 io_in_r_bypass_regNext_18_1_df_is_ws_29;
  reg                 io_in_r_bypass_regNext_18_1_stall_29;
  reg        [15:0]   io_in_r_bypass_regNext_18_2_data_29;
  reg                 io_in_r_bypass_regNext_18_2_load_store_29;
  reg                 io_in_r_bypass_regNext_18_2_df_is_ws_29;
  reg                 io_in_r_bypass_regNext_18_2_stall_29;
  reg        [15:0]   io_in_r_bypass_regNext_18_3_data_29;
  reg                 io_in_r_bypass_regNext_18_3_load_store_29;
  reg                 io_in_r_bypass_regNext_18_3_df_is_ws_29;
  reg                 io_in_r_bypass_regNext_18_3_stall_29;
  reg        [15:0]   io_in_r_bypass_regNext_19_0_data_29;
  reg                 io_in_r_bypass_regNext_19_0_load_store_29;
  reg                 io_in_r_bypass_regNext_19_0_df_is_ws_29;
  reg                 io_in_r_bypass_regNext_19_0_stall_29;
  reg        [15:0]   io_in_r_bypass_regNext_19_1_data_29;
  reg                 io_in_r_bypass_regNext_19_1_load_store_29;
  reg                 io_in_r_bypass_regNext_19_1_df_is_ws_29;
  reg                 io_in_r_bypass_regNext_19_1_stall_29;
  reg        [15:0]   io_in_r_bypass_regNext_19_2_data_29;
  reg                 io_in_r_bypass_regNext_19_2_load_store_29;
  reg                 io_in_r_bypass_regNext_19_2_df_is_ws_29;
  reg                 io_in_r_bypass_regNext_19_2_stall_29;
  reg        [15:0]   io_in_r_bypass_regNext_19_3_data_29;
  reg                 io_in_r_bypass_regNext_19_3_load_store_29;
  reg                 io_in_r_bypass_regNext_19_3_df_is_ws_29;
  reg                 io_in_r_bypass_regNext_19_3_stall_29;
  reg        [15:0]   io_in_r_bypass_regNext_20_0_data_29;
  reg                 io_in_r_bypass_regNext_20_0_load_store_29;
  reg                 io_in_r_bypass_regNext_20_0_df_is_ws_29;
  reg                 io_in_r_bypass_regNext_20_0_stall_29;
  reg        [15:0]   io_in_r_bypass_regNext_20_1_data_29;
  reg                 io_in_r_bypass_regNext_20_1_load_store_29;
  reg                 io_in_r_bypass_regNext_20_1_df_is_ws_29;
  reg                 io_in_r_bypass_regNext_20_1_stall_29;
  reg        [15:0]   io_in_r_bypass_regNext_20_2_data_29;
  reg                 io_in_r_bypass_regNext_20_2_load_store_29;
  reg                 io_in_r_bypass_regNext_20_2_df_is_ws_29;
  reg                 io_in_r_bypass_regNext_20_2_stall_29;
  reg        [15:0]   io_in_r_bypass_regNext_20_3_data_29;
  reg                 io_in_r_bypass_regNext_20_3_load_store_29;
  reg                 io_in_r_bypass_regNext_20_3_df_is_ws_29;
  reg                 io_in_r_bypass_regNext_20_3_stall_29;
  reg        [15:0]   io_in_r_bypass_regNext_21_0_data_29;
  reg                 io_in_r_bypass_regNext_21_0_load_store_29;
  reg                 io_in_r_bypass_regNext_21_0_df_is_ws_29;
  reg                 io_in_r_bypass_regNext_21_0_stall_29;
  reg        [15:0]   io_in_r_bypass_regNext_21_1_data_29;
  reg                 io_in_r_bypass_regNext_21_1_load_store_29;
  reg                 io_in_r_bypass_regNext_21_1_df_is_ws_29;
  reg                 io_in_r_bypass_regNext_21_1_stall_29;
  reg        [15:0]   io_in_r_bypass_regNext_21_2_data_29;
  reg                 io_in_r_bypass_regNext_21_2_load_store_29;
  reg                 io_in_r_bypass_regNext_21_2_df_is_ws_29;
  reg                 io_in_r_bypass_regNext_21_2_stall_29;
  reg        [15:0]   io_in_r_bypass_regNext_21_3_data_29;
  reg                 io_in_r_bypass_regNext_21_3_load_store_29;
  reg                 io_in_r_bypass_regNext_21_3_df_is_ws_29;
  reg                 io_in_r_bypass_regNext_21_3_stall_29;
  reg        [15:0]   io_in_r_bypass_regNext_22_0_data_29;
  reg                 io_in_r_bypass_regNext_22_0_load_store_29;
  reg                 io_in_r_bypass_regNext_22_0_df_is_ws_29;
  reg                 io_in_r_bypass_regNext_22_0_stall_29;
  reg        [15:0]   io_in_r_bypass_regNext_22_1_data_29;
  reg                 io_in_r_bypass_regNext_22_1_load_store_29;
  reg                 io_in_r_bypass_regNext_22_1_df_is_ws_29;
  reg                 io_in_r_bypass_regNext_22_1_stall_29;
  reg        [15:0]   io_in_r_bypass_regNext_22_2_data_29;
  reg                 io_in_r_bypass_regNext_22_2_load_store_29;
  reg                 io_in_r_bypass_regNext_22_2_df_is_ws_29;
  reg                 io_in_r_bypass_regNext_22_2_stall_29;
  reg        [15:0]   io_in_r_bypass_regNext_22_3_data_29;
  reg                 io_in_r_bypass_regNext_22_3_load_store_29;
  reg                 io_in_r_bypass_regNext_22_3_df_is_ws_29;
  reg                 io_in_r_bypass_regNext_22_3_stall_29;
  reg        [15:0]   io_in_r_bypass_regNext_23_0_data_29;
  reg                 io_in_r_bypass_regNext_23_0_load_store_29;
  reg                 io_in_r_bypass_regNext_23_0_df_is_ws_29;
  reg                 io_in_r_bypass_regNext_23_0_stall_29;
  reg        [15:0]   io_in_r_bypass_regNext_23_1_data_29;
  reg                 io_in_r_bypass_regNext_23_1_load_store_29;
  reg                 io_in_r_bypass_regNext_23_1_df_is_ws_29;
  reg                 io_in_r_bypass_regNext_23_1_stall_29;
  reg        [15:0]   io_in_r_bypass_regNext_23_2_data_29;
  reg                 io_in_r_bypass_regNext_23_2_load_store_29;
  reg                 io_in_r_bypass_regNext_23_2_df_is_ws_29;
  reg                 io_in_r_bypass_regNext_23_2_stall_29;
  reg        [15:0]   io_in_r_bypass_regNext_23_3_data_29;
  reg                 io_in_r_bypass_regNext_23_3_load_store_29;
  reg                 io_in_r_bypass_regNext_23_3_df_is_ws_29;
  reg                 io_in_r_bypass_regNext_23_3_stall_29;
  reg        [15:0]   io_in_r_bypass_regNext_24_0_data_29;
  reg                 io_in_r_bypass_regNext_24_0_load_store_29;
  reg                 io_in_r_bypass_regNext_24_0_df_is_ws_29;
  reg                 io_in_r_bypass_regNext_24_0_stall_29;
  reg        [15:0]   io_in_r_bypass_regNext_24_1_data_29;
  reg                 io_in_r_bypass_regNext_24_1_load_store_29;
  reg                 io_in_r_bypass_regNext_24_1_df_is_ws_29;
  reg                 io_in_r_bypass_regNext_24_1_stall_29;
  reg        [15:0]   io_in_r_bypass_regNext_24_2_data_29;
  reg                 io_in_r_bypass_regNext_24_2_load_store_29;
  reg                 io_in_r_bypass_regNext_24_2_df_is_ws_29;
  reg                 io_in_r_bypass_regNext_24_2_stall_29;
  reg        [15:0]   io_in_r_bypass_regNext_24_3_data_29;
  reg                 io_in_r_bypass_regNext_24_3_load_store_29;
  reg                 io_in_r_bypass_regNext_24_3_df_is_ws_29;
  reg                 io_in_r_bypass_regNext_24_3_stall_29;
  reg        [15:0]   io_in_r_bypass_regNext_25_0_data_29;
  reg                 io_in_r_bypass_regNext_25_0_load_store_29;
  reg                 io_in_r_bypass_regNext_25_0_df_is_ws_29;
  reg                 io_in_r_bypass_regNext_25_0_stall_29;
  reg        [15:0]   io_in_r_bypass_regNext_25_1_data_29;
  reg                 io_in_r_bypass_regNext_25_1_load_store_29;
  reg                 io_in_r_bypass_regNext_25_1_df_is_ws_29;
  reg                 io_in_r_bypass_regNext_25_1_stall_29;
  reg        [15:0]   io_in_r_bypass_regNext_25_2_data_29;
  reg                 io_in_r_bypass_regNext_25_2_load_store_29;
  reg                 io_in_r_bypass_regNext_25_2_df_is_ws_29;
  reg                 io_in_r_bypass_regNext_25_2_stall_29;
  reg        [15:0]   io_in_r_bypass_regNext_25_3_data_29;
  reg                 io_in_r_bypass_regNext_25_3_load_store_29;
  reg                 io_in_r_bypass_regNext_25_3_df_is_ws_29;
  reg                 io_in_r_bypass_regNext_25_3_stall_29;
  reg        [15:0]   io_in_r_bypass_regNext_26_0_data_29;
  reg                 io_in_r_bypass_regNext_26_0_load_store_29;
  reg                 io_in_r_bypass_regNext_26_0_df_is_ws_29;
  reg                 io_in_r_bypass_regNext_26_0_stall_29;
  reg        [15:0]   io_in_r_bypass_regNext_26_1_data_29;
  reg                 io_in_r_bypass_regNext_26_1_load_store_29;
  reg                 io_in_r_bypass_regNext_26_1_df_is_ws_29;
  reg                 io_in_r_bypass_regNext_26_1_stall_29;
  reg        [15:0]   io_in_r_bypass_regNext_26_2_data_29;
  reg                 io_in_r_bypass_regNext_26_2_load_store_29;
  reg                 io_in_r_bypass_regNext_26_2_df_is_ws_29;
  reg                 io_in_r_bypass_regNext_26_2_stall_29;
  reg        [15:0]   io_in_r_bypass_regNext_26_3_data_29;
  reg                 io_in_r_bypass_regNext_26_3_load_store_29;
  reg                 io_in_r_bypass_regNext_26_3_df_is_ws_29;
  reg                 io_in_r_bypass_regNext_26_3_stall_29;
  reg        [15:0]   io_in_r_bypass_regNext_27_0_data_29;
  reg                 io_in_r_bypass_regNext_27_0_load_store_29;
  reg                 io_in_r_bypass_regNext_27_0_df_is_ws_29;
  reg                 io_in_r_bypass_regNext_27_0_stall_29;
  reg        [15:0]   io_in_r_bypass_regNext_27_1_data_29;
  reg                 io_in_r_bypass_regNext_27_1_load_store_29;
  reg                 io_in_r_bypass_regNext_27_1_df_is_ws_29;
  reg                 io_in_r_bypass_regNext_27_1_stall_29;
  reg        [15:0]   io_in_r_bypass_regNext_27_2_data_29;
  reg                 io_in_r_bypass_regNext_27_2_load_store_29;
  reg                 io_in_r_bypass_regNext_27_2_df_is_ws_29;
  reg                 io_in_r_bypass_regNext_27_2_stall_29;
  reg        [15:0]   io_in_r_bypass_regNext_27_3_data_29;
  reg                 io_in_r_bypass_regNext_27_3_load_store_29;
  reg                 io_in_r_bypass_regNext_27_3_df_is_ws_29;
  reg                 io_in_r_bypass_regNext_27_3_stall_29;
  reg        [15:0]   io_in_r_bypass_regNext_28_0_data_29;
  reg                 io_in_r_bypass_regNext_28_0_load_store_29;
  reg                 io_in_r_bypass_regNext_28_0_df_is_ws_29;
  reg                 io_in_r_bypass_regNext_28_0_stall_29;
  reg        [15:0]   io_in_r_bypass_regNext_28_1_data_29;
  reg                 io_in_r_bypass_regNext_28_1_load_store_29;
  reg                 io_in_r_bypass_regNext_28_1_df_is_ws_29;
  reg                 io_in_r_bypass_regNext_28_1_stall_29;
  reg        [15:0]   io_in_r_bypass_regNext_28_2_data_29;
  reg                 io_in_r_bypass_regNext_28_2_load_store_29;
  reg                 io_in_r_bypass_regNext_28_2_df_is_ws_29;
  reg                 io_in_r_bypass_regNext_28_2_stall_29;
  reg        [15:0]   io_in_r_bypass_regNext_28_3_data_29;
  reg                 io_in_r_bypass_regNext_28_3_load_store_29;
  reg                 io_in_r_bypass_regNext_28_3_df_is_ws_29;
  reg                 io_in_r_bypass_regNext_28_3_stall_29;
  reg        [15:0]   io_in_r_bypass_regNext_29_0_data_29;
  reg                 io_in_r_bypass_regNext_29_0_load_store_29;
  reg                 io_in_r_bypass_regNext_29_0_df_is_ws_29;
  reg                 io_in_r_bypass_regNext_29_0_stall_29;
  reg        [15:0]   io_in_r_bypass_regNext_29_1_data_29;
  reg                 io_in_r_bypass_regNext_29_1_load_store_29;
  reg                 io_in_r_bypass_regNext_29_1_df_is_ws_29;
  reg                 io_in_r_bypass_regNext_29_1_stall_29;
  reg        [15:0]   io_in_r_bypass_regNext_29_2_data_29;
  reg                 io_in_r_bypass_regNext_29_2_load_store_29;
  reg                 io_in_r_bypass_regNext_29_2_df_is_ws_29;
  reg                 io_in_r_bypass_regNext_29_2_stall_29;
  reg        [15:0]   io_in_r_bypass_regNext_29_3_data_29;
  reg                 io_in_r_bypass_regNext_29_3_load_store_29;
  reg                 io_in_r_bypass_regNext_29_3_df_is_ws_29;
  reg                 io_in_r_bypass_regNext_29_3_stall_29;
  reg        [15:0]   io_in_r_bypass_regNext_30_0_data_29;
  reg                 io_in_r_bypass_regNext_30_0_load_store_29;
  reg                 io_in_r_bypass_regNext_30_0_df_is_ws_29;
  reg                 io_in_r_bypass_regNext_30_0_stall_29;
  reg        [15:0]   io_in_r_bypass_regNext_30_1_data_29;
  reg                 io_in_r_bypass_regNext_30_1_load_store_29;
  reg                 io_in_r_bypass_regNext_30_1_df_is_ws_29;
  reg                 io_in_r_bypass_regNext_30_1_stall_29;
  reg        [15:0]   io_in_r_bypass_regNext_30_2_data_29;
  reg                 io_in_r_bypass_regNext_30_2_load_store_29;
  reg                 io_in_r_bypass_regNext_30_2_df_is_ws_29;
  reg                 io_in_r_bypass_regNext_30_2_stall_29;
  reg        [15:0]   io_in_r_bypass_regNext_30_3_data_29;
  reg                 io_in_r_bypass_regNext_30_3_load_store_29;
  reg                 io_in_r_bypass_regNext_30_3_df_is_ws_29;
  reg                 io_in_r_bypass_regNext_30_3_stall_29;
  reg        [15:0]   io_in_r_bypass_regNext_31_0_data_29;
  reg                 io_in_r_bypass_regNext_31_0_load_store_29;
  reg                 io_in_r_bypass_regNext_31_0_df_is_ws_29;
  reg                 io_in_r_bypass_regNext_31_0_stall_29;
  reg        [15:0]   io_in_r_bypass_regNext_31_1_data_29;
  reg                 io_in_r_bypass_regNext_31_1_load_store_29;
  reg                 io_in_r_bypass_regNext_31_1_df_is_ws_29;
  reg                 io_in_r_bypass_regNext_31_1_stall_29;
  reg        [15:0]   io_in_r_bypass_regNext_31_2_data_29;
  reg                 io_in_r_bypass_regNext_31_2_load_store_29;
  reg                 io_in_r_bypass_regNext_31_2_df_is_ws_29;
  reg                 io_in_r_bypass_regNext_31_2_stall_29;
  reg        [15:0]   io_in_r_bypass_regNext_31_3_data_29;
  reg                 io_in_r_bypass_regNext_31_3_load_store_29;
  reg                 io_in_r_bypass_regNext_31_3_df_is_ws_29;
  reg                 io_in_r_bypass_regNext_31_3_stall_29;
  reg        [15:0]   io_in_r_bypass_regNext_0_0_data_30;
  reg                 io_in_r_bypass_regNext_0_0_load_store_30;
  reg                 io_in_r_bypass_regNext_0_0_df_is_ws_30;
  reg                 io_in_r_bypass_regNext_0_0_stall_30;
  reg        [15:0]   io_in_r_bypass_regNext_0_1_data_30;
  reg                 io_in_r_bypass_regNext_0_1_load_store_30;
  reg                 io_in_r_bypass_regNext_0_1_df_is_ws_30;
  reg                 io_in_r_bypass_regNext_0_1_stall_30;
  reg        [15:0]   io_in_r_bypass_regNext_0_2_data_30;
  reg                 io_in_r_bypass_regNext_0_2_load_store_30;
  reg                 io_in_r_bypass_regNext_0_2_df_is_ws_30;
  reg                 io_in_r_bypass_regNext_0_2_stall_30;
  reg        [15:0]   io_in_r_bypass_regNext_0_3_data_30;
  reg                 io_in_r_bypass_regNext_0_3_load_store_30;
  reg                 io_in_r_bypass_regNext_0_3_df_is_ws_30;
  reg                 io_in_r_bypass_regNext_0_3_stall_30;
  reg        [15:0]   io_in_r_bypass_regNext_1_0_data_30;
  reg                 io_in_r_bypass_regNext_1_0_load_store_30;
  reg                 io_in_r_bypass_regNext_1_0_df_is_ws_30;
  reg                 io_in_r_bypass_regNext_1_0_stall_30;
  reg        [15:0]   io_in_r_bypass_regNext_1_1_data_30;
  reg                 io_in_r_bypass_regNext_1_1_load_store_30;
  reg                 io_in_r_bypass_regNext_1_1_df_is_ws_30;
  reg                 io_in_r_bypass_regNext_1_1_stall_30;
  reg        [15:0]   io_in_r_bypass_regNext_1_2_data_30;
  reg                 io_in_r_bypass_regNext_1_2_load_store_30;
  reg                 io_in_r_bypass_regNext_1_2_df_is_ws_30;
  reg                 io_in_r_bypass_regNext_1_2_stall_30;
  reg        [15:0]   io_in_r_bypass_regNext_1_3_data_30;
  reg                 io_in_r_bypass_regNext_1_3_load_store_30;
  reg                 io_in_r_bypass_regNext_1_3_df_is_ws_30;
  reg                 io_in_r_bypass_regNext_1_3_stall_30;
  reg        [15:0]   io_in_r_bypass_regNext_2_0_data_30;
  reg                 io_in_r_bypass_regNext_2_0_load_store_30;
  reg                 io_in_r_bypass_regNext_2_0_df_is_ws_30;
  reg                 io_in_r_bypass_regNext_2_0_stall_30;
  reg        [15:0]   io_in_r_bypass_regNext_2_1_data_30;
  reg                 io_in_r_bypass_regNext_2_1_load_store_30;
  reg                 io_in_r_bypass_regNext_2_1_df_is_ws_30;
  reg                 io_in_r_bypass_regNext_2_1_stall_30;
  reg        [15:0]   io_in_r_bypass_regNext_2_2_data_30;
  reg                 io_in_r_bypass_regNext_2_2_load_store_30;
  reg                 io_in_r_bypass_regNext_2_2_df_is_ws_30;
  reg                 io_in_r_bypass_regNext_2_2_stall_30;
  reg        [15:0]   io_in_r_bypass_regNext_2_3_data_30;
  reg                 io_in_r_bypass_regNext_2_3_load_store_30;
  reg                 io_in_r_bypass_regNext_2_3_df_is_ws_30;
  reg                 io_in_r_bypass_regNext_2_3_stall_30;
  reg        [15:0]   io_in_r_bypass_regNext_3_0_data_30;
  reg                 io_in_r_bypass_regNext_3_0_load_store_30;
  reg                 io_in_r_bypass_regNext_3_0_df_is_ws_30;
  reg                 io_in_r_bypass_regNext_3_0_stall_30;
  reg        [15:0]   io_in_r_bypass_regNext_3_1_data_30;
  reg                 io_in_r_bypass_regNext_3_1_load_store_30;
  reg                 io_in_r_bypass_regNext_3_1_df_is_ws_30;
  reg                 io_in_r_bypass_regNext_3_1_stall_30;
  reg        [15:0]   io_in_r_bypass_regNext_3_2_data_30;
  reg                 io_in_r_bypass_regNext_3_2_load_store_30;
  reg                 io_in_r_bypass_regNext_3_2_df_is_ws_30;
  reg                 io_in_r_bypass_regNext_3_2_stall_30;
  reg        [15:0]   io_in_r_bypass_regNext_3_3_data_30;
  reg                 io_in_r_bypass_regNext_3_3_load_store_30;
  reg                 io_in_r_bypass_regNext_3_3_df_is_ws_30;
  reg                 io_in_r_bypass_regNext_3_3_stall_30;
  reg        [15:0]   io_in_r_bypass_regNext_4_0_data_30;
  reg                 io_in_r_bypass_regNext_4_0_load_store_30;
  reg                 io_in_r_bypass_regNext_4_0_df_is_ws_30;
  reg                 io_in_r_bypass_regNext_4_0_stall_30;
  reg        [15:0]   io_in_r_bypass_regNext_4_1_data_30;
  reg                 io_in_r_bypass_regNext_4_1_load_store_30;
  reg                 io_in_r_bypass_regNext_4_1_df_is_ws_30;
  reg                 io_in_r_bypass_regNext_4_1_stall_30;
  reg        [15:0]   io_in_r_bypass_regNext_4_2_data_30;
  reg                 io_in_r_bypass_regNext_4_2_load_store_30;
  reg                 io_in_r_bypass_regNext_4_2_df_is_ws_30;
  reg                 io_in_r_bypass_regNext_4_2_stall_30;
  reg        [15:0]   io_in_r_bypass_regNext_4_3_data_30;
  reg                 io_in_r_bypass_regNext_4_3_load_store_30;
  reg                 io_in_r_bypass_regNext_4_3_df_is_ws_30;
  reg                 io_in_r_bypass_regNext_4_3_stall_30;
  reg        [15:0]   io_in_r_bypass_regNext_5_0_data_30;
  reg                 io_in_r_bypass_regNext_5_0_load_store_30;
  reg                 io_in_r_bypass_regNext_5_0_df_is_ws_30;
  reg                 io_in_r_bypass_regNext_5_0_stall_30;
  reg        [15:0]   io_in_r_bypass_regNext_5_1_data_30;
  reg                 io_in_r_bypass_regNext_5_1_load_store_30;
  reg                 io_in_r_bypass_regNext_5_1_df_is_ws_30;
  reg                 io_in_r_bypass_regNext_5_1_stall_30;
  reg        [15:0]   io_in_r_bypass_regNext_5_2_data_30;
  reg                 io_in_r_bypass_regNext_5_2_load_store_30;
  reg                 io_in_r_bypass_regNext_5_2_df_is_ws_30;
  reg                 io_in_r_bypass_regNext_5_2_stall_30;
  reg        [15:0]   io_in_r_bypass_regNext_5_3_data_30;
  reg                 io_in_r_bypass_regNext_5_3_load_store_30;
  reg                 io_in_r_bypass_regNext_5_3_df_is_ws_30;
  reg                 io_in_r_bypass_regNext_5_3_stall_30;
  reg        [15:0]   io_in_r_bypass_regNext_6_0_data_30;
  reg                 io_in_r_bypass_regNext_6_0_load_store_30;
  reg                 io_in_r_bypass_regNext_6_0_df_is_ws_30;
  reg                 io_in_r_bypass_regNext_6_0_stall_30;
  reg        [15:0]   io_in_r_bypass_regNext_6_1_data_30;
  reg                 io_in_r_bypass_regNext_6_1_load_store_30;
  reg                 io_in_r_bypass_regNext_6_1_df_is_ws_30;
  reg                 io_in_r_bypass_regNext_6_1_stall_30;
  reg        [15:0]   io_in_r_bypass_regNext_6_2_data_30;
  reg                 io_in_r_bypass_regNext_6_2_load_store_30;
  reg                 io_in_r_bypass_regNext_6_2_df_is_ws_30;
  reg                 io_in_r_bypass_regNext_6_2_stall_30;
  reg        [15:0]   io_in_r_bypass_regNext_6_3_data_30;
  reg                 io_in_r_bypass_regNext_6_3_load_store_30;
  reg                 io_in_r_bypass_regNext_6_3_df_is_ws_30;
  reg                 io_in_r_bypass_regNext_6_3_stall_30;
  reg        [15:0]   io_in_r_bypass_regNext_7_0_data_30;
  reg                 io_in_r_bypass_regNext_7_0_load_store_30;
  reg                 io_in_r_bypass_regNext_7_0_df_is_ws_30;
  reg                 io_in_r_bypass_regNext_7_0_stall_30;
  reg        [15:0]   io_in_r_bypass_regNext_7_1_data_30;
  reg                 io_in_r_bypass_regNext_7_1_load_store_30;
  reg                 io_in_r_bypass_regNext_7_1_df_is_ws_30;
  reg                 io_in_r_bypass_regNext_7_1_stall_30;
  reg        [15:0]   io_in_r_bypass_regNext_7_2_data_30;
  reg                 io_in_r_bypass_regNext_7_2_load_store_30;
  reg                 io_in_r_bypass_regNext_7_2_df_is_ws_30;
  reg                 io_in_r_bypass_regNext_7_2_stall_30;
  reg        [15:0]   io_in_r_bypass_regNext_7_3_data_30;
  reg                 io_in_r_bypass_regNext_7_3_load_store_30;
  reg                 io_in_r_bypass_regNext_7_3_df_is_ws_30;
  reg                 io_in_r_bypass_regNext_7_3_stall_30;
  reg        [15:0]   io_in_r_bypass_regNext_8_0_data_30;
  reg                 io_in_r_bypass_regNext_8_0_load_store_30;
  reg                 io_in_r_bypass_regNext_8_0_df_is_ws_30;
  reg                 io_in_r_bypass_regNext_8_0_stall_30;
  reg        [15:0]   io_in_r_bypass_regNext_8_1_data_30;
  reg                 io_in_r_bypass_regNext_8_1_load_store_30;
  reg                 io_in_r_bypass_regNext_8_1_df_is_ws_30;
  reg                 io_in_r_bypass_regNext_8_1_stall_30;
  reg        [15:0]   io_in_r_bypass_regNext_8_2_data_30;
  reg                 io_in_r_bypass_regNext_8_2_load_store_30;
  reg                 io_in_r_bypass_regNext_8_2_df_is_ws_30;
  reg                 io_in_r_bypass_regNext_8_2_stall_30;
  reg        [15:0]   io_in_r_bypass_regNext_8_3_data_30;
  reg                 io_in_r_bypass_regNext_8_3_load_store_30;
  reg                 io_in_r_bypass_regNext_8_3_df_is_ws_30;
  reg                 io_in_r_bypass_regNext_8_3_stall_30;
  reg        [15:0]   io_in_r_bypass_regNext_9_0_data_30;
  reg                 io_in_r_bypass_regNext_9_0_load_store_30;
  reg                 io_in_r_bypass_regNext_9_0_df_is_ws_30;
  reg                 io_in_r_bypass_regNext_9_0_stall_30;
  reg        [15:0]   io_in_r_bypass_regNext_9_1_data_30;
  reg                 io_in_r_bypass_regNext_9_1_load_store_30;
  reg                 io_in_r_bypass_regNext_9_1_df_is_ws_30;
  reg                 io_in_r_bypass_regNext_9_1_stall_30;
  reg        [15:0]   io_in_r_bypass_regNext_9_2_data_30;
  reg                 io_in_r_bypass_regNext_9_2_load_store_30;
  reg                 io_in_r_bypass_regNext_9_2_df_is_ws_30;
  reg                 io_in_r_bypass_regNext_9_2_stall_30;
  reg        [15:0]   io_in_r_bypass_regNext_9_3_data_30;
  reg                 io_in_r_bypass_regNext_9_3_load_store_30;
  reg                 io_in_r_bypass_regNext_9_3_df_is_ws_30;
  reg                 io_in_r_bypass_regNext_9_3_stall_30;
  reg        [15:0]   io_in_r_bypass_regNext_10_0_data_30;
  reg                 io_in_r_bypass_regNext_10_0_load_store_30;
  reg                 io_in_r_bypass_regNext_10_0_df_is_ws_30;
  reg                 io_in_r_bypass_regNext_10_0_stall_30;
  reg        [15:0]   io_in_r_bypass_regNext_10_1_data_30;
  reg                 io_in_r_bypass_regNext_10_1_load_store_30;
  reg                 io_in_r_bypass_regNext_10_1_df_is_ws_30;
  reg                 io_in_r_bypass_regNext_10_1_stall_30;
  reg        [15:0]   io_in_r_bypass_regNext_10_2_data_30;
  reg                 io_in_r_bypass_regNext_10_2_load_store_30;
  reg                 io_in_r_bypass_regNext_10_2_df_is_ws_30;
  reg                 io_in_r_bypass_regNext_10_2_stall_30;
  reg        [15:0]   io_in_r_bypass_regNext_10_3_data_30;
  reg                 io_in_r_bypass_regNext_10_3_load_store_30;
  reg                 io_in_r_bypass_regNext_10_3_df_is_ws_30;
  reg                 io_in_r_bypass_regNext_10_3_stall_30;
  reg        [15:0]   io_in_r_bypass_regNext_11_0_data_30;
  reg                 io_in_r_bypass_regNext_11_0_load_store_30;
  reg                 io_in_r_bypass_regNext_11_0_df_is_ws_30;
  reg                 io_in_r_bypass_regNext_11_0_stall_30;
  reg        [15:0]   io_in_r_bypass_regNext_11_1_data_30;
  reg                 io_in_r_bypass_regNext_11_1_load_store_30;
  reg                 io_in_r_bypass_regNext_11_1_df_is_ws_30;
  reg                 io_in_r_bypass_regNext_11_1_stall_30;
  reg        [15:0]   io_in_r_bypass_regNext_11_2_data_30;
  reg                 io_in_r_bypass_regNext_11_2_load_store_30;
  reg                 io_in_r_bypass_regNext_11_2_df_is_ws_30;
  reg                 io_in_r_bypass_regNext_11_2_stall_30;
  reg        [15:0]   io_in_r_bypass_regNext_11_3_data_30;
  reg                 io_in_r_bypass_regNext_11_3_load_store_30;
  reg                 io_in_r_bypass_regNext_11_3_df_is_ws_30;
  reg                 io_in_r_bypass_regNext_11_3_stall_30;
  reg        [15:0]   io_in_r_bypass_regNext_12_0_data_30;
  reg                 io_in_r_bypass_regNext_12_0_load_store_30;
  reg                 io_in_r_bypass_regNext_12_0_df_is_ws_30;
  reg                 io_in_r_bypass_regNext_12_0_stall_30;
  reg        [15:0]   io_in_r_bypass_regNext_12_1_data_30;
  reg                 io_in_r_bypass_regNext_12_1_load_store_30;
  reg                 io_in_r_bypass_regNext_12_1_df_is_ws_30;
  reg                 io_in_r_bypass_regNext_12_1_stall_30;
  reg        [15:0]   io_in_r_bypass_regNext_12_2_data_30;
  reg                 io_in_r_bypass_regNext_12_2_load_store_30;
  reg                 io_in_r_bypass_regNext_12_2_df_is_ws_30;
  reg                 io_in_r_bypass_regNext_12_2_stall_30;
  reg        [15:0]   io_in_r_bypass_regNext_12_3_data_30;
  reg                 io_in_r_bypass_regNext_12_3_load_store_30;
  reg                 io_in_r_bypass_regNext_12_3_df_is_ws_30;
  reg                 io_in_r_bypass_regNext_12_3_stall_30;
  reg        [15:0]   io_in_r_bypass_regNext_13_0_data_30;
  reg                 io_in_r_bypass_regNext_13_0_load_store_30;
  reg                 io_in_r_bypass_regNext_13_0_df_is_ws_30;
  reg                 io_in_r_bypass_regNext_13_0_stall_30;
  reg        [15:0]   io_in_r_bypass_regNext_13_1_data_30;
  reg                 io_in_r_bypass_regNext_13_1_load_store_30;
  reg                 io_in_r_bypass_regNext_13_1_df_is_ws_30;
  reg                 io_in_r_bypass_regNext_13_1_stall_30;
  reg        [15:0]   io_in_r_bypass_regNext_13_2_data_30;
  reg                 io_in_r_bypass_regNext_13_2_load_store_30;
  reg                 io_in_r_bypass_regNext_13_2_df_is_ws_30;
  reg                 io_in_r_bypass_regNext_13_2_stall_30;
  reg        [15:0]   io_in_r_bypass_regNext_13_3_data_30;
  reg                 io_in_r_bypass_regNext_13_3_load_store_30;
  reg                 io_in_r_bypass_regNext_13_3_df_is_ws_30;
  reg                 io_in_r_bypass_regNext_13_3_stall_30;
  reg        [15:0]   io_in_r_bypass_regNext_14_0_data_30;
  reg                 io_in_r_bypass_regNext_14_0_load_store_30;
  reg                 io_in_r_bypass_regNext_14_0_df_is_ws_30;
  reg                 io_in_r_bypass_regNext_14_0_stall_30;
  reg        [15:0]   io_in_r_bypass_regNext_14_1_data_30;
  reg                 io_in_r_bypass_regNext_14_1_load_store_30;
  reg                 io_in_r_bypass_regNext_14_1_df_is_ws_30;
  reg                 io_in_r_bypass_regNext_14_1_stall_30;
  reg        [15:0]   io_in_r_bypass_regNext_14_2_data_30;
  reg                 io_in_r_bypass_regNext_14_2_load_store_30;
  reg                 io_in_r_bypass_regNext_14_2_df_is_ws_30;
  reg                 io_in_r_bypass_regNext_14_2_stall_30;
  reg        [15:0]   io_in_r_bypass_regNext_14_3_data_30;
  reg                 io_in_r_bypass_regNext_14_3_load_store_30;
  reg                 io_in_r_bypass_regNext_14_3_df_is_ws_30;
  reg                 io_in_r_bypass_regNext_14_3_stall_30;
  reg        [15:0]   io_in_r_bypass_regNext_15_0_data_30;
  reg                 io_in_r_bypass_regNext_15_0_load_store_30;
  reg                 io_in_r_bypass_regNext_15_0_df_is_ws_30;
  reg                 io_in_r_bypass_regNext_15_0_stall_30;
  reg        [15:0]   io_in_r_bypass_regNext_15_1_data_30;
  reg                 io_in_r_bypass_regNext_15_1_load_store_30;
  reg                 io_in_r_bypass_regNext_15_1_df_is_ws_30;
  reg                 io_in_r_bypass_regNext_15_1_stall_30;
  reg        [15:0]   io_in_r_bypass_regNext_15_2_data_30;
  reg                 io_in_r_bypass_regNext_15_2_load_store_30;
  reg                 io_in_r_bypass_regNext_15_2_df_is_ws_30;
  reg                 io_in_r_bypass_regNext_15_2_stall_30;
  reg        [15:0]   io_in_r_bypass_regNext_15_3_data_30;
  reg                 io_in_r_bypass_regNext_15_3_load_store_30;
  reg                 io_in_r_bypass_regNext_15_3_df_is_ws_30;
  reg                 io_in_r_bypass_regNext_15_3_stall_30;
  reg        [15:0]   io_in_r_bypass_regNext_16_0_data_30;
  reg                 io_in_r_bypass_regNext_16_0_load_store_30;
  reg                 io_in_r_bypass_regNext_16_0_df_is_ws_30;
  reg                 io_in_r_bypass_regNext_16_0_stall_30;
  reg        [15:0]   io_in_r_bypass_regNext_16_1_data_30;
  reg                 io_in_r_bypass_regNext_16_1_load_store_30;
  reg                 io_in_r_bypass_regNext_16_1_df_is_ws_30;
  reg                 io_in_r_bypass_regNext_16_1_stall_30;
  reg        [15:0]   io_in_r_bypass_regNext_16_2_data_30;
  reg                 io_in_r_bypass_regNext_16_2_load_store_30;
  reg                 io_in_r_bypass_regNext_16_2_df_is_ws_30;
  reg                 io_in_r_bypass_regNext_16_2_stall_30;
  reg        [15:0]   io_in_r_bypass_regNext_16_3_data_30;
  reg                 io_in_r_bypass_regNext_16_3_load_store_30;
  reg                 io_in_r_bypass_regNext_16_3_df_is_ws_30;
  reg                 io_in_r_bypass_regNext_16_3_stall_30;
  reg        [15:0]   io_in_r_bypass_regNext_17_0_data_30;
  reg                 io_in_r_bypass_regNext_17_0_load_store_30;
  reg                 io_in_r_bypass_regNext_17_0_df_is_ws_30;
  reg                 io_in_r_bypass_regNext_17_0_stall_30;
  reg        [15:0]   io_in_r_bypass_regNext_17_1_data_30;
  reg                 io_in_r_bypass_regNext_17_1_load_store_30;
  reg                 io_in_r_bypass_regNext_17_1_df_is_ws_30;
  reg                 io_in_r_bypass_regNext_17_1_stall_30;
  reg        [15:0]   io_in_r_bypass_regNext_17_2_data_30;
  reg                 io_in_r_bypass_regNext_17_2_load_store_30;
  reg                 io_in_r_bypass_regNext_17_2_df_is_ws_30;
  reg                 io_in_r_bypass_regNext_17_2_stall_30;
  reg        [15:0]   io_in_r_bypass_regNext_17_3_data_30;
  reg                 io_in_r_bypass_regNext_17_3_load_store_30;
  reg                 io_in_r_bypass_regNext_17_3_df_is_ws_30;
  reg                 io_in_r_bypass_regNext_17_3_stall_30;
  reg        [15:0]   io_in_r_bypass_regNext_18_0_data_30;
  reg                 io_in_r_bypass_regNext_18_0_load_store_30;
  reg                 io_in_r_bypass_regNext_18_0_df_is_ws_30;
  reg                 io_in_r_bypass_regNext_18_0_stall_30;
  reg        [15:0]   io_in_r_bypass_regNext_18_1_data_30;
  reg                 io_in_r_bypass_regNext_18_1_load_store_30;
  reg                 io_in_r_bypass_regNext_18_1_df_is_ws_30;
  reg                 io_in_r_bypass_regNext_18_1_stall_30;
  reg        [15:0]   io_in_r_bypass_regNext_18_2_data_30;
  reg                 io_in_r_bypass_regNext_18_2_load_store_30;
  reg                 io_in_r_bypass_regNext_18_2_df_is_ws_30;
  reg                 io_in_r_bypass_regNext_18_2_stall_30;
  reg        [15:0]   io_in_r_bypass_regNext_18_3_data_30;
  reg                 io_in_r_bypass_regNext_18_3_load_store_30;
  reg                 io_in_r_bypass_regNext_18_3_df_is_ws_30;
  reg                 io_in_r_bypass_regNext_18_3_stall_30;
  reg        [15:0]   io_in_r_bypass_regNext_19_0_data_30;
  reg                 io_in_r_bypass_regNext_19_0_load_store_30;
  reg                 io_in_r_bypass_regNext_19_0_df_is_ws_30;
  reg                 io_in_r_bypass_regNext_19_0_stall_30;
  reg        [15:0]   io_in_r_bypass_regNext_19_1_data_30;
  reg                 io_in_r_bypass_regNext_19_1_load_store_30;
  reg                 io_in_r_bypass_regNext_19_1_df_is_ws_30;
  reg                 io_in_r_bypass_regNext_19_1_stall_30;
  reg        [15:0]   io_in_r_bypass_regNext_19_2_data_30;
  reg                 io_in_r_bypass_regNext_19_2_load_store_30;
  reg                 io_in_r_bypass_regNext_19_2_df_is_ws_30;
  reg                 io_in_r_bypass_regNext_19_2_stall_30;
  reg        [15:0]   io_in_r_bypass_regNext_19_3_data_30;
  reg                 io_in_r_bypass_regNext_19_3_load_store_30;
  reg                 io_in_r_bypass_regNext_19_3_df_is_ws_30;
  reg                 io_in_r_bypass_regNext_19_3_stall_30;
  reg        [15:0]   io_in_r_bypass_regNext_20_0_data_30;
  reg                 io_in_r_bypass_regNext_20_0_load_store_30;
  reg                 io_in_r_bypass_regNext_20_0_df_is_ws_30;
  reg                 io_in_r_bypass_regNext_20_0_stall_30;
  reg        [15:0]   io_in_r_bypass_regNext_20_1_data_30;
  reg                 io_in_r_bypass_regNext_20_1_load_store_30;
  reg                 io_in_r_bypass_regNext_20_1_df_is_ws_30;
  reg                 io_in_r_bypass_regNext_20_1_stall_30;
  reg        [15:0]   io_in_r_bypass_regNext_20_2_data_30;
  reg                 io_in_r_bypass_regNext_20_2_load_store_30;
  reg                 io_in_r_bypass_regNext_20_2_df_is_ws_30;
  reg                 io_in_r_bypass_regNext_20_2_stall_30;
  reg        [15:0]   io_in_r_bypass_regNext_20_3_data_30;
  reg                 io_in_r_bypass_regNext_20_3_load_store_30;
  reg                 io_in_r_bypass_regNext_20_3_df_is_ws_30;
  reg                 io_in_r_bypass_regNext_20_3_stall_30;
  reg        [15:0]   io_in_r_bypass_regNext_21_0_data_30;
  reg                 io_in_r_bypass_regNext_21_0_load_store_30;
  reg                 io_in_r_bypass_regNext_21_0_df_is_ws_30;
  reg                 io_in_r_bypass_regNext_21_0_stall_30;
  reg        [15:0]   io_in_r_bypass_regNext_21_1_data_30;
  reg                 io_in_r_bypass_regNext_21_1_load_store_30;
  reg                 io_in_r_bypass_regNext_21_1_df_is_ws_30;
  reg                 io_in_r_bypass_regNext_21_1_stall_30;
  reg        [15:0]   io_in_r_bypass_regNext_21_2_data_30;
  reg                 io_in_r_bypass_regNext_21_2_load_store_30;
  reg                 io_in_r_bypass_regNext_21_2_df_is_ws_30;
  reg                 io_in_r_bypass_regNext_21_2_stall_30;
  reg        [15:0]   io_in_r_bypass_regNext_21_3_data_30;
  reg                 io_in_r_bypass_regNext_21_3_load_store_30;
  reg                 io_in_r_bypass_regNext_21_3_df_is_ws_30;
  reg                 io_in_r_bypass_regNext_21_3_stall_30;
  reg        [15:0]   io_in_r_bypass_regNext_22_0_data_30;
  reg                 io_in_r_bypass_regNext_22_0_load_store_30;
  reg                 io_in_r_bypass_regNext_22_0_df_is_ws_30;
  reg                 io_in_r_bypass_regNext_22_0_stall_30;
  reg        [15:0]   io_in_r_bypass_regNext_22_1_data_30;
  reg                 io_in_r_bypass_regNext_22_1_load_store_30;
  reg                 io_in_r_bypass_regNext_22_1_df_is_ws_30;
  reg                 io_in_r_bypass_regNext_22_1_stall_30;
  reg        [15:0]   io_in_r_bypass_regNext_22_2_data_30;
  reg                 io_in_r_bypass_regNext_22_2_load_store_30;
  reg                 io_in_r_bypass_regNext_22_2_df_is_ws_30;
  reg                 io_in_r_bypass_regNext_22_2_stall_30;
  reg        [15:0]   io_in_r_bypass_regNext_22_3_data_30;
  reg                 io_in_r_bypass_regNext_22_3_load_store_30;
  reg                 io_in_r_bypass_regNext_22_3_df_is_ws_30;
  reg                 io_in_r_bypass_regNext_22_3_stall_30;
  reg        [15:0]   io_in_r_bypass_regNext_23_0_data_30;
  reg                 io_in_r_bypass_regNext_23_0_load_store_30;
  reg                 io_in_r_bypass_regNext_23_0_df_is_ws_30;
  reg                 io_in_r_bypass_regNext_23_0_stall_30;
  reg        [15:0]   io_in_r_bypass_regNext_23_1_data_30;
  reg                 io_in_r_bypass_regNext_23_1_load_store_30;
  reg                 io_in_r_bypass_regNext_23_1_df_is_ws_30;
  reg                 io_in_r_bypass_regNext_23_1_stall_30;
  reg        [15:0]   io_in_r_bypass_regNext_23_2_data_30;
  reg                 io_in_r_bypass_regNext_23_2_load_store_30;
  reg                 io_in_r_bypass_regNext_23_2_df_is_ws_30;
  reg                 io_in_r_bypass_regNext_23_2_stall_30;
  reg        [15:0]   io_in_r_bypass_regNext_23_3_data_30;
  reg                 io_in_r_bypass_regNext_23_3_load_store_30;
  reg                 io_in_r_bypass_regNext_23_3_df_is_ws_30;
  reg                 io_in_r_bypass_regNext_23_3_stall_30;
  reg        [15:0]   io_in_r_bypass_regNext_24_0_data_30;
  reg                 io_in_r_bypass_regNext_24_0_load_store_30;
  reg                 io_in_r_bypass_regNext_24_0_df_is_ws_30;
  reg                 io_in_r_bypass_regNext_24_0_stall_30;
  reg        [15:0]   io_in_r_bypass_regNext_24_1_data_30;
  reg                 io_in_r_bypass_regNext_24_1_load_store_30;
  reg                 io_in_r_bypass_regNext_24_1_df_is_ws_30;
  reg                 io_in_r_bypass_regNext_24_1_stall_30;
  reg        [15:0]   io_in_r_bypass_regNext_24_2_data_30;
  reg                 io_in_r_bypass_regNext_24_2_load_store_30;
  reg                 io_in_r_bypass_regNext_24_2_df_is_ws_30;
  reg                 io_in_r_bypass_regNext_24_2_stall_30;
  reg        [15:0]   io_in_r_bypass_regNext_24_3_data_30;
  reg                 io_in_r_bypass_regNext_24_3_load_store_30;
  reg                 io_in_r_bypass_regNext_24_3_df_is_ws_30;
  reg                 io_in_r_bypass_regNext_24_3_stall_30;
  reg        [15:0]   io_in_r_bypass_regNext_25_0_data_30;
  reg                 io_in_r_bypass_regNext_25_0_load_store_30;
  reg                 io_in_r_bypass_regNext_25_0_df_is_ws_30;
  reg                 io_in_r_bypass_regNext_25_0_stall_30;
  reg        [15:0]   io_in_r_bypass_regNext_25_1_data_30;
  reg                 io_in_r_bypass_regNext_25_1_load_store_30;
  reg                 io_in_r_bypass_regNext_25_1_df_is_ws_30;
  reg                 io_in_r_bypass_regNext_25_1_stall_30;
  reg        [15:0]   io_in_r_bypass_regNext_25_2_data_30;
  reg                 io_in_r_bypass_regNext_25_2_load_store_30;
  reg                 io_in_r_bypass_regNext_25_2_df_is_ws_30;
  reg                 io_in_r_bypass_regNext_25_2_stall_30;
  reg        [15:0]   io_in_r_bypass_regNext_25_3_data_30;
  reg                 io_in_r_bypass_regNext_25_3_load_store_30;
  reg                 io_in_r_bypass_regNext_25_3_df_is_ws_30;
  reg                 io_in_r_bypass_regNext_25_3_stall_30;
  reg        [15:0]   io_in_r_bypass_regNext_26_0_data_30;
  reg                 io_in_r_bypass_regNext_26_0_load_store_30;
  reg                 io_in_r_bypass_regNext_26_0_df_is_ws_30;
  reg                 io_in_r_bypass_regNext_26_0_stall_30;
  reg        [15:0]   io_in_r_bypass_regNext_26_1_data_30;
  reg                 io_in_r_bypass_regNext_26_1_load_store_30;
  reg                 io_in_r_bypass_regNext_26_1_df_is_ws_30;
  reg                 io_in_r_bypass_regNext_26_1_stall_30;
  reg        [15:0]   io_in_r_bypass_regNext_26_2_data_30;
  reg                 io_in_r_bypass_regNext_26_2_load_store_30;
  reg                 io_in_r_bypass_regNext_26_2_df_is_ws_30;
  reg                 io_in_r_bypass_regNext_26_2_stall_30;
  reg        [15:0]   io_in_r_bypass_regNext_26_3_data_30;
  reg                 io_in_r_bypass_regNext_26_3_load_store_30;
  reg                 io_in_r_bypass_regNext_26_3_df_is_ws_30;
  reg                 io_in_r_bypass_regNext_26_3_stall_30;
  reg        [15:0]   io_in_r_bypass_regNext_27_0_data_30;
  reg                 io_in_r_bypass_regNext_27_0_load_store_30;
  reg                 io_in_r_bypass_regNext_27_0_df_is_ws_30;
  reg                 io_in_r_bypass_regNext_27_0_stall_30;
  reg        [15:0]   io_in_r_bypass_regNext_27_1_data_30;
  reg                 io_in_r_bypass_regNext_27_1_load_store_30;
  reg                 io_in_r_bypass_regNext_27_1_df_is_ws_30;
  reg                 io_in_r_bypass_regNext_27_1_stall_30;
  reg        [15:0]   io_in_r_bypass_regNext_27_2_data_30;
  reg                 io_in_r_bypass_regNext_27_2_load_store_30;
  reg                 io_in_r_bypass_regNext_27_2_df_is_ws_30;
  reg                 io_in_r_bypass_regNext_27_2_stall_30;
  reg        [15:0]   io_in_r_bypass_regNext_27_3_data_30;
  reg                 io_in_r_bypass_regNext_27_3_load_store_30;
  reg                 io_in_r_bypass_regNext_27_3_df_is_ws_30;
  reg                 io_in_r_bypass_regNext_27_3_stall_30;
  reg        [15:0]   io_in_r_bypass_regNext_28_0_data_30;
  reg                 io_in_r_bypass_regNext_28_0_load_store_30;
  reg                 io_in_r_bypass_regNext_28_0_df_is_ws_30;
  reg                 io_in_r_bypass_regNext_28_0_stall_30;
  reg        [15:0]   io_in_r_bypass_regNext_28_1_data_30;
  reg                 io_in_r_bypass_regNext_28_1_load_store_30;
  reg                 io_in_r_bypass_regNext_28_1_df_is_ws_30;
  reg                 io_in_r_bypass_regNext_28_1_stall_30;
  reg        [15:0]   io_in_r_bypass_regNext_28_2_data_30;
  reg                 io_in_r_bypass_regNext_28_2_load_store_30;
  reg                 io_in_r_bypass_regNext_28_2_df_is_ws_30;
  reg                 io_in_r_bypass_regNext_28_2_stall_30;
  reg        [15:0]   io_in_r_bypass_regNext_28_3_data_30;
  reg                 io_in_r_bypass_regNext_28_3_load_store_30;
  reg                 io_in_r_bypass_regNext_28_3_df_is_ws_30;
  reg                 io_in_r_bypass_regNext_28_3_stall_30;
  reg        [15:0]   io_in_r_bypass_regNext_29_0_data_30;
  reg                 io_in_r_bypass_regNext_29_0_load_store_30;
  reg                 io_in_r_bypass_regNext_29_0_df_is_ws_30;
  reg                 io_in_r_bypass_regNext_29_0_stall_30;
  reg        [15:0]   io_in_r_bypass_regNext_29_1_data_30;
  reg                 io_in_r_bypass_regNext_29_1_load_store_30;
  reg                 io_in_r_bypass_regNext_29_1_df_is_ws_30;
  reg                 io_in_r_bypass_regNext_29_1_stall_30;
  reg        [15:0]   io_in_r_bypass_regNext_29_2_data_30;
  reg                 io_in_r_bypass_regNext_29_2_load_store_30;
  reg                 io_in_r_bypass_regNext_29_2_df_is_ws_30;
  reg                 io_in_r_bypass_regNext_29_2_stall_30;
  reg        [15:0]   io_in_r_bypass_regNext_29_3_data_30;
  reg                 io_in_r_bypass_regNext_29_3_load_store_30;
  reg                 io_in_r_bypass_regNext_29_3_df_is_ws_30;
  reg                 io_in_r_bypass_regNext_29_3_stall_30;
  reg        [15:0]   io_in_r_bypass_regNext_30_0_data_30;
  reg                 io_in_r_bypass_regNext_30_0_load_store_30;
  reg                 io_in_r_bypass_regNext_30_0_df_is_ws_30;
  reg                 io_in_r_bypass_regNext_30_0_stall_30;
  reg        [15:0]   io_in_r_bypass_regNext_30_1_data_30;
  reg                 io_in_r_bypass_regNext_30_1_load_store_30;
  reg                 io_in_r_bypass_regNext_30_1_df_is_ws_30;
  reg                 io_in_r_bypass_regNext_30_1_stall_30;
  reg        [15:0]   io_in_r_bypass_regNext_30_2_data_30;
  reg                 io_in_r_bypass_regNext_30_2_load_store_30;
  reg                 io_in_r_bypass_regNext_30_2_df_is_ws_30;
  reg                 io_in_r_bypass_regNext_30_2_stall_30;
  reg        [15:0]   io_in_r_bypass_regNext_30_3_data_30;
  reg                 io_in_r_bypass_regNext_30_3_load_store_30;
  reg                 io_in_r_bypass_regNext_30_3_df_is_ws_30;
  reg                 io_in_r_bypass_regNext_30_3_stall_30;
  reg        [15:0]   io_in_r_bypass_regNext_31_0_data_30;
  reg                 io_in_r_bypass_regNext_31_0_load_store_30;
  reg                 io_in_r_bypass_regNext_31_0_df_is_ws_30;
  reg                 io_in_r_bypass_regNext_31_0_stall_30;
  reg        [15:0]   io_in_r_bypass_regNext_31_1_data_30;
  reg                 io_in_r_bypass_regNext_31_1_load_store_30;
  reg                 io_in_r_bypass_regNext_31_1_df_is_ws_30;
  reg                 io_in_r_bypass_regNext_31_1_stall_30;
  reg        [15:0]   io_in_r_bypass_regNext_31_2_data_30;
  reg                 io_in_r_bypass_regNext_31_2_load_store_30;
  reg                 io_in_r_bypass_regNext_31_2_df_is_ws_30;
  reg                 io_in_r_bypass_regNext_31_2_stall_30;
  reg        [15:0]   io_in_r_bypass_regNext_31_3_data_30;
  reg                 io_in_r_bypass_regNext_31_3_load_store_30;
  reg                 io_in_r_bypass_regNext_31_3_df_is_ws_30;
  reg                 io_in_r_bypass_regNext_31_3_stall_30;
  reg        [15:0]   io_in_c_bypass_regNext_0_0_data;
  reg                 io_in_c_bypass_regNext_0_0_is_stationary;
  reg        [15:0]   io_in_c_bypass_regNext_0_1_data;
  reg                 io_in_c_bypass_regNext_0_1_is_stationary;
  reg        [15:0]   io_in_c_bypass_regNext_0_2_data;
  reg                 io_in_c_bypass_regNext_0_2_is_stationary;
  reg        [15:0]   io_in_c_bypass_regNext_0_3_data;
  reg                 io_in_c_bypass_regNext_0_3_is_stationary;
  reg        [15:0]   io_in_c_bypass_regNext_1_0_data;
  reg                 io_in_c_bypass_regNext_1_0_is_stationary;
  reg        [15:0]   io_in_c_bypass_regNext_1_1_data;
  reg                 io_in_c_bypass_regNext_1_1_is_stationary;
  reg        [15:0]   io_in_c_bypass_regNext_1_2_data;
  reg                 io_in_c_bypass_regNext_1_2_is_stationary;
  reg        [15:0]   io_in_c_bypass_regNext_1_3_data;
  reg                 io_in_c_bypass_regNext_1_3_is_stationary;
  reg        [15:0]   io_in_c_bypass_regNext_2_0_data;
  reg                 io_in_c_bypass_regNext_2_0_is_stationary;
  reg        [15:0]   io_in_c_bypass_regNext_2_1_data;
  reg                 io_in_c_bypass_regNext_2_1_is_stationary;
  reg        [15:0]   io_in_c_bypass_regNext_2_2_data;
  reg                 io_in_c_bypass_regNext_2_2_is_stationary;
  reg        [15:0]   io_in_c_bypass_regNext_2_3_data;
  reg                 io_in_c_bypass_regNext_2_3_is_stationary;
  reg        [15:0]   io_in_c_bypass_regNext_3_0_data;
  reg                 io_in_c_bypass_regNext_3_0_is_stationary;
  reg        [15:0]   io_in_c_bypass_regNext_3_1_data;
  reg                 io_in_c_bypass_regNext_3_1_is_stationary;
  reg        [15:0]   io_in_c_bypass_regNext_3_2_data;
  reg                 io_in_c_bypass_regNext_3_2_is_stationary;
  reg        [15:0]   io_in_c_bypass_regNext_3_3_data;
  reg                 io_in_c_bypass_regNext_3_3_is_stationary;
  reg        [15:0]   io_in_c_bypass_regNext_4_0_data;
  reg                 io_in_c_bypass_regNext_4_0_is_stationary;
  reg        [15:0]   io_in_c_bypass_regNext_4_1_data;
  reg                 io_in_c_bypass_regNext_4_1_is_stationary;
  reg        [15:0]   io_in_c_bypass_regNext_4_2_data;
  reg                 io_in_c_bypass_regNext_4_2_is_stationary;
  reg        [15:0]   io_in_c_bypass_regNext_4_3_data;
  reg                 io_in_c_bypass_regNext_4_3_is_stationary;
  reg        [15:0]   io_in_c_bypass_regNext_5_0_data;
  reg                 io_in_c_bypass_regNext_5_0_is_stationary;
  reg        [15:0]   io_in_c_bypass_regNext_5_1_data;
  reg                 io_in_c_bypass_regNext_5_1_is_stationary;
  reg        [15:0]   io_in_c_bypass_regNext_5_2_data;
  reg                 io_in_c_bypass_regNext_5_2_is_stationary;
  reg        [15:0]   io_in_c_bypass_regNext_5_3_data;
  reg                 io_in_c_bypass_regNext_5_3_is_stationary;
  reg        [15:0]   io_in_c_bypass_regNext_6_0_data;
  reg                 io_in_c_bypass_regNext_6_0_is_stationary;
  reg        [15:0]   io_in_c_bypass_regNext_6_1_data;
  reg                 io_in_c_bypass_regNext_6_1_is_stationary;
  reg        [15:0]   io_in_c_bypass_regNext_6_2_data;
  reg                 io_in_c_bypass_regNext_6_2_is_stationary;
  reg        [15:0]   io_in_c_bypass_regNext_6_3_data;
  reg                 io_in_c_bypass_regNext_6_3_is_stationary;
  reg        [15:0]   io_in_c_bypass_regNext_7_0_data;
  reg                 io_in_c_bypass_regNext_7_0_is_stationary;
  reg        [15:0]   io_in_c_bypass_regNext_7_1_data;
  reg                 io_in_c_bypass_regNext_7_1_is_stationary;
  reg        [15:0]   io_in_c_bypass_regNext_7_2_data;
  reg                 io_in_c_bypass_regNext_7_2_is_stationary;
  reg        [15:0]   io_in_c_bypass_regNext_7_3_data;
  reg                 io_in_c_bypass_regNext_7_3_is_stationary;
  reg        [15:0]   io_in_c_bypass_regNext_8_0_data;
  reg                 io_in_c_bypass_regNext_8_0_is_stationary;
  reg        [15:0]   io_in_c_bypass_regNext_8_1_data;
  reg                 io_in_c_bypass_regNext_8_1_is_stationary;
  reg        [15:0]   io_in_c_bypass_regNext_8_2_data;
  reg                 io_in_c_bypass_regNext_8_2_is_stationary;
  reg        [15:0]   io_in_c_bypass_regNext_8_3_data;
  reg                 io_in_c_bypass_regNext_8_3_is_stationary;
  reg        [15:0]   io_in_c_bypass_regNext_9_0_data;
  reg                 io_in_c_bypass_regNext_9_0_is_stationary;
  reg        [15:0]   io_in_c_bypass_regNext_9_1_data;
  reg                 io_in_c_bypass_regNext_9_1_is_stationary;
  reg        [15:0]   io_in_c_bypass_regNext_9_2_data;
  reg                 io_in_c_bypass_regNext_9_2_is_stationary;
  reg        [15:0]   io_in_c_bypass_regNext_9_3_data;
  reg                 io_in_c_bypass_regNext_9_3_is_stationary;
  reg        [15:0]   io_in_c_bypass_regNext_10_0_data;
  reg                 io_in_c_bypass_regNext_10_0_is_stationary;
  reg        [15:0]   io_in_c_bypass_regNext_10_1_data;
  reg                 io_in_c_bypass_regNext_10_1_is_stationary;
  reg        [15:0]   io_in_c_bypass_regNext_10_2_data;
  reg                 io_in_c_bypass_regNext_10_2_is_stationary;
  reg        [15:0]   io_in_c_bypass_regNext_10_3_data;
  reg                 io_in_c_bypass_regNext_10_3_is_stationary;
  reg        [15:0]   io_in_c_bypass_regNext_11_0_data;
  reg                 io_in_c_bypass_regNext_11_0_is_stationary;
  reg        [15:0]   io_in_c_bypass_regNext_11_1_data;
  reg                 io_in_c_bypass_regNext_11_1_is_stationary;
  reg        [15:0]   io_in_c_bypass_regNext_11_2_data;
  reg                 io_in_c_bypass_regNext_11_2_is_stationary;
  reg        [15:0]   io_in_c_bypass_regNext_11_3_data;
  reg                 io_in_c_bypass_regNext_11_3_is_stationary;
  reg        [15:0]   io_in_c_bypass_regNext_12_0_data;
  reg                 io_in_c_bypass_regNext_12_0_is_stationary;
  reg        [15:0]   io_in_c_bypass_regNext_12_1_data;
  reg                 io_in_c_bypass_regNext_12_1_is_stationary;
  reg        [15:0]   io_in_c_bypass_regNext_12_2_data;
  reg                 io_in_c_bypass_regNext_12_2_is_stationary;
  reg        [15:0]   io_in_c_bypass_regNext_12_3_data;
  reg                 io_in_c_bypass_regNext_12_3_is_stationary;
  reg        [15:0]   io_in_c_bypass_regNext_13_0_data;
  reg                 io_in_c_bypass_regNext_13_0_is_stationary;
  reg        [15:0]   io_in_c_bypass_regNext_13_1_data;
  reg                 io_in_c_bypass_regNext_13_1_is_stationary;
  reg        [15:0]   io_in_c_bypass_regNext_13_2_data;
  reg                 io_in_c_bypass_regNext_13_2_is_stationary;
  reg        [15:0]   io_in_c_bypass_regNext_13_3_data;
  reg                 io_in_c_bypass_regNext_13_3_is_stationary;
  reg        [15:0]   io_in_c_bypass_regNext_14_0_data;
  reg                 io_in_c_bypass_regNext_14_0_is_stationary;
  reg        [15:0]   io_in_c_bypass_regNext_14_1_data;
  reg                 io_in_c_bypass_regNext_14_1_is_stationary;
  reg        [15:0]   io_in_c_bypass_regNext_14_2_data;
  reg                 io_in_c_bypass_regNext_14_2_is_stationary;
  reg        [15:0]   io_in_c_bypass_regNext_14_3_data;
  reg                 io_in_c_bypass_regNext_14_3_is_stationary;
  reg        [15:0]   io_in_c_bypass_regNext_15_0_data;
  reg                 io_in_c_bypass_regNext_15_0_is_stationary;
  reg        [15:0]   io_in_c_bypass_regNext_15_1_data;
  reg                 io_in_c_bypass_regNext_15_1_is_stationary;
  reg        [15:0]   io_in_c_bypass_regNext_15_2_data;
  reg                 io_in_c_bypass_regNext_15_2_is_stationary;
  reg        [15:0]   io_in_c_bypass_regNext_15_3_data;
  reg                 io_in_c_bypass_regNext_15_3_is_stationary;
  reg        [15:0]   io_in_c_bypass_regNext_16_0_data;
  reg                 io_in_c_bypass_regNext_16_0_is_stationary;
  reg        [15:0]   io_in_c_bypass_regNext_16_1_data;
  reg                 io_in_c_bypass_regNext_16_1_is_stationary;
  reg        [15:0]   io_in_c_bypass_regNext_16_2_data;
  reg                 io_in_c_bypass_regNext_16_2_is_stationary;
  reg        [15:0]   io_in_c_bypass_regNext_16_3_data;
  reg                 io_in_c_bypass_regNext_16_3_is_stationary;
  reg        [15:0]   io_in_c_bypass_regNext_17_0_data;
  reg                 io_in_c_bypass_regNext_17_0_is_stationary;
  reg        [15:0]   io_in_c_bypass_regNext_17_1_data;
  reg                 io_in_c_bypass_regNext_17_1_is_stationary;
  reg        [15:0]   io_in_c_bypass_regNext_17_2_data;
  reg                 io_in_c_bypass_regNext_17_2_is_stationary;
  reg        [15:0]   io_in_c_bypass_regNext_17_3_data;
  reg                 io_in_c_bypass_regNext_17_3_is_stationary;
  reg        [15:0]   io_in_c_bypass_regNext_18_0_data;
  reg                 io_in_c_bypass_regNext_18_0_is_stationary;
  reg        [15:0]   io_in_c_bypass_regNext_18_1_data;
  reg                 io_in_c_bypass_regNext_18_1_is_stationary;
  reg        [15:0]   io_in_c_bypass_regNext_18_2_data;
  reg                 io_in_c_bypass_regNext_18_2_is_stationary;
  reg        [15:0]   io_in_c_bypass_regNext_18_3_data;
  reg                 io_in_c_bypass_regNext_18_3_is_stationary;
  reg        [15:0]   io_in_c_bypass_regNext_19_0_data;
  reg                 io_in_c_bypass_regNext_19_0_is_stationary;
  reg        [15:0]   io_in_c_bypass_regNext_19_1_data;
  reg                 io_in_c_bypass_regNext_19_1_is_stationary;
  reg        [15:0]   io_in_c_bypass_regNext_19_2_data;
  reg                 io_in_c_bypass_regNext_19_2_is_stationary;
  reg        [15:0]   io_in_c_bypass_regNext_19_3_data;
  reg                 io_in_c_bypass_regNext_19_3_is_stationary;
  reg        [15:0]   io_in_c_bypass_regNext_20_0_data;
  reg                 io_in_c_bypass_regNext_20_0_is_stationary;
  reg        [15:0]   io_in_c_bypass_regNext_20_1_data;
  reg                 io_in_c_bypass_regNext_20_1_is_stationary;
  reg        [15:0]   io_in_c_bypass_regNext_20_2_data;
  reg                 io_in_c_bypass_regNext_20_2_is_stationary;
  reg        [15:0]   io_in_c_bypass_regNext_20_3_data;
  reg                 io_in_c_bypass_regNext_20_3_is_stationary;
  reg        [15:0]   io_in_c_bypass_regNext_21_0_data;
  reg                 io_in_c_bypass_regNext_21_0_is_stationary;
  reg        [15:0]   io_in_c_bypass_regNext_21_1_data;
  reg                 io_in_c_bypass_regNext_21_1_is_stationary;
  reg        [15:0]   io_in_c_bypass_regNext_21_2_data;
  reg                 io_in_c_bypass_regNext_21_2_is_stationary;
  reg        [15:0]   io_in_c_bypass_regNext_21_3_data;
  reg                 io_in_c_bypass_regNext_21_3_is_stationary;
  reg        [15:0]   io_in_c_bypass_regNext_22_0_data;
  reg                 io_in_c_bypass_regNext_22_0_is_stationary;
  reg        [15:0]   io_in_c_bypass_regNext_22_1_data;
  reg                 io_in_c_bypass_regNext_22_1_is_stationary;
  reg        [15:0]   io_in_c_bypass_regNext_22_2_data;
  reg                 io_in_c_bypass_regNext_22_2_is_stationary;
  reg        [15:0]   io_in_c_bypass_regNext_22_3_data;
  reg                 io_in_c_bypass_regNext_22_3_is_stationary;
  reg        [15:0]   io_in_c_bypass_regNext_23_0_data;
  reg                 io_in_c_bypass_regNext_23_0_is_stationary;
  reg        [15:0]   io_in_c_bypass_regNext_23_1_data;
  reg                 io_in_c_bypass_regNext_23_1_is_stationary;
  reg        [15:0]   io_in_c_bypass_regNext_23_2_data;
  reg                 io_in_c_bypass_regNext_23_2_is_stationary;
  reg        [15:0]   io_in_c_bypass_regNext_23_3_data;
  reg                 io_in_c_bypass_regNext_23_3_is_stationary;
  reg        [15:0]   io_in_c_bypass_regNext_24_0_data;
  reg                 io_in_c_bypass_regNext_24_0_is_stationary;
  reg        [15:0]   io_in_c_bypass_regNext_24_1_data;
  reg                 io_in_c_bypass_regNext_24_1_is_stationary;
  reg        [15:0]   io_in_c_bypass_regNext_24_2_data;
  reg                 io_in_c_bypass_regNext_24_2_is_stationary;
  reg        [15:0]   io_in_c_bypass_regNext_24_3_data;
  reg                 io_in_c_bypass_regNext_24_3_is_stationary;
  reg        [15:0]   io_in_c_bypass_regNext_25_0_data;
  reg                 io_in_c_bypass_regNext_25_0_is_stationary;
  reg        [15:0]   io_in_c_bypass_regNext_25_1_data;
  reg                 io_in_c_bypass_regNext_25_1_is_stationary;
  reg        [15:0]   io_in_c_bypass_regNext_25_2_data;
  reg                 io_in_c_bypass_regNext_25_2_is_stationary;
  reg        [15:0]   io_in_c_bypass_regNext_25_3_data;
  reg                 io_in_c_bypass_regNext_25_3_is_stationary;
  reg        [15:0]   io_in_c_bypass_regNext_26_0_data;
  reg                 io_in_c_bypass_regNext_26_0_is_stationary;
  reg        [15:0]   io_in_c_bypass_regNext_26_1_data;
  reg                 io_in_c_bypass_regNext_26_1_is_stationary;
  reg        [15:0]   io_in_c_bypass_regNext_26_2_data;
  reg                 io_in_c_bypass_regNext_26_2_is_stationary;
  reg        [15:0]   io_in_c_bypass_regNext_26_3_data;
  reg                 io_in_c_bypass_regNext_26_3_is_stationary;
  reg        [15:0]   io_in_c_bypass_regNext_27_0_data;
  reg                 io_in_c_bypass_regNext_27_0_is_stationary;
  reg        [15:0]   io_in_c_bypass_regNext_27_1_data;
  reg                 io_in_c_bypass_regNext_27_1_is_stationary;
  reg        [15:0]   io_in_c_bypass_regNext_27_2_data;
  reg                 io_in_c_bypass_regNext_27_2_is_stationary;
  reg        [15:0]   io_in_c_bypass_regNext_27_3_data;
  reg                 io_in_c_bypass_regNext_27_3_is_stationary;
  reg        [15:0]   io_in_c_bypass_regNext_28_0_data;
  reg                 io_in_c_bypass_regNext_28_0_is_stationary;
  reg        [15:0]   io_in_c_bypass_regNext_28_1_data;
  reg                 io_in_c_bypass_regNext_28_1_is_stationary;
  reg        [15:0]   io_in_c_bypass_regNext_28_2_data;
  reg                 io_in_c_bypass_regNext_28_2_is_stationary;
  reg        [15:0]   io_in_c_bypass_regNext_28_3_data;
  reg                 io_in_c_bypass_regNext_28_3_is_stationary;
  reg        [15:0]   io_in_c_bypass_regNext_29_0_data;
  reg                 io_in_c_bypass_regNext_29_0_is_stationary;
  reg        [15:0]   io_in_c_bypass_regNext_29_1_data;
  reg                 io_in_c_bypass_regNext_29_1_is_stationary;
  reg        [15:0]   io_in_c_bypass_regNext_29_2_data;
  reg                 io_in_c_bypass_regNext_29_2_is_stationary;
  reg        [15:0]   io_in_c_bypass_regNext_29_3_data;
  reg                 io_in_c_bypass_regNext_29_3_is_stationary;
  reg        [15:0]   io_in_c_bypass_regNext_30_0_data;
  reg                 io_in_c_bypass_regNext_30_0_is_stationary;
  reg        [15:0]   io_in_c_bypass_regNext_30_1_data;
  reg                 io_in_c_bypass_regNext_30_1_is_stationary;
  reg        [15:0]   io_in_c_bypass_regNext_30_2_data;
  reg                 io_in_c_bypass_regNext_30_2_is_stationary;
  reg        [15:0]   io_in_c_bypass_regNext_30_3_data;
  reg                 io_in_c_bypass_regNext_30_3_is_stationary;
  reg        [15:0]   io_in_c_bypass_regNext_31_0_data;
  reg                 io_in_c_bypass_regNext_31_0_is_stationary;
  reg        [15:0]   io_in_c_bypass_regNext_31_1_data;
  reg                 io_in_c_bypass_regNext_31_1_is_stationary;
  reg        [15:0]   io_in_c_bypass_regNext_31_2_data;
  reg                 io_in_c_bypass_regNext_31_2_is_stationary;
  reg        [15:0]   io_in_c_bypass_regNext_31_3_data;
  reg                 io_in_c_bypass_regNext_31_3_is_stationary;
  reg        [15:0]   io_in_c_bypass_regNext_0_0_data_1;
  reg                 io_in_c_bypass_regNext_0_0_is_stationary_1;
  reg        [15:0]   io_in_c_bypass_regNext_0_1_data_1;
  reg                 io_in_c_bypass_regNext_0_1_is_stationary_1;
  reg        [15:0]   io_in_c_bypass_regNext_0_2_data_1;
  reg                 io_in_c_bypass_regNext_0_2_is_stationary_1;
  reg        [15:0]   io_in_c_bypass_regNext_0_3_data_1;
  reg                 io_in_c_bypass_regNext_0_3_is_stationary_1;
  reg        [15:0]   io_in_c_bypass_regNext_1_0_data_1;
  reg                 io_in_c_bypass_regNext_1_0_is_stationary_1;
  reg        [15:0]   io_in_c_bypass_regNext_1_1_data_1;
  reg                 io_in_c_bypass_regNext_1_1_is_stationary_1;
  reg        [15:0]   io_in_c_bypass_regNext_1_2_data_1;
  reg                 io_in_c_bypass_regNext_1_2_is_stationary_1;
  reg        [15:0]   io_in_c_bypass_regNext_1_3_data_1;
  reg                 io_in_c_bypass_regNext_1_3_is_stationary_1;
  reg        [15:0]   io_in_c_bypass_regNext_2_0_data_1;
  reg                 io_in_c_bypass_regNext_2_0_is_stationary_1;
  reg        [15:0]   io_in_c_bypass_regNext_2_1_data_1;
  reg                 io_in_c_bypass_regNext_2_1_is_stationary_1;
  reg        [15:0]   io_in_c_bypass_regNext_2_2_data_1;
  reg                 io_in_c_bypass_regNext_2_2_is_stationary_1;
  reg        [15:0]   io_in_c_bypass_regNext_2_3_data_1;
  reg                 io_in_c_bypass_regNext_2_3_is_stationary_1;
  reg        [15:0]   io_in_c_bypass_regNext_3_0_data_1;
  reg                 io_in_c_bypass_regNext_3_0_is_stationary_1;
  reg        [15:0]   io_in_c_bypass_regNext_3_1_data_1;
  reg                 io_in_c_bypass_regNext_3_1_is_stationary_1;
  reg        [15:0]   io_in_c_bypass_regNext_3_2_data_1;
  reg                 io_in_c_bypass_regNext_3_2_is_stationary_1;
  reg        [15:0]   io_in_c_bypass_regNext_3_3_data_1;
  reg                 io_in_c_bypass_regNext_3_3_is_stationary_1;
  reg        [15:0]   io_in_c_bypass_regNext_4_0_data_1;
  reg                 io_in_c_bypass_regNext_4_0_is_stationary_1;
  reg        [15:0]   io_in_c_bypass_regNext_4_1_data_1;
  reg                 io_in_c_bypass_regNext_4_1_is_stationary_1;
  reg        [15:0]   io_in_c_bypass_regNext_4_2_data_1;
  reg                 io_in_c_bypass_regNext_4_2_is_stationary_1;
  reg        [15:0]   io_in_c_bypass_regNext_4_3_data_1;
  reg                 io_in_c_bypass_regNext_4_3_is_stationary_1;
  reg        [15:0]   io_in_c_bypass_regNext_5_0_data_1;
  reg                 io_in_c_bypass_regNext_5_0_is_stationary_1;
  reg        [15:0]   io_in_c_bypass_regNext_5_1_data_1;
  reg                 io_in_c_bypass_regNext_5_1_is_stationary_1;
  reg        [15:0]   io_in_c_bypass_regNext_5_2_data_1;
  reg                 io_in_c_bypass_regNext_5_2_is_stationary_1;
  reg        [15:0]   io_in_c_bypass_regNext_5_3_data_1;
  reg                 io_in_c_bypass_regNext_5_3_is_stationary_1;
  reg        [15:0]   io_in_c_bypass_regNext_6_0_data_1;
  reg                 io_in_c_bypass_regNext_6_0_is_stationary_1;
  reg        [15:0]   io_in_c_bypass_regNext_6_1_data_1;
  reg                 io_in_c_bypass_regNext_6_1_is_stationary_1;
  reg        [15:0]   io_in_c_bypass_regNext_6_2_data_1;
  reg                 io_in_c_bypass_regNext_6_2_is_stationary_1;
  reg        [15:0]   io_in_c_bypass_regNext_6_3_data_1;
  reg                 io_in_c_bypass_regNext_6_3_is_stationary_1;
  reg        [15:0]   io_in_c_bypass_regNext_7_0_data_1;
  reg                 io_in_c_bypass_regNext_7_0_is_stationary_1;
  reg        [15:0]   io_in_c_bypass_regNext_7_1_data_1;
  reg                 io_in_c_bypass_regNext_7_1_is_stationary_1;
  reg        [15:0]   io_in_c_bypass_regNext_7_2_data_1;
  reg                 io_in_c_bypass_regNext_7_2_is_stationary_1;
  reg        [15:0]   io_in_c_bypass_regNext_7_3_data_1;
  reg                 io_in_c_bypass_regNext_7_3_is_stationary_1;
  reg        [15:0]   io_in_c_bypass_regNext_8_0_data_1;
  reg                 io_in_c_bypass_regNext_8_0_is_stationary_1;
  reg        [15:0]   io_in_c_bypass_regNext_8_1_data_1;
  reg                 io_in_c_bypass_regNext_8_1_is_stationary_1;
  reg        [15:0]   io_in_c_bypass_regNext_8_2_data_1;
  reg                 io_in_c_bypass_regNext_8_2_is_stationary_1;
  reg        [15:0]   io_in_c_bypass_regNext_8_3_data_1;
  reg                 io_in_c_bypass_regNext_8_3_is_stationary_1;
  reg        [15:0]   io_in_c_bypass_regNext_9_0_data_1;
  reg                 io_in_c_bypass_regNext_9_0_is_stationary_1;
  reg        [15:0]   io_in_c_bypass_regNext_9_1_data_1;
  reg                 io_in_c_bypass_regNext_9_1_is_stationary_1;
  reg        [15:0]   io_in_c_bypass_regNext_9_2_data_1;
  reg                 io_in_c_bypass_regNext_9_2_is_stationary_1;
  reg        [15:0]   io_in_c_bypass_regNext_9_3_data_1;
  reg                 io_in_c_bypass_regNext_9_3_is_stationary_1;
  reg        [15:0]   io_in_c_bypass_regNext_10_0_data_1;
  reg                 io_in_c_bypass_regNext_10_0_is_stationary_1;
  reg        [15:0]   io_in_c_bypass_regNext_10_1_data_1;
  reg                 io_in_c_bypass_regNext_10_1_is_stationary_1;
  reg        [15:0]   io_in_c_bypass_regNext_10_2_data_1;
  reg                 io_in_c_bypass_regNext_10_2_is_stationary_1;
  reg        [15:0]   io_in_c_bypass_regNext_10_3_data_1;
  reg                 io_in_c_bypass_regNext_10_3_is_stationary_1;
  reg        [15:0]   io_in_c_bypass_regNext_11_0_data_1;
  reg                 io_in_c_bypass_regNext_11_0_is_stationary_1;
  reg        [15:0]   io_in_c_bypass_regNext_11_1_data_1;
  reg                 io_in_c_bypass_regNext_11_1_is_stationary_1;
  reg        [15:0]   io_in_c_bypass_regNext_11_2_data_1;
  reg                 io_in_c_bypass_regNext_11_2_is_stationary_1;
  reg        [15:0]   io_in_c_bypass_regNext_11_3_data_1;
  reg                 io_in_c_bypass_regNext_11_3_is_stationary_1;
  reg        [15:0]   io_in_c_bypass_regNext_12_0_data_1;
  reg                 io_in_c_bypass_regNext_12_0_is_stationary_1;
  reg        [15:0]   io_in_c_bypass_regNext_12_1_data_1;
  reg                 io_in_c_bypass_regNext_12_1_is_stationary_1;
  reg        [15:0]   io_in_c_bypass_regNext_12_2_data_1;
  reg                 io_in_c_bypass_regNext_12_2_is_stationary_1;
  reg        [15:0]   io_in_c_bypass_regNext_12_3_data_1;
  reg                 io_in_c_bypass_regNext_12_3_is_stationary_1;
  reg        [15:0]   io_in_c_bypass_regNext_13_0_data_1;
  reg                 io_in_c_bypass_regNext_13_0_is_stationary_1;
  reg        [15:0]   io_in_c_bypass_regNext_13_1_data_1;
  reg                 io_in_c_bypass_regNext_13_1_is_stationary_1;
  reg        [15:0]   io_in_c_bypass_regNext_13_2_data_1;
  reg                 io_in_c_bypass_regNext_13_2_is_stationary_1;
  reg        [15:0]   io_in_c_bypass_regNext_13_3_data_1;
  reg                 io_in_c_bypass_regNext_13_3_is_stationary_1;
  reg        [15:0]   io_in_c_bypass_regNext_14_0_data_1;
  reg                 io_in_c_bypass_regNext_14_0_is_stationary_1;
  reg        [15:0]   io_in_c_bypass_regNext_14_1_data_1;
  reg                 io_in_c_bypass_regNext_14_1_is_stationary_1;
  reg        [15:0]   io_in_c_bypass_regNext_14_2_data_1;
  reg                 io_in_c_bypass_regNext_14_2_is_stationary_1;
  reg        [15:0]   io_in_c_bypass_regNext_14_3_data_1;
  reg                 io_in_c_bypass_regNext_14_3_is_stationary_1;
  reg        [15:0]   io_in_c_bypass_regNext_15_0_data_1;
  reg                 io_in_c_bypass_regNext_15_0_is_stationary_1;
  reg        [15:0]   io_in_c_bypass_regNext_15_1_data_1;
  reg                 io_in_c_bypass_regNext_15_1_is_stationary_1;
  reg        [15:0]   io_in_c_bypass_regNext_15_2_data_1;
  reg                 io_in_c_bypass_regNext_15_2_is_stationary_1;
  reg        [15:0]   io_in_c_bypass_regNext_15_3_data_1;
  reg                 io_in_c_bypass_regNext_15_3_is_stationary_1;
  reg        [15:0]   io_in_c_bypass_regNext_16_0_data_1;
  reg                 io_in_c_bypass_regNext_16_0_is_stationary_1;
  reg        [15:0]   io_in_c_bypass_regNext_16_1_data_1;
  reg                 io_in_c_bypass_regNext_16_1_is_stationary_1;
  reg        [15:0]   io_in_c_bypass_regNext_16_2_data_1;
  reg                 io_in_c_bypass_regNext_16_2_is_stationary_1;
  reg        [15:0]   io_in_c_bypass_regNext_16_3_data_1;
  reg                 io_in_c_bypass_regNext_16_3_is_stationary_1;
  reg        [15:0]   io_in_c_bypass_regNext_17_0_data_1;
  reg                 io_in_c_bypass_regNext_17_0_is_stationary_1;
  reg        [15:0]   io_in_c_bypass_regNext_17_1_data_1;
  reg                 io_in_c_bypass_regNext_17_1_is_stationary_1;
  reg        [15:0]   io_in_c_bypass_regNext_17_2_data_1;
  reg                 io_in_c_bypass_regNext_17_2_is_stationary_1;
  reg        [15:0]   io_in_c_bypass_regNext_17_3_data_1;
  reg                 io_in_c_bypass_regNext_17_3_is_stationary_1;
  reg        [15:0]   io_in_c_bypass_regNext_18_0_data_1;
  reg                 io_in_c_bypass_regNext_18_0_is_stationary_1;
  reg        [15:0]   io_in_c_bypass_regNext_18_1_data_1;
  reg                 io_in_c_bypass_regNext_18_1_is_stationary_1;
  reg        [15:0]   io_in_c_bypass_regNext_18_2_data_1;
  reg                 io_in_c_bypass_regNext_18_2_is_stationary_1;
  reg        [15:0]   io_in_c_bypass_regNext_18_3_data_1;
  reg                 io_in_c_bypass_regNext_18_3_is_stationary_1;
  reg        [15:0]   io_in_c_bypass_regNext_19_0_data_1;
  reg                 io_in_c_bypass_regNext_19_0_is_stationary_1;
  reg        [15:0]   io_in_c_bypass_regNext_19_1_data_1;
  reg                 io_in_c_bypass_regNext_19_1_is_stationary_1;
  reg        [15:0]   io_in_c_bypass_regNext_19_2_data_1;
  reg                 io_in_c_bypass_regNext_19_2_is_stationary_1;
  reg        [15:0]   io_in_c_bypass_regNext_19_3_data_1;
  reg                 io_in_c_bypass_regNext_19_3_is_stationary_1;
  reg        [15:0]   io_in_c_bypass_regNext_20_0_data_1;
  reg                 io_in_c_bypass_regNext_20_0_is_stationary_1;
  reg        [15:0]   io_in_c_bypass_regNext_20_1_data_1;
  reg                 io_in_c_bypass_regNext_20_1_is_stationary_1;
  reg        [15:0]   io_in_c_bypass_regNext_20_2_data_1;
  reg                 io_in_c_bypass_regNext_20_2_is_stationary_1;
  reg        [15:0]   io_in_c_bypass_regNext_20_3_data_1;
  reg                 io_in_c_bypass_regNext_20_3_is_stationary_1;
  reg        [15:0]   io_in_c_bypass_regNext_21_0_data_1;
  reg                 io_in_c_bypass_regNext_21_0_is_stationary_1;
  reg        [15:0]   io_in_c_bypass_regNext_21_1_data_1;
  reg                 io_in_c_bypass_regNext_21_1_is_stationary_1;
  reg        [15:0]   io_in_c_bypass_regNext_21_2_data_1;
  reg                 io_in_c_bypass_regNext_21_2_is_stationary_1;
  reg        [15:0]   io_in_c_bypass_regNext_21_3_data_1;
  reg                 io_in_c_bypass_regNext_21_3_is_stationary_1;
  reg        [15:0]   io_in_c_bypass_regNext_22_0_data_1;
  reg                 io_in_c_bypass_regNext_22_0_is_stationary_1;
  reg        [15:0]   io_in_c_bypass_regNext_22_1_data_1;
  reg                 io_in_c_bypass_regNext_22_1_is_stationary_1;
  reg        [15:0]   io_in_c_bypass_regNext_22_2_data_1;
  reg                 io_in_c_bypass_regNext_22_2_is_stationary_1;
  reg        [15:0]   io_in_c_bypass_regNext_22_3_data_1;
  reg                 io_in_c_bypass_regNext_22_3_is_stationary_1;
  reg        [15:0]   io_in_c_bypass_regNext_23_0_data_1;
  reg                 io_in_c_bypass_regNext_23_0_is_stationary_1;
  reg        [15:0]   io_in_c_bypass_regNext_23_1_data_1;
  reg                 io_in_c_bypass_regNext_23_1_is_stationary_1;
  reg        [15:0]   io_in_c_bypass_regNext_23_2_data_1;
  reg                 io_in_c_bypass_regNext_23_2_is_stationary_1;
  reg        [15:0]   io_in_c_bypass_regNext_23_3_data_1;
  reg                 io_in_c_bypass_regNext_23_3_is_stationary_1;
  reg        [15:0]   io_in_c_bypass_regNext_24_0_data_1;
  reg                 io_in_c_bypass_regNext_24_0_is_stationary_1;
  reg        [15:0]   io_in_c_bypass_regNext_24_1_data_1;
  reg                 io_in_c_bypass_regNext_24_1_is_stationary_1;
  reg        [15:0]   io_in_c_bypass_regNext_24_2_data_1;
  reg                 io_in_c_bypass_regNext_24_2_is_stationary_1;
  reg        [15:0]   io_in_c_bypass_regNext_24_3_data_1;
  reg                 io_in_c_bypass_regNext_24_3_is_stationary_1;
  reg        [15:0]   io_in_c_bypass_regNext_25_0_data_1;
  reg                 io_in_c_bypass_regNext_25_0_is_stationary_1;
  reg        [15:0]   io_in_c_bypass_regNext_25_1_data_1;
  reg                 io_in_c_bypass_regNext_25_1_is_stationary_1;
  reg        [15:0]   io_in_c_bypass_regNext_25_2_data_1;
  reg                 io_in_c_bypass_regNext_25_2_is_stationary_1;
  reg        [15:0]   io_in_c_bypass_regNext_25_3_data_1;
  reg                 io_in_c_bypass_regNext_25_3_is_stationary_1;
  reg        [15:0]   io_in_c_bypass_regNext_26_0_data_1;
  reg                 io_in_c_bypass_regNext_26_0_is_stationary_1;
  reg        [15:0]   io_in_c_bypass_regNext_26_1_data_1;
  reg                 io_in_c_bypass_regNext_26_1_is_stationary_1;
  reg        [15:0]   io_in_c_bypass_regNext_26_2_data_1;
  reg                 io_in_c_bypass_regNext_26_2_is_stationary_1;
  reg        [15:0]   io_in_c_bypass_regNext_26_3_data_1;
  reg                 io_in_c_bypass_regNext_26_3_is_stationary_1;
  reg        [15:0]   io_in_c_bypass_regNext_27_0_data_1;
  reg                 io_in_c_bypass_regNext_27_0_is_stationary_1;
  reg        [15:0]   io_in_c_bypass_regNext_27_1_data_1;
  reg                 io_in_c_bypass_regNext_27_1_is_stationary_1;
  reg        [15:0]   io_in_c_bypass_regNext_27_2_data_1;
  reg                 io_in_c_bypass_regNext_27_2_is_stationary_1;
  reg        [15:0]   io_in_c_bypass_regNext_27_3_data_1;
  reg                 io_in_c_bypass_regNext_27_3_is_stationary_1;
  reg        [15:0]   io_in_c_bypass_regNext_28_0_data_1;
  reg                 io_in_c_bypass_regNext_28_0_is_stationary_1;
  reg        [15:0]   io_in_c_bypass_regNext_28_1_data_1;
  reg                 io_in_c_bypass_regNext_28_1_is_stationary_1;
  reg        [15:0]   io_in_c_bypass_regNext_28_2_data_1;
  reg                 io_in_c_bypass_regNext_28_2_is_stationary_1;
  reg        [15:0]   io_in_c_bypass_regNext_28_3_data_1;
  reg                 io_in_c_bypass_regNext_28_3_is_stationary_1;
  reg        [15:0]   io_in_c_bypass_regNext_29_0_data_1;
  reg                 io_in_c_bypass_regNext_29_0_is_stationary_1;
  reg        [15:0]   io_in_c_bypass_regNext_29_1_data_1;
  reg                 io_in_c_bypass_regNext_29_1_is_stationary_1;
  reg        [15:0]   io_in_c_bypass_regNext_29_2_data_1;
  reg                 io_in_c_bypass_regNext_29_2_is_stationary_1;
  reg        [15:0]   io_in_c_bypass_regNext_29_3_data_1;
  reg                 io_in_c_bypass_regNext_29_3_is_stationary_1;
  reg        [15:0]   io_in_c_bypass_regNext_30_0_data_1;
  reg                 io_in_c_bypass_regNext_30_0_is_stationary_1;
  reg        [15:0]   io_in_c_bypass_regNext_30_1_data_1;
  reg                 io_in_c_bypass_regNext_30_1_is_stationary_1;
  reg        [15:0]   io_in_c_bypass_regNext_30_2_data_1;
  reg                 io_in_c_bypass_regNext_30_2_is_stationary_1;
  reg        [15:0]   io_in_c_bypass_regNext_30_3_data_1;
  reg                 io_in_c_bypass_regNext_30_3_is_stationary_1;
  reg        [15:0]   io_in_c_bypass_regNext_31_0_data_1;
  reg                 io_in_c_bypass_regNext_31_0_is_stationary_1;
  reg        [15:0]   io_in_c_bypass_regNext_31_1_data_1;
  reg                 io_in_c_bypass_regNext_31_1_is_stationary_1;
  reg        [15:0]   io_in_c_bypass_regNext_31_2_data_1;
  reg                 io_in_c_bypass_regNext_31_2_is_stationary_1;
  reg        [15:0]   io_in_c_bypass_regNext_31_3_data_1;
  reg                 io_in_c_bypass_regNext_31_3_is_stationary_1;
  reg        [15:0]   io_in_c_bypass_regNext_0_0_data_2;
  reg                 io_in_c_bypass_regNext_0_0_is_stationary_2;
  reg        [15:0]   io_in_c_bypass_regNext_0_1_data_2;
  reg                 io_in_c_bypass_regNext_0_1_is_stationary_2;
  reg        [15:0]   io_in_c_bypass_regNext_0_2_data_2;
  reg                 io_in_c_bypass_regNext_0_2_is_stationary_2;
  reg        [15:0]   io_in_c_bypass_regNext_0_3_data_2;
  reg                 io_in_c_bypass_regNext_0_3_is_stationary_2;
  reg        [15:0]   io_in_c_bypass_regNext_1_0_data_2;
  reg                 io_in_c_bypass_regNext_1_0_is_stationary_2;
  reg        [15:0]   io_in_c_bypass_regNext_1_1_data_2;
  reg                 io_in_c_bypass_regNext_1_1_is_stationary_2;
  reg        [15:0]   io_in_c_bypass_regNext_1_2_data_2;
  reg                 io_in_c_bypass_regNext_1_2_is_stationary_2;
  reg        [15:0]   io_in_c_bypass_regNext_1_3_data_2;
  reg                 io_in_c_bypass_regNext_1_3_is_stationary_2;
  reg        [15:0]   io_in_c_bypass_regNext_2_0_data_2;
  reg                 io_in_c_bypass_regNext_2_0_is_stationary_2;
  reg        [15:0]   io_in_c_bypass_regNext_2_1_data_2;
  reg                 io_in_c_bypass_regNext_2_1_is_stationary_2;
  reg        [15:0]   io_in_c_bypass_regNext_2_2_data_2;
  reg                 io_in_c_bypass_regNext_2_2_is_stationary_2;
  reg        [15:0]   io_in_c_bypass_regNext_2_3_data_2;
  reg                 io_in_c_bypass_regNext_2_3_is_stationary_2;
  reg        [15:0]   io_in_c_bypass_regNext_3_0_data_2;
  reg                 io_in_c_bypass_regNext_3_0_is_stationary_2;
  reg        [15:0]   io_in_c_bypass_regNext_3_1_data_2;
  reg                 io_in_c_bypass_regNext_3_1_is_stationary_2;
  reg        [15:0]   io_in_c_bypass_regNext_3_2_data_2;
  reg                 io_in_c_bypass_regNext_3_2_is_stationary_2;
  reg        [15:0]   io_in_c_bypass_regNext_3_3_data_2;
  reg                 io_in_c_bypass_regNext_3_3_is_stationary_2;
  reg        [15:0]   io_in_c_bypass_regNext_4_0_data_2;
  reg                 io_in_c_bypass_regNext_4_0_is_stationary_2;
  reg        [15:0]   io_in_c_bypass_regNext_4_1_data_2;
  reg                 io_in_c_bypass_regNext_4_1_is_stationary_2;
  reg        [15:0]   io_in_c_bypass_regNext_4_2_data_2;
  reg                 io_in_c_bypass_regNext_4_2_is_stationary_2;
  reg        [15:0]   io_in_c_bypass_regNext_4_3_data_2;
  reg                 io_in_c_bypass_regNext_4_3_is_stationary_2;
  reg        [15:0]   io_in_c_bypass_regNext_5_0_data_2;
  reg                 io_in_c_bypass_regNext_5_0_is_stationary_2;
  reg        [15:0]   io_in_c_bypass_regNext_5_1_data_2;
  reg                 io_in_c_bypass_regNext_5_1_is_stationary_2;
  reg        [15:0]   io_in_c_bypass_regNext_5_2_data_2;
  reg                 io_in_c_bypass_regNext_5_2_is_stationary_2;
  reg        [15:0]   io_in_c_bypass_regNext_5_3_data_2;
  reg                 io_in_c_bypass_regNext_5_3_is_stationary_2;
  reg        [15:0]   io_in_c_bypass_regNext_6_0_data_2;
  reg                 io_in_c_bypass_regNext_6_0_is_stationary_2;
  reg        [15:0]   io_in_c_bypass_regNext_6_1_data_2;
  reg                 io_in_c_bypass_regNext_6_1_is_stationary_2;
  reg        [15:0]   io_in_c_bypass_regNext_6_2_data_2;
  reg                 io_in_c_bypass_regNext_6_2_is_stationary_2;
  reg        [15:0]   io_in_c_bypass_regNext_6_3_data_2;
  reg                 io_in_c_bypass_regNext_6_3_is_stationary_2;
  reg        [15:0]   io_in_c_bypass_regNext_7_0_data_2;
  reg                 io_in_c_bypass_regNext_7_0_is_stationary_2;
  reg        [15:0]   io_in_c_bypass_regNext_7_1_data_2;
  reg                 io_in_c_bypass_regNext_7_1_is_stationary_2;
  reg        [15:0]   io_in_c_bypass_regNext_7_2_data_2;
  reg                 io_in_c_bypass_regNext_7_2_is_stationary_2;
  reg        [15:0]   io_in_c_bypass_regNext_7_3_data_2;
  reg                 io_in_c_bypass_regNext_7_3_is_stationary_2;
  reg        [15:0]   io_in_c_bypass_regNext_8_0_data_2;
  reg                 io_in_c_bypass_regNext_8_0_is_stationary_2;
  reg        [15:0]   io_in_c_bypass_regNext_8_1_data_2;
  reg                 io_in_c_bypass_regNext_8_1_is_stationary_2;
  reg        [15:0]   io_in_c_bypass_regNext_8_2_data_2;
  reg                 io_in_c_bypass_regNext_8_2_is_stationary_2;
  reg        [15:0]   io_in_c_bypass_regNext_8_3_data_2;
  reg                 io_in_c_bypass_regNext_8_3_is_stationary_2;
  reg        [15:0]   io_in_c_bypass_regNext_9_0_data_2;
  reg                 io_in_c_bypass_regNext_9_0_is_stationary_2;
  reg        [15:0]   io_in_c_bypass_regNext_9_1_data_2;
  reg                 io_in_c_bypass_regNext_9_1_is_stationary_2;
  reg        [15:0]   io_in_c_bypass_regNext_9_2_data_2;
  reg                 io_in_c_bypass_regNext_9_2_is_stationary_2;
  reg        [15:0]   io_in_c_bypass_regNext_9_3_data_2;
  reg                 io_in_c_bypass_regNext_9_3_is_stationary_2;
  reg        [15:0]   io_in_c_bypass_regNext_10_0_data_2;
  reg                 io_in_c_bypass_regNext_10_0_is_stationary_2;
  reg        [15:0]   io_in_c_bypass_regNext_10_1_data_2;
  reg                 io_in_c_bypass_regNext_10_1_is_stationary_2;
  reg        [15:0]   io_in_c_bypass_regNext_10_2_data_2;
  reg                 io_in_c_bypass_regNext_10_2_is_stationary_2;
  reg        [15:0]   io_in_c_bypass_regNext_10_3_data_2;
  reg                 io_in_c_bypass_regNext_10_3_is_stationary_2;
  reg        [15:0]   io_in_c_bypass_regNext_11_0_data_2;
  reg                 io_in_c_bypass_regNext_11_0_is_stationary_2;
  reg        [15:0]   io_in_c_bypass_regNext_11_1_data_2;
  reg                 io_in_c_bypass_regNext_11_1_is_stationary_2;
  reg        [15:0]   io_in_c_bypass_regNext_11_2_data_2;
  reg                 io_in_c_bypass_regNext_11_2_is_stationary_2;
  reg        [15:0]   io_in_c_bypass_regNext_11_3_data_2;
  reg                 io_in_c_bypass_regNext_11_3_is_stationary_2;
  reg        [15:0]   io_in_c_bypass_regNext_12_0_data_2;
  reg                 io_in_c_bypass_regNext_12_0_is_stationary_2;
  reg        [15:0]   io_in_c_bypass_regNext_12_1_data_2;
  reg                 io_in_c_bypass_regNext_12_1_is_stationary_2;
  reg        [15:0]   io_in_c_bypass_regNext_12_2_data_2;
  reg                 io_in_c_bypass_regNext_12_2_is_stationary_2;
  reg        [15:0]   io_in_c_bypass_regNext_12_3_data_2;
  reg                 io_in_c_bypass_regNext_12_3_is_stationary_2;
  reg        [15:0]   io_in_c_bypass_regNext_13_0_data_2;
  reg                 io_in_c_bypass_regNext_13_0_is_stationary_2;
  reg        [15:0]   io_in_c_bypass_regNext_13_1_data_2;
  reg                 io_in_c_bypass_regNext_13_1_is_stationary_2;
  reg        [15:0]   io_in_c_bypass_regNext_13_2_data_2;
  reg                 io_in_c_bypass_regNext_13_2_is_stationary_2;
  reg        [15:0]   io_in_c_bypass_regNext_13_3_data_2;
  reg                 io_in_c_bypass_regNext_13_3_is_stationary_2;
  reg        [15:0]   io_in_c_bypass_regNext_14_0_data_2;
  reg                 io_in_c_bypass_regNext_14_0_is_stationary_2;
  reg        [15:0]   io_in_c_bypass_regNext_14_1_data_2;
  reg                 io_in_c_bypass_regNext_14_1_is_stationary_2;
  reg        [15:0]   io_in_c_bypass_regNext_14_2_data_2;
  reg                 io_in_c_bypass_regNext_14_2_is_stationary_2;
  reg        [15:0]   io_in_c_bypass_regNext_14_3_data_2;
  reg                 io_in_c_bypass_regNext_14_3_is_stationary_2;
  reg        [15:0]   io_in_c_bypass_regNext_15_0_data_2;
  reg                 io_in_c_bypass_regNext_15_0_is_stationary_2;
  reg        [15:0]   io_in_c_bypass_regNext_15_1_data_2;
  reg                 io_in_c_bypass_regNext_15_1_is_stationary_2;
  reg        [15:0]   io_in_c_bypass_regNext_15_2_data_2;
  reg                 io_in_c_bypass_regNext_15_2_is_stationary_2;
  reg        [15:0]   io_in_c_bypass_regNext_15_3_data_2;
  reg                 io_in_c_bypass_regNext_15_3_is_stationary_2;
  reg        [15:0]   io_in_c_bypass_regNext_16_0_data_2;
  reg                 io_in_c_bypass_regNext_16_0_is_stationary_2;
  reg        [15:0]   io_in_c_bypass_regNext_16_1_data_2;
  reg                 io_in_c_bypass_regNext_16_1_is_stationary_2;
  reg        [15:0]   io_in_c_bypass_regNext_16_2_data_2;
  reg                 io_in_c_bypass_regNext_16_2_is_stationary_2;
  reg        [15:0]   io_in_c_bypass_regNext_16_3_data_2;
  reg                 io_in_c_bypass_regNext_16_3_is_stationary_2;
  reg        [15:0]   io_in_c_bypass_regNext_17_0_data_2;
  reg                 io_in_c_bypass_regNext_17_0_is_stationary_2;
  reg        [15:0]   io_in_c_bypass_regNext_17_1_data_2;
  reg                 io_in_c_bypass_regNext_17_1_is_stationary_2;
  reg        [15:0]   io_in_c_bypass_regNext_17_2_data_2;
  reg                 io_in_c_bypass_regNext_17_2_is_stationary_2;
  reg        [15:0]   io_in_c_bypass_regNext_17_3_data_2;
  reg                 io_in_c_bypass_regNext_17_3_is_stationary_2;
  reg        [15:0]   io_in_c_bypass_regNext_18_0_data_2;
  reg                 io_in_c_bypass_regNext_18_0_is_stationary_2;
  reg        [15:0]   io_in_c_bypass_regNext_18_1_data_2;
  reg                 io_in_c_bypass_regNext_18_1_is_stationary_2;
  reg        [15:0]   io_in_c_bypass_regNext_18_2_data_2;
  reg                 io_in_c_bypass_regNext_18_2_is_stationary_2;
  reg        [15:0]   io_in_c_bypass_regNext_18_3_data_2;
  reg                 io_in_c_bypass_regNext_18_3_is_stationary_2;
  reg        [15:0]   io_in_c_bypass_regNext_19_0_data_2;
  reg                 io_in_c_bypass_regNext_19_0_is_stationary_2;
  reg        [15:0]   io_in_c_bypass_regNext_19_1_data_2;
  reg                 io_in_c_bypass_regNext_19_1_is_stationary_2;
  reg        [15:0]   io_in_c_bypass_regNext_19_2_data_2;
  reg                 io_in_c_bypass_regNext_19_2_is_stationary_2;
  reg        [15:0]   io_in_c_bypass_regNext_19_3_data_2;
  reg                 io_in_c_bypass_regNext_19_3_is_stationary_2;
  reg        [15:0]   io_in_c_bypass_regNext_20_0_data_2;
  reg                 io_in_c_bypass_regNext_20_0_is_stationary_2;
  reg        [15:0]   io_in_c_bypass_regNext_20_1_data_2;
  reg                 io_in_c_bypass_regNext_20_1_is_stationary_2;
  reg        [15:0]   io_in_c_bypass_regNext_20_2_data_2;
  reg                 io_in_c_bypass_regNext_20_2_is_stationary_2;
  reg        [15:0]   io_in_c_bypass_regNext_20_3_data_2;
  reg                 io_in_c_bypass_regNext_20_3_is_stationary_2;
  reg        [15:0]   io_in_c_bypass_regNext_21_0_data_2;
  reg                 io_in_c_bypass_regNext_21_0_is_stationary_2;
  reg        [15:0]   io_in_c_bypass_regNext_21_1_data_2;
  reg                 io_in_c_bypass_regNext_21_1_is_stationary_2;
  reg        [15:0]   io_in_c_bypass_regNext_21_2_data_2;
  reg                 io_in_c_bypass_regNext_21_2_is_stationary_2;
  reg        [15:0]   io_in_c_bypass_regNext_21_3_data_2;
  reg                 io_in_c_bypass_regNext_21_3_is_stationary_2;
  reg        [15:0]   io_in_c_bypass_regNext_22_0_data_2;
  reg                 io_in_c_bypass_regNext_22_0_is_stationary_2;
  reg        [15:0]   io_in_c_bypass_regNext_22_1_data_2;
  reg                 io_in_c_bypass_regNext_22_1_is_stationary_2;
  reg        [15:0]   io_in_c_bypass_regNext_22_2_data_2;
  reg                 io_in_c_bypass_regNext_22_2_is_stationary_2;
  reg        [15:0]   io_in_c_bypass_regNext_22_3_data_2;
  reg                 io_in_c_bypass_regNext_22_3_is_stationary_2;
  reg        [15:0]   io_in_c_bypass_regNext_23_0_data_2;
  reg                 io_in_c_bypass_regNext_23_0_is_stationary_2;
  reg        [15:0]   io_in_c_bypass_regNext_23_1_data_2;
  reg                 io_in_c_bypass_regNext_23_1_is_stationary_2;
  reg        [15:0]   io_in_c_bypass_regNext_23_2_data_2;
  reg                 io_in_c_bypass_regNext_23_2_is_stationary_2;
  reg        [15:0]   io_in_c_bypass_regNext_23_3_data_2;
  reg                 io_in_c_bypass_regNext_23_3_is_stationary_2;
  reg        [15:0]   io_in_c_bypass_regNext_24_0_data_2;
  reg                 io_in_c_bypass_regNext_24_0_is_stationary_2;
  reg        [15:0]   io_in_c_bypass_regNext_24_1_data_2;
  reg                 io_in_c_bypass_regNext_24_1_is_stationary_2;
  reg        [15:0]   io_in_c_bypass_regNext_24_2_data_2;
  reg                 io_in_c_bypass_regNext_24_2_is_stationary_2;
  reg        [15:0]   io_in_c_bypass_regNext_24_3_data_2;
  reg                 io_in_c_bypass_regNext_24_3_is_stationary_2;
  reg        [15:0]   io_in_c_bypass_regNext_25_0_data_2;
  reg                 io_in_c_bypass_regNext_25_0_is_stationary_2;
  reg        [15:0]   io_in_c_bypass_regNext_25_1_data_2;
  reg                 io_in_c_bypass_regNext_25_1_is_stationary_2;
  reg        [15:0]   io_in_c_bypass_regNext_25_2_data_2;
  reg                 io_in_c_bypass_regNext_25_2_is_stationary_2;
  reg        [15:0]   io_in_c_bypass_regNext_25_3_data_2;
  reg                 io_in_c_bypass_regNext_25_3_is_stationary_2;
  reg        [15:0]   io_in_c_bypass_regNext_26_0_data_2;
  reg                 io_in_c_bypass_regNext_26_0_is_stationary_2;
  reg        [15:0]   io_in_c_bypass_regNext_26_1_data_2;
  reg                 io_in_c_bypass_regNext_26_1_is_stationary_2;
  reg        [15:0]   io_in_c_bypass_regNext_26_2_data_2;
  reg                 io_in_c_bypass_regNext_26_2_is_stationary_2;
  reg        [15:0]   io_in_c_bypass_regNext_26_3_data_2;
  reg                 io_in_c_bypass_regNext_26_3_is_stationary_2;
  reg        [15:0]   io_in_c_bypass_regNext_27_0_data_2;
  reg                 io_in_c_bypass_regNext_27_0_is_stationary_2;
  reg        [15:0]   io_in_c_bypass_regNext_27_1_data_2;
  reg                 io_in_c_bypass_regNext_27_1_is_stationary_2;
  reg        [15:0]   io_in_c_bypass_regNext_27_2_data_2;
  reg                 io_in_c_bypass_regNext_27_2_is_stationary_2;
  reg        [15:0]   io_in_c_bypass_regNext_27_3_data_2;
  reg                 io_in_c_bypass_regNext_27_3_is_stationary_2;
  reg        [15:0]   io_in_c_bypass_regNext_28_0_data_2;
  reg                 io_in_c_bypass_regNext_28_0_is_stationary_2;
  reg        [15:0]   io_in_c_bypass_regNext_28_1_data_2;
  reg                 io_in_c_bypass_regNext_28_1_is_stationary_2;
  reg        [15:0]   io_in_c_bypass_regNext_28_2_data_2;
  reg                 io_in_c_bypass_regNext_28_2_is_stationary_2;
  reg        [15:0]   io_in_c_bypass_regNext_28_3_data_2;
  reg                 io_in_c_bypass_regNext_28_3_is_stationary_2;
  reg        [15:0]   io_in_c_bypass_regNext_29_0_data_2;
  reg                 io_in_c_bypass_regNext_29_0_is_stationary_2;
  reg        [15:0]   io_in_c_bypass_regNext_29_1_data_2;
  reg                 io_in_c_bypass_regNext_29_1_is_stationary_2;
  reg        [15:0]   io_in_c_bypass_regNext_29_2_data_2;
  reg                 io_in_c_bypass_regNext_29_2_is_stationary_2;
  reg        [15:0]   io_in_c_bypass_regNext_29_3_data_2;
  reg                 io_in_c_bypass_regNext_29_3_is_stationary_2;
  reg        [15:0]   io_in_c_bypass_regNext_30_0_data_2;
  reg                 io_in_c_bypass_regNext_30_0_is_stationary_2;
  reg        [15:0]   io_in_c_bypass_regNext_30_1_data_2;
  reg                 io_in_c_bypass_regNext_30_1_is_stationary_2;
  reg        [15:0]   io_in_c_bypass_regNext_30_2_data_2;
  reg                 io_in_c_bypass_regNext_30_2_is_stationary_2;
  reg        [15:0]   io_in_c_bypass_regNext_30_3_data_2;
  reg                 io_in_c_bypass_regNext_30_3_is_stationary_2;
  reg        [15:0]   io_in_c_bypass_regNext_31_0_data_2;
  reg                 io_in_c_bypass_regNext_31_0_is_stationary_2;
  reg        [15:0]   io_in_c_bypass_regNext_31_1_data_2;
  reg                 io_in_c_bypass_regNext_31_1_is_stationary_2;
  reg        [15:0]   io_in_c_bypass_regNext_31_2_data_2;
  reg                 io_in_c_bypass_regNext_31_2_is_stationary_2;
  reg        [15:0]   io_in_c_bypass_regNext_31_3_data_2;
  reg                 io_in_c_bypass_regNext_31_3_is_stationary_2;
  reg        [15:0]   io_in_c_bypass_regNext_0_0_data_3;
  reg                 io_in_c_bypass_regNext_0_0_is_stationary_3;
  reg        [15:0]   io_in_c_bypass_regNext_0_1_data_3;
  reg                 io_in_c_bypass_regNext_0_1_is_stationary_3;
  reg        [15:0]   io_in_c_bypass_regNext_0_2_data_3;
  reg                 io_in_c_bypass_regNext_0_2_is_stationary_3;
  reg        [15:0]   io_in_c_bypass_regNext_0_3_data_3;
  reg                 io_in_c_bypass_regNext_0_3_is_stationary_3;
  reg        [15:0]   io_in_c_bypass_regNext_1_0_data_3;
  reg                 io_in_c_bypass_regNext_1_0_is_stationary_3;
  reg        [15:0]   io_in_c_bypass_regNext_1_1_data_3;
  reg                 io_in_c_bypass_regNext_1_1_is_stationary_3;
  reg        [15:0]   io_in_c_bypass_regNext_1_2_data_3;
  reg                 io_in_c_bypass_regNext_1_2_is_stationary_3;
  reg        [15:0]   io_in_c_bypass_regNext_1_3_data_3;
  reg                 io_in_c_bypass_regNext_1_3_is_stationary_3;
  reg        [15:0]   io_in_c_bypass_regNext_2_0_data_3;
  reg                 io_in_c_bypass_regNext_2_0_is_stationary_3;
  reg        [15:0]   io_in_c_bypass_regNext_2_1_data_3;
  reg                 io_in_c_bypass_regNext_2_1_is_stationary_3;
  reg        [15:0]   io_in_c_bypass_regNext_2_2_data_3;
  reg                 io_in_c_bypass_regNext_2_2_is_stationary_3;
  reg        [15:0]   io_in_c_bypass_regNext_2_3_data_3;
  reg                 io_in_c_bypass_regNext_2_3_is_stationary_3;
  reg        [15:0]   io_in_c_bypass_regNext_3_0_data_3;
  reg                 io_in_c_bypass_regNext_3_0_is_stationary_3;
  reg        [15:0]   io_in_c_bypass_regNext_3_1_data_3;
  reg                 io_in_c_bypass_regNext_3_1_is_stationary_3;
  reg        [15:0]   io_in_c_bypass_regNext_3_2_data_3;
  reg                 io_in_c_bypass_regNext_3_2_is_stationary_3;
  reg        [15:0]   io_in_c_bypass_regNext_3_3_data_3;
  reg                 io_in_c_bypass_regNext_3_3_is_stationary_3;
  reg        [15:0]   io_in_c_bypass_regNext_4_0_data_3;
  reg                 io_in_c_bypass_regNext_4_0_is_stationary_3;
  reg        [15:0]   io_in_c_bypass_regNext_4_1_data_3;
  reg                 io_in_c_bypass_regNext_4_1_is_stationary_3;
  reg        [15:0]   io_in_c_bypass_regNext_4_2_data_3;
  reg                 io_in_c_bypass_regNext_4_2_is_stationary_3;
  reg        [15:0]   io_in_c_bypass_regNext_4_3_data_3;
  reg                 io_in_c_bypass_regNext_4_3_is_stationary_3;
  reg        [15:0]   io_in_c_bypass_regNext_5_0_data_3;
  reg                 io_in_c_bypass_regNext_5_0_is_stationary_3;
  reg        [15:0]   io_in_c_bypass_regNext_5_1_data_3;
  reg                 io_in_c_bypass_regNext_5_1_is_stationary_3;
  reg        [15:0]   io_in_c_bypass_regNext_5_2_data_3;
  reg                 io_in_c_bypass_regNext_5_2_is_stationary_3;
  reg        [15:0]   io_in_c_bypass_regNext_5_3_data_3;
  reg                 io_in_c_bypass_regNext_5_3_is_stationary_3;
  reg        [15:0]   io_in_c_bypass_regNext_6_0_data_3;
  reg                 io_in_c_bypass_regNext_6_0_is_stationary_3;
  reg        [15:0]   io_in_c_bypass_regNext_6_1_data_3;
  reg                 io_in_c_bypass_regNext_6_1_is_stationary_3;
  reg        [15:0]   io_in_c_bypass_regNext_6_2_data_3;
  reg                 io_in_c_bypass_regNext_6_2_is_stationary_3;
  reg        [15:0]   io_in_c_bypass_regNext_6_3_data_3;
  reg                 io_in_c_bypass_regNext_6_3_is_stationary_3;
  reg        [15:0]   io_in_c_bypass_regNext_7_0_data_3;
  reg                 io_in_c_bypass_regNext_7_0_is_stationary_3;
  reg        [15:0]   io_in_c_bypass_regNext_7_1_data_3;
  reg                 io_in_c_bypass_regNext_7_1_is_stationary_3;
  reg        [15:0]   io_in_c_bypass_regNext_7_2_data_3;
  reg                 io_in_c_bypass_regNext_7_2_is_stationary_3;
  reg        [15:0]   io_in_c_bypass_regNext_7_3_data_3;
  reg                 io_in_c_bypass_regNext_7_3_is_stationary_3;
  reg        [15:0]   io_in_c_bypass_regNext_8_0_data_3;
  reg                 io_in_c_bypass_regNext_8_0_is_stationary_3;
  reg        [15:0]   io_in_c_bypass_regNext_8_1_data_3;
  reg                 io_in_c_bypass_regNext_8_1_is_stationary_3;
  reg        [15:0]   io_in_c_bypass_regNext_8_2_data_3;
  reg                 io_in_c_bypass_regNext_8_2_is_stationary_3;
  reg        [15:0]   io_in_c_bypass_regNext_8_3_data_3;
  reg                 io_in_c_bypass_regNext_8_3_is_stationary_3;
  reg        [15:0]   io_in_c_bypass_regNext_9_0_data_3;
  reg                 io_in_c_bypass_regNext_9_0_is_stationary_3;
  reg        [15:0]   io_in_c_bypass_regNext_9_1_data_3;
  reg                 io_in_c_bypass_regNext_9_1_is_stationary_3;
  reg        [15:0]   io_in_c_bypass_regNext_9_2_data_3;
  reg                 io_in_c_bypass_regNext_9_2_is_stationary_3;
  reg        [15:0]   io_in_c_bypass_regNext_9_3_data_3;
  reg                 io_in_c_bypass_regNext_9_3_is_stationary_3;
  reg        [15:0]   io_in_c_bypass_regNext_10_0_data_3;
  reg                 io_in_c_bypass_regNext_10_0_is_stationary_3;
  reg        [15:0]   io_in_c_bypass_regNext_10_1_data_3;
  reg                 io_in_c_bypass_regNext_10_1_is_stationary_3;
  reg        [15:0]   io_in_c_bypass_regNext_10_2_data_3;
  reg                 io_in_c_bypass_regNext_10_2_is_stationary_3;
  reg        [15:0]   io_in_c_bypass_regNext_10_3_data_3;
  reg                 io_in_c_bypass_regNext_10_3_is_stationary_3;
  reg        [15:0]   io_in_c_bypass_regNext_11_0_data_3;
  reg                 io_in_c_bypass_regNext_11_0_is_stationary_3;
  reg        [15:0]   io_in_c_bypass_regNext_11_1_data_3;
  reg                 io_in_c_bypass_regNext_11_1_is_stationary_3;
  reg        [15:0]   io_in_c_bypass_regNext_11_2_data_3;
  reg                 io_in_c_bypass_regNext_11_2_is_stationary_3;
  reg        [15:0]   io_in_c_bypass_regNext_11_3_data_3;
  reg                 io_in_c_bypass_regNext_11_3_is_stationary_3;
  reg        [15:0]   io_in_c_bypass_regNext_12_0_data_3;
  reg                 io_in_c_bypass_regNext_12_0_is_stationary_3;
  reg        [15:0]   io_in_c_bypass_regNext_12_1_data_3;
  reg                 io_in_c_bypass_regNext_12_1_is_stationary_3;
  reg        [15:0]   io_in_c_bypass_regNext_12_2_data_3;
  reg                 io_in_c_bypass_regNext_12_2_is_stationary_3;
  reg        [15:0]   io_in_c_bypass_regNext_12_3_data_3;
  reg                 io_in_c_bypass_regNext_12_3_is_stationary_3;
  reg        [15:0]   io_in_c_bypass_regNext_13_0_data_3;
  reg                 io_in_c_bypass_regNext_13_0_is_stationary_3;
  reg        [15:0]   io_in_c_bypass_regNext_13_1_data_3;
  reg                 io_in_c_bypass_regNext_13_1_is_stationary_3;
  reg        [15:0]   io_in_c_bypass_regNext_13_2_data_3;
  reg                 io_in_c_bypass_regNext_13_2_is_stationary_3;
  reg        [15:0]   io_in_c_bypass_regNext_13_3_data_3;
  reg                 io_in_c_bypass_regNext_13_3_is_stationary_3;
  reg        [15:0]   io_in_c_bypass_regNext_14_0_data_3;
  reg                 io_in_c_bypass_regNext_14_0_is_stationary_3;
  reg        [15:0]   io_in_c_bypass_regNext_14_1_data_3;
  reg                 io_in_c_bypass_regNext_14_1_is_stationary_3;
  reg        [15:0]   io_in_c_bypass_regNext_14_2_data_3;
  reg                 io_in_c_bypass_regNext_14_2_is_stationary_3;
  reg        [15:0]   io_in_c_bypass_regNext_14_3_data_3;
  reg                 io_in_c_bypass_regNext_14_3_is_stationary_3;
  reg        [15:0]   io_in_c_bypass_regNext_15_0_data_3;
  reg                 io_in_c_bypass_regNext_15_0_is_stationary_3;
  reg        [15:0]   io_in_c_bypass_regNext_15_1_data_3;
  reg                 io_in_c_bypass_regNext_15_1_is_stationary_3;
  reg        [15:0]   io_in_c_bypass_regNext_15_2_data_3;
  reg                 io_in_c_bypass_regNext_15_2_is_stationary_3;
  reg        [15:0]   io_in_c_bypass_regNext_15_3_data_3;
  reg                 io_in_c_bypass_regNext_15_3_is_stationary_3;
  reg        [15:0]   io_in_c_bypass_regNext_16_0_data_3;
  reg                 io_in_c_bypass_regNext_16_0_is_stationary_3;
  reg        [15:0]   io_in_c_bypass_regNext_16_1_data_3;
  reg                 io_in_c_bypass_regNext_16_1_is_stationary_3;
  reg        [15:0]   io_in_c_bypass_regNext_16_2_data_3;
  reg                 io_in_c_bypass_regNext_16_2_is_stationary_3;
  reg        [15:0]   io_in_c_bypass_regNext_16_3_data_3;
  reg                 io_in_c_bypass_regNext_16_3_is_stationary_3;
  reg        [15:0]   io_in_c_bypass_regNext_17_0_data_3;
  reg                 io_in_c_bypass_regNext_17_0_is_stationary_3;
  reg        [15:0]   io_in_c_bypass_regNext_17_1_data_3;
  reg                 io_in_c_bypass_regNext_17_1_is_stationary_3;
  reg        [15:0]   io_in_c_bypass_regNext_17_2_data_3;
  reg                 io_in_c_bypass_regNext_17_2_is_stationary_3;
  reg        [15:0]   io_in_c_bypass_regNext_17_3_data_3;
  reg                 io_in_c_bypass_regNext_17_3_is_stationary_3;
  reg        [15:0]   io_in_c_bypass_regNext_18_0_data_3;
  reg                 io_in_c_bypass_regNext_18_0_is_stationary_3;
  reg        [15:0]   io_in_c_bypass_regNext_18_1_data_3;
  reg                 io_in_c_bypass_regNext_18_1_is_stationary_3;
  reg        [15:0]   io_in_c_bypass_regNext_18_2_data_3;
  reg                 io_in_c_bypass_regNext_18_2_is_stationary_3;
  reg        [15:0]   io_in_c_bypass_regNext_18_3_data_3;
  reg                 io_in_c_bypass_regNext_18_3_is_stationary_3;
  reg        [15:0]   io_in_c_bypass_regNext_19_0_data_3;
  reg                 io_in_c_bypass_regNext_19_0_is_stationary_3;
  reg        [15:0]   io_in_c_bypass_regNext_19_1_data_3;
  reg                 io_in_c_bypass_regNext_19_1_is_stationary_3;
  reg        [15:0]   io_in_c_bypass_regNext_19_2_data_3;
  reg                 io_in_c_bypass_regNext_19_2_is_stationary_3;
  reg        [15:0]   io_in_c_bypass_regNext_19_3_data_3;
  reg                 io_in_c_bypass_regNext_19_3_is_stationary_3;
  reg        [15:0]   io_in_c_bypass_regNext_20_0_data_3;
  reg                 io_in_c_bypass_regNext_20_0_is_stationary_3;
  reg        [15:0]   io_in_c_bypass_regNext_20_1_data_3;
  reg                 io_in_c_bypass_regNext_20_1_is_stationary_3;
  reg        [15:0]   io_in_c_bypass_regNext_20_2_data_3;
  reg                 io_in_c_bypass_regNext_20_2_is_stationary_3;
  reg        [15:0]   io_in_c_bypass_regNext_20_3_data_3;
  reg                 io_in_c_bypass_regNext_20_3_is_stationary_3;
  reg        [15:0]   io_in_c_bypass_regNext_21_0_data_3;
  reg                 io_in_c_bypass_regNext_21_0_is_stationary_3;
  reg        [15:0]   io_in_c_bypass_regNext_21_1_data_3;
  reg                 io_in_c_bypass_regNext_21_1_is_stationary_3;
  reg        [15:0]   io_in_c_bypass_regNext_21_2_data_3;
  reg                 io_in_c_bypass_regNext_21_2_is_stationary_3;
  reg        [15:0]   io_in_c_bypass_regNext_21_3_data_3;
  reg                 io_in_c_bypass_regNext_21_3_is_stationary_3;
  reg        [15:0]   io_in_c_bypass_regNext_22_0_data_3;
  reg                 io_in_c_bypass_regNext_22_0_is_stationary_3;
  reg        [15:0]   io_in_c_bypass_regNext_22_1_data_3;
  reg                 io_in_c_bypass_regNext_22_1_is_stationary_3;
  reg        [15:0]   io_in_c_bypass_regNext_22_2_data_3;
  reg                 io_in_c_bypass_regNext_22_2_is_stationary_3;
  reg        [15:0]   io_in_c_bypass_regNext_22_3_data_3;
  reg                 io_in_c_bypass_regNext_22_3_is_stationary_3;
  reg        [15:0]   io_in_c_bypass_regNext_23_0_data_3;
  reg                 io_in_c_bypass_regNext_23_0_is_stationary_3;
  reg        [15:0]   io_in_c_bypass_regNext_23_1_data_3;
  reg                 io_in_c_bypass_regNext_23_1_is_stationary_3;
  reg        [15:0]   io_in_c_bypass_regNext_23_2_data_3;
  reg                 io_in_c_bypass_regNext_23_2_is_stationary_3;
  reg        [15:0]   io_in_c_bypass_regNext_23_3_data_3;
  reg                 io_in_c_bypass_regNext_23_3_is_stationary_3;
  reg        [15:0]   io_in_c_bypass_regNext_24_0_data_3;
  reg                 io_in_c_bypass_regNext_24_0_is_stationary_3;
  reg        [15:0]   io_in_c_bypass_regNext_24_1_data_3;
  reg                 io_in_c_bypass_regNext_24_1_is_stationary_3;
  reg        [15:0]   io_in_c_bypass_regNext_24_2_data_3;
  reg                 io_in_c_bypass_regNext_24_2_is_stationary_3;
  reg        [15:0]   io_in_c_bypass_regNext_24_3_data_3;
  reg                 io_in_c_bypass_regNext_24_3_is_stationary_3;
  reg        [15:0]   io_in_c_bypass_regNext_25_0_data_3;
  reg                 io_in_c_bypass_regNext_25_0_is_stationary_3;
  reg        [15:0]   io_in_c_bypass_regNext_25_1_data_3;
  reg                 io_in_c_bypass_regNext_25_1_is_stationary_3;
  reg        [15:0]   io_in_c_bypass_regNext_25_2_data_3;
  reg                 io_in_c_bypass_regNext_25_2_is_stationary_3;
  reg        [15:0]   io_in_c_bypass_regNext_25_3_data_3;
  reg                 io_in_c_bypass_regNext_25_3_is_stationary_3;
  reg        [15:0]   io_in_c_bypass_regNext_26_0_data_3;
  reg                 io_in_c_bypass_regNext_26_0_is_stationary_3;
  reg        [15:0]   io_in_c_bypass_regNext_26_1_data_3;
  reg                 io_in_c_bypass_regNext_26_1_is_stationary_3;
  reg        [15:0]   io_in_c_bypass_regNext_26_2_data_3;
  reg                 io_in_c_bypass_regNext_26_2_is_stationary_3;
  reg        [15:0]   io_in_c_bypass_regNext_26_3_data_3;
  reg                 io_in_c_bypass_regNext_26_3_is_stationary_3;
  reg        [15:0]   io_in_c_bypass_regNext_27_0_data_3;
  reg                 io_in_c_bypass_regNext_27_0_is_stationary_3;
  reg        [15:0]   io_in_c_bypass_regNext_27_1_data_3;
  reg                 io_in_c_bypass_regNext_27_1_is_stationary_3;
  reg        [15:0]   io_in_c_bypass_regNext_27_2_data_3;
  reg                 io_in_c_bypass_regNext_27_2_is_stationary_3;
  reg        [15:0]   io_in_c_bypass_regNext_27_3_data_3;
  reg                 io_in_c_bypass_regNext_27_3_is_stationary_3;
  reg        [15:0]   io_in_c_bypass_regNext_28_0_data_3;
  reg                 io_in_c_bypass_regNext_28_0_is_stationary_3;
  reg        [15:0]   io_in_c_bypass_regNext_28_1_data_3;
  reg                 io_in_c_bypass_regNext_28_1_is_stationary_3;
  reg        [15:0]   io_in_c_bypass_regNext_28_2_data_3;
  reg                 io_in_c_bypass_regNext_28_2_is_stationary_3;
  reg        [15:0]   io_in_c_bypass_regNext_28_3_data_3;
  reg                 io_in_c_bypass_regNext_28_3_is_stationary_3;
  reg        [15:0]   io_in_c_bypass_regNext_29_0_data_3;
  reg                 io_in_c_bypass_regNext_29_0_is_stationary_3;
  reg        [15:0]   io_in_c_bypass_regNext_29_1_data_3;
  reg                 io_in_c_bypass_regNext_29_1_is_stationary_3;
  reg        [15:0]   io_in_c_bypass_regNext_29_2_data_3;
  reg                 io_in_c_bypass_regNext_29_2_is_stationary_3;
  reg        [15:0]   io_in_c_bypass_regNext_29_3_data_3;
  reg                 io_in_c_bypass_regNext_29_3_is_stationary_3;
  reg        [15:0]   io_in_c_bypass_regNext_30_0_data_3;
  reg                 io_in_c_bypass_regNext_30_0_is_stationary_3;
  reg        [15:0]   io_in_c_bypass_regNext_30_1_data_3;
  reg                 io_in_c_bypass_regNext_30_1_is_stationary_3;
  reg        [15:0]   io_in_c_bypass_regNext_30_2_data_3;
  reg                 io_in_c_bypass_regNext_30_2_is_stationary_3;
  reg        [15:0]   io_in_c_bypass_regNext_30_3_data_3;
  reg                 io_in_c_bypass_regNext_30_3_is_stationary_3;
  reg        [15:0]   io_in_c_bypass_regNext_31_0_data_3;
  reg                 io_in_c_bypass_regNext_31_0_is_stationary_3;
  reg        [15:0]   io_in_c_bypass_regNext_31_1_data_3;
  reg                 io_in_c_bypass_regNext_31_1_is_stationary_3;
  reg        [15:0]   io_in_c_bypass_regNext_31_2_data_3;
  reg                 io_in_c_bypass_regNext_31_2_is_stationary_3;
  reg        [15:0]   io_in_c_bypass_regNext_31_3_data_3;
  reg                 io_in_c_bypass_regNext_31_3_is_stationary_3;
  reg        [15:0]   io_in_c_bypass_regNext_0_0_data_4;
  reg                 io_in_c_bypass_regNext_0_0_is_stationary_4;
  reg        [15:0]   io_in_c_bypass_regNext_0_1_data_4;
  reg                 io_in_c_bypass_regNext_0_1_is_stationary_4;
  reg        [15:0]   io_in_c_bypass_regNext_0_2_data_4;
  reg                 io_in_c_bypass_regNext_0_2_is_stationary_4;
  reg        [15:0]   io_in_c_bypass_regNext_0_3_data_4;
  reg                 io_in_c_bypass_regNext_0_3_is_stationary_4;
  reg        [15:0]   io_in_c_bypass_regNext_1_0_data_4;
  reg                 io_in_c_bypass_regNext_1_0_is_stationary_4;
  reg        [15:0]   io_in_c_bypass_regNext_1_1_data_4;
  reg                 io_in_c_bypass_regNext_1_1_is_stationary_4;
  reg        [15:0]   io_in_c_bypass_regNext_1_2_data_4;
  reg                 io_in_c_bypass_regNext_1_2_is_stationary_4;
  reg        [15:0]   io_in_c_bypass_regNext_1_3_data_4;
  reg                 io_in_c_bypass_regNext_1_3_is_stationary_4;
  reg        [15:0]   io_in_c_bypass_regNext_2_0_data_4;
  reg                 io_in_c_bypass_regNext_2_0_is_stationary_4;
  reg        [15:0]   io_in_c_bypass_regNext_2_1_data_4;
  reg                 io_in_c_bypass_regNext_2_1_is_stationary_4;
  reg        [15:0]   io_in_c_bypass_regNext_2_2_data_4;
  reg                 io_in_c_bypass_regNext_2_2_is_stationary_4;
  reg        [15:0]   io_in_c_bypass_regNext_2_3_data_4;
  reg                 io_in_c_bypass_regNext_2_3_is_stationary_4;
  reg        [15:0]   io_in_c_bypass_regNext_3_0_data_4;
  reg                 io_in_c_bypass_regNext_3_0_is_stationary_4;
  reg        [15:0]   io_in_c_bypass_regNext_3_1_data_4;
  reg                 io_in_c_bypass_regNext_3_1_is_stationary_4;
  reg        [15:0]   io_in_c_bypass_regNext_3_2_data_4;
  reg                 io_in_c_bypass_regNext_3_2_is_stationary_4;
  reg        [15:0]   io_in_c_bypass_regNext_3_3_data_4;
  reg                 io_in_c_bypass_regNext_3_3_is_stationary_4;
  reg        [15:0]   io_in_c_bypass_regNext_4_0_data_4;
  reg                 io_in_c_bypass_regNext_4_0_is_stationary_4;
  reg        [15:0]   io_in_c_bypass_regNext_4_1_data_4;
  reg                 io_in_c_bypass_regNext_4_1_is_stationary_4;
  reg        [15:0]   io_in_c_bypass_regNext_4_2_data_4;
  reg                 io_in_c_bypass_regNext_4_2_is_stationary_4;
  reg        [15:0]   io_in_c_bypass_regNext_4_3_data_4;
  reg                 io_in_c_bypass_regNext_4_3_is_stationary_4;
  reg        [15:0]   io_in_c_bypass_regNext_5_0_data_4;
  reg                 io_in_c_bypass_regNext_5_0_is_stationary_4;
  reg        [15:0]   io_in_c_bypass_regNext_5_1_data_4;
  reg                 io_in_c_bypass_regNext_5_1_is_stationary_4;
  reg        [15:0]   io_in_c_bypass_regNext_5_2_data_4;
  reg                 io_in_c_bypass_regNext_5_2_is_stationary_4;
  reg        [15:0]   io_in_c_bypass_regNext_5_3_data_4;
  reg                 io_in_c_bypass_regNext_5_3_is_stationary_4;
  reg        [15:0]   io_in_c_bypass_regNext_6_0_data_4;
  reg                 io_in_c_bypass_regNext_6_0_is_stationary_4;
  reg        [15:0]   io_in_c_bypass_regNext_6_1_data_4;
  reg                 io_in_c_bypass_regNext_6_1_is_stationary_4;
  reg        [15:0]   io_in_c_bypass_regNext_6_2_data_4;
  reg                 io_in_c_bypass_regNext_6_2_is_stationary_4;
  reg        [15:0]   io_in_c_bypass_regNext_6_3_data_4;
  reg                 io_in_c_bypass_regNext_6_3_is_stationary_4;
  reg        [15:0]   io_in_c_bypass_regNext_7_0_data_4;
  reg                 io_in_c_bypass_regNext_7_0_is_stationary_4;
  reg        [15:0]   io_in_c_bypass_regNext_7_1_data_4;
  reg                 io_in_c_bypass_regNext_7_1_is_stationary_4;
  reg        [15:0]   io_in_c_bypass_regNext_7_2_data_4;
  reg                 io_in_c_bypass_regNext_7_2_is_stationary_4;
  reg        [15:0]   io_in_c_bypass_regNext_7_3_data_4;
  reg                 io_in_c_bypass_regNext_7_3_is_stationary_4;
  reg        [15:0]   io_in_c_bypass_regNext_8_0_data_4;
  reg                 io_in_c_bypass_regNext_8_0_is_stationary_4;
  reg        [15:0]   io_in_c_bypass_regNext_8_1_data_4;
  reg                 io_in_c_bypass_regNext_8_1_is_stationary_4;
  reg        [15:0]   io_in_c_bypass_regNext_8_2_data_4;
  reg                 io_in_c_bypass_regNext_8_2_is_stationary_4;
  reg        [15:0]   io_in_c_bypass_regNext_8_3_data_4;
  reg                 io_in_c_bypass_regNext_8_3_is_stationary_4;
  reg        [15:0]   io_in_c_bypass_regNext_9_0_data_4;
  reg                 io_in_c_bypass_regNext_9_0_is_stationary_4;
  reg        [15:0]   io_in_c_bypass_regNext_9_1_data_4;
  reg                 io_in_c_bypass_regNext_9_1_is_stationary_4;
  reg        [15:0]   io_in_c_bypass_regNext_9_2_data_4;
  reg                 io_in_c_bypass_regNext_9_2_is_stationary_4;
  reg        [15:0]   io_in_c_bypass_regNext_9_3_data_4;
  reg                 io_in_c_bypass_regNext_9_3_is_stationary_4;
  reg        [15:0]   io_in_c_bypass_regNext_10_0_data_4;
  reg                 io_in_c_bypass_regNext_10_0_is_stationary_4;
  reg        [15:0]   io_in_c_bypass_regNext_10_1_data_4;
  reg                 io_in_c_bypass_regNext_10_1_is_stationary_4;
  reg        [15:0]   io_in_c_bypass_regNext_10_2_data_4;
  reg                 io_in_c_bypass_regNext_10_2_is_stationary_4;
  reg        [15:0]   io_in_c_bypass_regNext_10_3_data_4;
  reg                 io_in_c_bypass_regNext_10_3_is_stationary_4;
  reg        [15:0]   io_in_c_bypass_regNext_11_0_data_4;
  reg                 io_in_c_bypass_regNext_11_0_is_stationary_4;
  reg        [15:0]   io_in_c_bypass_regNext_11_1_data_4;
  reg                 io_in_c_bypass_regNext_11_1_is_stationary_4;
  reg        [15:0]   io_in_c_bypass_regNext_11_2_data_4;
  reg                 io_in_c_bypass_regNext_11_2_is_stationary_4;
  reg        [15:0]   io_in_c_bypass_regNext_11_3_data_4;
  reg                 io_in_c_bypass_regNext_11_3_is_stationary_4;
  reg        [15:0]   io_in_c_bypass_regNext_12_0_data_4;
  reg                 io_in_c_bypass_regNext_12_0_is_stationary_4;
  reg        [15:0]   io_in_c_bypass_regNext_12_1_data_4;
  reg                 io_in_c_bypass_regNext_12_1_is_stationary_4;
  reg        [15:0]   io_in_c_bypass_regNext_12_2_data_4;
  reg                 io_in_c_bypass_regNext_12_2_is_stationary_4;
  reg        [15:0]   io_in_c_bypass_regNext_12_3_data_4;
  reg                 io_in_c_bypass_regNext_12_3_is_stationary_4;
  reg        [15:0]   io_in_c_bypass_regNext_13_0_data_4;
  reg                 io_in_c_bypass_regNext_13_0_is_stationary_4;
  reg        [15:0]   io_in_c_bypass_regNext_13_1_data_4;
  reg                 io_in_c_bypass_regNext_13_1_is_stationary_4;
  reg        [15:0]   io_in_c_bypass_regNext_13_2_data_4;
  reg                 io_in_c_bypass_regNext_13_2_is_stationary_4;
  reg        [15:0]   io_in_c_bypass_regNext_13_3_data_4;
  reg                 io_in_c_bypass_regNext_13_3_is_stationary_4;
  reg        [15:0]   io_in_c_bypass_regNext_14_0_data_4;
  reg                 io_in_c_bypass_regNext_14_0_is_stationary_4;
  reg        [15:0]   io_in_c_bypass_regNext_14_1_data_4;
  reg                 io_in_c_bypass_regNext_14_1_is_stationary_4;
  reg        [15:0]   io_in_c_bypass_regNext_14_2_data_4;
  reg                 io_in_c_bypass_regNext_14_2_is_stationary_4;
  reg        [15:0]   io_in_c_bypass_regNext_14_3_data_4;
  reg                 io_in_c_bypass_regNext_14_3_is_stationary_4;
  reg        [15:0]   io_in_c_bypass_regNext_15_0_data_4;
  reg                 io_in_c_bypass_regNext_15_0_is_stationary_4;
  reg        [15:0]   io_in_c_bypass_regNext_15_1_data_4;
  reg                 io_in_c_bypass_regNext_15_1_is_stationary_4;
  reg        [15:0]   io_in_c_bypass_regNext_15_2_data_4;
  reg                 io_in_c_bypass_regNext_15_2_is_stationary_4;
  reg        [15:0]   io_in_c_bypass_regNext_15_3_data_4;
  reg                 io_in_c_bypass_regNext_15_3_is_stationary_4;
  reg        [15:0]   io_in_c_bypass_regNext_16_0_data_4;
  reg                 io_in_c_bypass_regNext_16_0_is_stationary_4;
  reg        [15:0]   io_in_c_bypass_regNext_16_1_data_4;
  reg                 io_in_c_bypass_regNext_16_1_is_stationary_4;
  reg        [15:0]   io_in_c_bypass_regNext_16_2_data_4;
  reg                 io_in_c_bypass_regNext_16_2_is_stationary_4;
  reg        [15:0]   io_in_c_bypass_regNext_16_3_data_4;
  reg                 io_in_c_bypass_regNext_16_3_is_stationary_4;
  reg        [15:0]   io_in_c_bypass_regNext_17_0_data_4;
  reg                 io_in_c_bypass_regNext_17_0_is_stationary_4;
  reg        [15:0]   io_in_c_bypass_regNext_17_1_data_4;
  reg                 io_in_c_bypass_regNext_17_1_is_stationary_4;
  reg        [15:0]   io_in_c_bypass_regNext_17_2_data_4;
  reg                 io_in_c_bypass_regNext_17_2_is_stationary_4;
  reg        [15:0]   io_in_c_bypass_regNext_17_3_data_4;
  reg                 io_in_c_bypass_regNext_17_3_is_stationary_4;
  reg        [15:0]   io_in_c_bypass_regNext_18_0_data_4;
  reg                 io_in_c_bypass_regNext_18_0_is_stationary_4;
  reg        [15:0]   io_in_c_bypass_regNext_18_1_data_4;
  reg                 io_in_c_bypass_regNext_18_1_is_stationary_4;
  reg        [15:0]   io_in_c_bypass_regNext_18_2_data_4;
  reg                 io_in_c_bypass_regNext_18_2_is_stationary_4;
  reg        [15:0]   io_in_c_bypass_regNext_18_3_data_4;
  reg                 io_in_c_bypass_regNext_18_3_is_stationary_4;
  reg        [15:0]   io_in_c_bypass_regNext_19_0_data_4;
  reg                 io_in_c_bypass_regNext_19_0_is_stationary_4;
  reg        [15:0]   io_in_c_bypass_regNext_19_1_data_4;
  reg                 io_in_c_bypass_regNext_19_1_is_stationary_4;
  reg        [15:0]   io_in_c_bypass_regNext_19_2_data_4;
  reg                 io_in_c_bypass_regNext_19_2_is_stationary_4;
  reg        [15:0]   io_in_c_bypass_regNext_19_3_data_4;
  reg                 io_in_c_bypass_regNext_19_3_is_stationary_4;
  reg        [15:0]   io_in_c_bypass_regNext_20_0_data_4;
  reg                 io_in_c_bypass_regNext_20_0_is_stationary_4;
  reg        [15:0]   io_in_c_bypass_regNext_20_1_data_4;
  reg                 io_in_c_bypass_regNext_20_1_is_stationary_4;
  reg        [15:0]   io_in_c_bypass_regNext_20_2_data_4;
  reg                 io_in_c_bypass_regNext_20_2_is_stationary_4;
  reg        [15:0]   io_in_c_bypass_regNext_20_3_data_4;
  reg                 io_in_c_bypass_regNext_20_3_is_stationary_4;
  reg        [15:0]   io_in_c_bypass_regNext_21_0_data_4;
  reg                 io_in_c_bypass_regNext_21_0_is_stationary_4;
  reg        [15:0]   io_in_c_bypass_regNext_21_1_data_4;
  reg                 io_in_c_bypass_regNext_21_1_is_stationary_4;
  reg        [15:0]   io_in_c_bypass_regNext_21_2_data_4;
  reg                 io_in_c_bypass_regNext_21_2_is_stationary_4;
  reg        [15:0]   io_in_c_bypass_regNext_21_3_data_4;
  reg                 io_in_c_bypass_regNext_21_3_is_stationary_4;
  reg        [15:0]   io_in_c_bypass_regNext_22_0_data_4;
  reg                 io_in_c_bypass_regNext_22_0_is_stationary_4;
  reg        [15:0]   io_in_c_bypass_regNext_22_1_data_4;
  reg                 io_in_c_bypass_regNext_22_1_is_stationary_4;
  reg        [15:0]   io_in_c_bypass_regNext_22_2_data_4;
  reg                 io_in_c_bypass_regNext_22_2_is_stationary_4;
  reg        [15:0]   io_in_c_bypass_regNext_22_3_data_4;
  reg                 io_in_c_bypass_regNext_22_3_is_stationary_4;
  reg        [15:0]   io_in_c_bypass_regNext_23_0_data_4;
  reg                 io_in_c_bypass_regNext_23_0_is_stationary_4;
  reg        [15:0]   io_in_c_bypass_regNext_23_1_data_4;
  reg                 io_in_c_bypass_regNext_23_1_is_stationary_4;
  reg        [15:0]   io_in_c_bypass_regNext_23_2_data_4;
  reg                 io_in_c_bypass_regNext_23_2_is_stationary_4;
  reg        [15:0]   io_in_c_bypass_regNext_23_3_data_4;
  reg                 io_in_c_bypass_regNext_23_3_is_stationary_4;
  reg        [15:0]   io_in_c_bypass_regNext_24_0_data_4;
  reg                 io_in_c_bypass_regNext_24_0_is_stationary_4;
  reg        [15:0]   io_in_c_bypass_regNext_24_1_data_4;
  reg                 io_in_c_bypass_regNext_24_1_is_stationary_4;
  reg        [15:0]   io_in_c_bypass_regNext_24_2_data_4;
  reg                 io_in_c_bypass_regNext_24_2_is_stationary_4;
  reg        [15:0]   io_in_c_bypass_regNext_24_3_data_4;
  reg                 io_in_c_bypass_regNext_24_3_is_stationary_4;
  reg        [15:0]   io_in_c_bypass_regNext_25_0_data_4;
  reg                 io_in_c_bypass_regNext_25_0_is_stationary_4;
  reg        [15:0]   io_in_c_bypass_regNext_25_1_data_4;
  reg                 io_in_c_bypass_regNext_25_1_is_stationary_4;
  reg        [15:0]   io_in_c_bypass_regNext_25_2_data_4;
  reg                 io_in_c_bypass_regNext_25_2_is_stationary_4;
  reg        [15:0]   io_in_c_bypass_regNext_25_3_data_4;
  reg                 io_in_c_bypass_regNext_25_3_is_stationary_4;
  reg        [15:0]   io_in_c_bypass_regNext_26_0_data_4;
  reg                 io_in_c_bypass_regNext_26_0_is_stationary_4;
  reg        [15:0]   io_in_c_bypass_regNext_26_1_data_4;
  reg                 io_in_c_bypass_regNext_26_1_is_stationary_4;
  reg        [15:0]   io_in_c_bypass_regNext_26_2_data_4;
  reg                 io_in_c_bypass_regNext_26_2_is_stationary_4;
  reg        [15:0]   io_in_c_bypass_regNext_26_3_data_4;
  reg                 io_in_c_bypass_regNext_26_3_is_stationary_4;
  reg        [15:0]   io_in_c_bypass_regNext_27_0_data_4;
  reg                 io_in_c_bypass_regNext_27_0_is_stationary_4;
  reg        [15:0]   io_in_c_bypass_regNext_27_1_data_4;
  reg                 io_in_c_bypass_regNext_27_1_is_stationary_4;
  reg        [15:0]   io_in_c_bypass_regNext_27_2_data_4;
  reg                 io_in_c_bypass_regNext_27_2_is_stationary_4;
  reg        [15:0]   io_in_c_bypass_regNext_27_3_data_4;
  reg                 io_in_c_bypass_regNext_27_3_is_stationary_4;
  reg        [15:0]   io_in_c_bypass_regNext_28_0_data_4;
  reg                 io_in_c_bypass_regNext_28_0_is_stationary_4;
  reg        [15:0]   io_in_c_bypass_regNext_28_1_data_4;
  reg                 io_in_c_bypass_regNext_28_1_is_stationary_4;
  reg        [15:0]   io_in_c_bypass_regNext_28_2_data_4;
  reg                 io_in_c_bypass_regNext_28_2_is_stationary_4;
  reg        [15:0]   io_in_c_bypass_regNext_28_3_data_4;
  reg                 io_in_c_bypass_regNext_28_3_is_stationary_4;
  reg        [15:0]   io_in_c_bypass_regNext_29_0_data_4;
  reg                 io_in_c_bypass_regNext_29_0_is_stationary_4;
  reg        [15:0]   io_in_c_bypass_regNext_29_1_data_4;
  reg                 io_in_c_bypass_regNext_29_1_is_stationary_4;
  reg        [15:0]   io_in_c_bypass_regNext_29_2_data_4;
  reg                 io_in_c_bypass_regNext_29_2_is_stationary_4;
  reg        [15:0]   io_in_c_bypass_regNext_29_3_data_4;
  reg                 io_in_c_bypass_regNext_29_3_is_stationary_4;
  reg        [15:0]   io_in_c_bypass_regNext_30_0_data_4;
  reg                 io_in_c_bypass_regNext_30_0_is_stationary_4;
  reg        [15:0]   io_in_c_bypass_regNext_30_1_data_4;
  reg                 io_in_c_bypass_regNext_30_1_is_stationary_4;
  reg        [15:0]   io_in_c_bypass_regNext_30_2_data_4;
  reg                 io_in_c_bypass_regNext_30_2_is_stationary_4;
  reg        [15:0]   io_in_c_bypass_regNext_30_3_data_4;
  reg                 io_in_c_bypass_regNext_30_3_is_stationary_4;
  reg        [15:0]   io_in_c_bypass_regNext_31_0_data_4;
  reg                 io_in_c_bypass_regNext_31_0_is_stationary_4;
  reg        [15:0]   io_in_c_bypass_regNext_31_1_data_4;
  reg                 io_in_c_bypass_regNext_31_1_is_stationary_4;
  reg        [15:0]   io_in_c_bypass_regNext_31_2_data_4;
  reg                 io_in_c_bypass_regNext_31_2_is_stationary_4;
  reg        [15:0]   io_in_c_bypass_regNext_31_3_data_4;
  reg                 io_in_c_bypass_regNext_31_3_is_stationary_4;
  reg        [15:0]   io_in_c_bypass_regNext_0_0_data_5;
  reg                 io_in_c_bypass_regNext_0_0_is_stationary_5;
  reg        [15:0]   io_in_c_bypass_regNext_0_1_data_5;
  reg                 io_in_c_bypass_regNext_0_1_is_stationary_5;
  reg        [15:0]   io_in_c_bypass_regNext_0_2_data_5;
  reg                 io_in_c_bypass_regNext_0_2_is_stationary_5;
  reg        [15:0]   io_in_c_bypass_regNext_0_3_data_5;
  reg                 io_in_c_bypass_regNext_0_3_is_stationary_5;
  reg        [15:0]   io_in_c_bypass_regNext_1_0_data_5;
  reg                 io_in_c_bypass_regNext_1_0_is_stationary_5;
  reg        [15:0]   io_in_c_bypass_regNext_1_1_data_5;
  reg                 io_in_c_bypass_regNext_1_1_is_stationary_5;
  reg        [15:0]   io_in_c_bypass_regNext_1_2_data_5;
  reg                 io_in_c_bypass_regNext_1_2_is_stationary_5;
  reg        [15:0]   io_in_c_bypass_regNext_1_3_data_5;
  reg                 io_in_c_bypass_regNext_1_3_is_stationary_5;
  reg        [15:0]   io_in_c_bypass_regNext_2_0_data_5;
  reg                 io_in_c_bypass_regNext_2_0_is_stationary_5;
  reg        [15:0]   io_in_c_bypass_regNext_2_1_data_5;
  reg                 io_in_c_bypass_regNext_2_1_is_stationary_5;
  reg        [15:0]   io_in_c_bypass_regNext_2_2_data_5;
  reg                 io_in_c_bypass_regNext_2_2_is_stationary_5;
  reg        [15:0]   io_in_c_bypass_regNext_2_3_data_5;
  reg                 io_in_c_bypass_regNext_2_3_is_stationary_5;
  reg        [15:0]   io_in_c_bypass_regNext_3_0_data_5;
  reg                 io_in_c_bypass_regNext_3_0_is_stationary_5;
  reg        [15:0]   io_in_c_bypass_regNext_3_1_data_5;
  reg                 io_in_c_bypass_regNext_3_1_is_stationary_5;
  reg        [15:0]   io_in_c_bypass_regNext_3_2_data_5;
  reg                 io_in_c_bypass_regNext_3_2_is_stationary_5;
  reg        [15:0]   io_in_c_bypass_regNext_3_3_data_5;
  reg                 io_in_c_bypass_regNext_3_3_is_stationary_5;
  reg        [15:0]   io_in_c_bypass_regNext_4_0_data_5;
  reg                 io_in_c_bypass_regNext_4_0_is_stationary_5;
  reg        [15:0]   io_in_c_bypass_regNext_4_1_data_5;
  reg                 io_in_c_bypass_regNext_4_1_is_stationary_5;
  reg        [15:0]   io_in_c_bypass_regNext_4_2_data_5;
  reg                 io_in_c_bypass_regNext_4_2_is_stationary_5;
  reg        [15:0]   io_in_c_bypass_regNext_4_3_data_5;
  reg                 io_in_c_bypass_regNext_4_3_is_stationary_5;
  reg        [15:0]   io_in_c_bypass_regNext_5_0_data_5;
  reg                 io_in_c_bypass_regNext_5_0_is_stationary_5;
  reg        [15:0]   io_in_c_bypass_regNext_5_1_data_5;
  reg                 io_in_c_bypass_regNext_5_1_is_stationary_5;
  reg        [15:0]   io_in_c_bypass_regNext_5_2_data_5;
  reg                 io_in_c_bypass_regNext_5_2_is_stationary_5;
  reg        [15:0]   io_in_c_bypass_regNext_5_3_data_5;
  reg                 io_in_c_bypass_regNext_5_3_is_stationary_5;
  reg        [15:0]   io_in_c_bypass_regNext_6_0_data_5;
  reg                 io_in_c_bypass_regNext_6_0_is_stationary_5;
  reg        [15:0]   io_in_c_bypass_regNext_6_1_data_5;
  reg                 io_in_c_bypass_regNext_6_1_is_stationary_5;
  reg        [15:0]   io_in_c_bypass_regNext_6_2_data_5;
  reg                 io_in_c_bypass_regNext_6_2_is_stationary_5;
  reg        [15:0]   io_in_c_bypass_regNext_6_3_data_5;
  reg                 io_in_c_bypass_regNext_6_3_is_stationary_5;
  reg        [15:0]   io_in_c_bypass_regNext_7_0_data_5;
  reg                 io_in_c_bypass_regNext_7_0_is_stationary_5;
  reg        [15:0]   io_in_c_bypass_regNext_7_1_data_5;
  reg                 io_in_c_bypass_regNext_7_1_is_stationary_5;
  reg        [15:0]   io_in_c_bypass_regNext_7_2_data_5;
  reg                 io_in_c_bypass_regNext_7_2_is_stationary_5;
  reg        [15:0]   io_in_c_bypass_regNext_7_3_data_5;
  reg                 io_in_c_bypass_regNext_7_3_is_stationary_5;
  reg        [15:0]   io_in_c_bypass_regNext_8_0_data_5;
  reg                 io_in_c_bypass_regNext_8_0_is_stationary_5;
  reg        [15:0]   io_in_c_bypass_regNext_8_1_data_5;
  reg                 io_in_c_bypass_regNext_8_1_is_stationary_5;
  reg        [15:0]   io_in_c_bypass_regNext_8_2_data_5;
  reg                 io_in_c_bypass_regNext_8_2_is_stationary_5;
  reg        [15:0]   io_in_c_bypass_regNext_8_3_data_5;
  reg                 io_in_c_bypass_regNext_8_3_is_stationary_5;
  reg        [15:0]   io_in_c_bypass_regNext_9_0_data_5;
  reg                 io_in_c_bypass_regNext_9_0_is_stationary_5;
  reg        [15:0]   io_in_c_bypass_regNext_9_1_data_5;
  reg                 io_in_c_bypass_regNext_9_1_is_stationary_5;
  reg        [15:0]   io_in_c_bypass_regNext_9_2_data_5;
  reg                 io_in_c_bypass_regNext_9_2_is_stationary_5;
  reg        [15:0]   io_in_c_bypass_regNext_9_3_data_5;
  reg                 io_in_c_bypass_regNext_9_3_is_stationary_5;
  reg        [15:0]   io_in_c_bypass_regNext_10_0_data_5;
  reg                 io_in_c_bypass_regNext_10_0_is_stationary_5;
  reg        [15:0]   io_in_c_bypass_regNext_10_1_data_5;
  reg                 io_in_c_bypass_regNext_10_1_is_stationary_5;
  reg        [15:0]   io_in_c_bypass_regNext_10_2_data_5;
  reg                 io_in_c_bypass_regNext_10_2_is_stationary_5;
  reg        [15:0]   io_in_c_bypass_regNext_10_3_data_5;
  reg                 io_in_c_bypass_regNext_10_3_is_stationary_5;
  reg        [15:0]   io_in_c_bypass_regNext_11_0_data_5;
  reg                 io_in_c_bypass_regNext_11_0_is_stationary_5;
  reg        [15:0]   io_in_c_bypass_regNext_11_1_data_5;
  reg                 io_in_c_bypass_regNext_11_1_is_stationary_5;
  reg        [15:0]   io_in_c_bypass_regNext_11_2_data_5;
  reg                 io_in_c_bypass_regNext_11_2_is_stationary_5;
  reg        [15:0]   io_in_c_bypass_regNext_11_3_data_5;
  reg                 io_in_c_bypass_regNext_11_3_is_stationary_5;
  reg        [15:0]   io_in_c_bypass_regNext_12_0_data_5;
  reg                 io_in_c_bypass_regNext_12_0_is_stationary_5;
  reg        [15:0]   io_in_c_bypass_regNext_12_1_data_5;
  reg                 io_in_c_bypass_regNext_12_1_is_stationary_5;
  reg        [15:0]   io_in_c_bypass_regNext_12_2_data_5;
  reg                 io_in_c_bypass_regNext_12_2_is_stationary_5;
  reg        [15:0]   io_in_c_bypass_regNext_12_3_data_5;
  reg                 io_in_c_bypass_regNext_12_3_is_stationary_5;
  reg        [15:0]   io_in_c_bypass_regNext_13_0_data_5;
  reg                 io_in_c_bypass_regNext_13_0_is_stationary_5;
  reg        [15:0]   io_in_c_bypass_regNext_13_1_data_5;
  reg                 io_in_c_bypass_regNext_13_1_is_stationary_5;
  reg        [15:0]   io_in_c_bypass_regNext_13_2_data_5;
  reg                 io_in_c_bypass_regNext_13_2_is_stationary_5;
  reg        [15:0]   io_in_c_bypass_regNext_13_3_data_5;
  reg                 io_in_c_bypass_regNext_13_3_is_stationary_5;
  reg        [15:0]   io_in_c_bypass_regNext_14_0_data_5;
  reg                 io_in_c_bypass_regNext_14_0_is_stationary_5;
  reg        [15:0]   io_in_c_bypass_regNext_14_1_data_5;
  reg                 io_in_c_bypass_regNext_14_1_is_stationary_5;
  reg        [15:0]   io_in_c_bypass_regNext_14_2_data_5;
  reg                 io_in_c_bypass_regNext_14_2_is_stationary_5;
  reg        [15:0]   io_in_c_bypass_regNext_14_3_data_5;
  reg                 io_in_c_bypass_regNext_14_3_is_stationary_5;
  reg        [15:0]   io_in_c_bypass_regNext_15_0_data_5;
  reg                 io_in_c_bypass_regNext_15_0_is_stationary_5;
  reg        [15:0]   io_in_c_bypass_regNext_15_1_data_5;
  reg                 io_in_c_bypass_regNext_15_1_is_stationary_5;
  reg        [15:0]   io_in_c_bypass_regNext_15_2_data_5;
  reg                 io_in_c_bypass_regNext_15_2_is_stationary_5;
  reg        [15:0]   io_in_c_bypass_regNext_15_3_data_5;
  reg                 io_in_c_bypass_regNext_15_3_is_stationary_5;
  reg        [15:0]   io_in_c_bypass_regNext_16_0_data_5;
  reg                 io_in_c_bypass_regNext_16_0_is_stationary_5;
  reg        [15:0]   io_in_c_bypass_regNext_16_1_data_5;
  reg                 io_in_c_bypass_regNext_16_1_is_stationary_5;
  reg        [15:0]   io_in_c_bypass_regNext_16_2_data_5;
  reg                 io_in_c_bypass_regNext_16_2_is_stationary_5;
  reg        [15:0]   io_in_c_bypass_regNext_16_3_data_5;
  reg                 io_in_c_bypass_regNext_16_3_is_stationary_5;
  reg        [15:0]   io_in_c_bypass_regNext_17_0_data_5;
  reg                 io_in_c_bypass_regNext_17_0_is_stationary_5;
  reg        [15:0]   io_in_c_bypass_regNext_17_1_data_5;
  reg                 io_in_c_bypass_regNext_17_1_is_stationary_5;
  reg        [15:0]   io_in_c_bypass_regNext_17_2_data_5;
  reg                 io_in_c_bypass_regNext_17_2_is_stationary_5;
  reg        [15:0]   io_in_c_bypass_regNext_17_3_data_5;
  reg                 io_in_c_bypass_regNext_17_3_is_stationary_5;
  reg        [15:0]   io_in_c_bypass_regNext_18_0_data_5;
  reg                 io_in_c_bypass_regNext_18_0_is_stationary_5;
  reg        [15:0]   io_in_c_bypass_regNext_18_1_data_5;
  reg                 io_in_c_bypass_regNext_18_1_is_stationary_5;
  reg        [15:0]   io_in_c_bypass_regNext_18_2_data_5;
  reg                 io_in_c_bypass_regNext_18_2_is_stationary_5;
  reg        [15:0]   io_in_c_bypass_regNext_18_3_data_5;
  reg                 io_in_c_bypass_regNext_18_3_is_stationary_5;
  reg        [15:0]   io_in_c_bypass_regNext_19_0_data_5;
  reg                 io_in_c_bypass_regNext_19_0_is_stationary_5;
  reg        [15:0]   io_in_c_bypass_regNext_19_1_data_5;
  reg                 io_in_c_bypass_regNext_19_1_is_stationary_5;
  reg        [15:0]   io_in_c_bypass_regNext_19_2_data_5;
  reg                 io_in_c_bypass_regNext_19_2_is_stationary_5;
  reg        [15:0]   io_in_c_bypass_regNext_19_3_data_5;
  reg                 io_in_c_bypass_regNext_19_3_is_stationary_5;
  reg        [15:0]   io_in_c_bypass_regNext_20_0_data_5;
  reg                 io_in_c_bypass_regNext_20_0_is_stationary_5;
  reg        [15:0]   io_in_c_bypass_regNext_20_1_data_5;
  reg                 io_in_c_bypass_regNext_20_1_is_stationary_5;
  reg        [15:0]   io_in_c_bypass_regNext_20_2_data_5;
  reg                 io_in_c_bypass_regNext_20_2_is_stationary_5;
  reg        [15:0]   io_in_c_bypass_regNext_20_3_data_5;
  reg                 io_in_c_bypass_regNext_20_3_is_stationary_5;
  reg        [15:0]   io_in_c_bypass_regNext_21_0_data_5;
  reg                 io_in_c_bypass_regNext_21_0_is_stationary_5;
  reg        [15:0]   io_in_c_bypass_regNext_21_1_data_5;
  reg                 io_in_c_bypass_regNext_21_1_is_stationary_5;
  reg        [15:0]   io_in_c_bypass_regNext_21_2_data_5;
  reg                 io_in_c_bypass_regNext_21_2_is_stationary_5;
  reg        [15:0]   io_in_c_bypass_regNext_21_3_data_5;
  reg                 io_in_c_bypass_regNext_21_3_is_stationary_5;
  reg        [15:0]   io_in_c_bypass_regNext_22_0_data_5;
  reg                 io_in_c_bypass_regNext_22_0_is_stationary_5;
  reg        [15:0]   io_in_c_bypass_regNext_22_1_data_5;
  reg                 io_in_c_bypass_regNext_22_1_is_stationary_5;
  reg        [15:0]   io_in_c_bypass_regNext_22_2_data_5;
  reg                 io_in_c_bypass_regNext_22_2_is_stationary_5;
  reg        [15:0]   io_in_c_bypass_regNext_22_3_data_5;
  reg                 io_in_c_bypass_regNext_22_3_is_stationary_5;
  reg        [15:0]   io_in_c_bypass_regNext_23_0_data_5;
  reg                 io_in_c_bypass_regNext_23_0_is_stationary_5;
  reg        [15:0]   io_in_c_bypass_regNext_23_1_data_5;
  reg                 io_in_c_bypass_regNext_23_1_is_stationary_5;
  reg        [15:0]   io_in_c_bypass_regNext_23_2_data_5;
  reg                 io_in_c_bypass_regNext_23_2_is_stationary_5;
  reg        [15:0]   io_in_c_bypass_regNext_23_3_data_5;
  reg                 io_in_c_bypass_regNext_23_3_is_stationary_5;
  reg        [15:0]   io_in_c_bypass_regNext_24_0_data_5;
  reg                 io_in_c_bypass_regNext_24_0_is_stationary_5;
  reg        [15:0]   io_in_c_bypass_regNext_24_1_data_5;
  reg                 io_in_c_bypass_regNext_24_1_is_stationary_5;
  reg        [15:0]   io_in_c_bypass_regNext_24_2_data_5;
  reg                 io_in_c_bypass_regNext_24_2_is_stationary_5;
  reg        [15:0]   io_in_c_bypass_regNext_24_3_data_5;
  reg                 io_in_c_bypass_regNext_24_3_is_stationary_5;
  reg        [15:0]   io_in_c_bypass_regNext_25_0_data_5;
  reg                 io_in_c_bypass_regNext_25_0_is_stationary_5;
  reg        [15:0]   io_in_c_bypass_regNext_25_1_data_5;
  reg                 io_in_c_bypass_regNext_25_1_is_stationary_5;
  reg        [15:0]   io_in_c_bypass_regNext_25_2_data_5;
  reg                 io_in_c_bypass_regNext_25_2_is_stationary_5;
  reg        [15:0]   io_in_c_bypass_regNext_25_3_data_5;
  reg                 io_in_c_bypass_regNext_25_3_is_stationary_5;
  reg        [15:0]   io_in_c_bypass_regNext_26_0_data_5;
  reg                 io_in_c_bypass_regNext_26_0_is_stationary_5;
  reg        [15:0]   io_in_c_bypass_regNext_26_1_data_5;
  reg                 io_in_c_bypass_regNext_26_1_is_stationary_5;
  reg        [15:0]   io_in_c_bypass_regNext_26_2_data_5;
  reg                 io_in_c_bypass_regNext_26_2_is_stationary_5;
  reg        [15:0]   io_in_c_bypass_regNext_26_3_data_5;
  reg                 io_in_c_bypass_regNext_26_3_is_stationary_5;
  reg        [15:0]   io_in_c_bypass_regNext_27_0_data_5;
  reg                 io_in_c_bypass_regNext_27_0_is_stationary_5;
  reg        [15:0]   io_in_c_bypass_regNext_27_1_data_5;
  reg                 io_in_c_bypass_regNext_27_1_is_stationary_5;
  reg        [15:0]   io_in_c_bypass_regNext_27_2_data_5;
  reg                 io_in_c_bypass_regNext_27_2_is_stationary_5;
  reg        [15:0]   io_in_c_bypass_regNext_27_3_data_5;
  reg                 io_in_c_bypass_regNext_27_3_is_stationary_5;
  reg        [15:0]   io_in_c_bypass_regNext_28_0_data_5;
  reg                 io_in_c_bypass_regNext_28_0_is_stationary_5;
  reg        [15:0]   io_in_c_bypass_regNext_28_1_data_5;
  reg                 io_in_c_bypass_regNext_28_1_is_stationary_5;
  reg        [15:0]   io_in_c_bypass_regNext_28_2_data_5;
  reg                 io_in_c_bypass_regNext_28_2_is_stationary_5;
  reg        [15:0]   io_in_c_bypass_regNext_28_3_data_5;
  reg                 io_in_c_bypass_regNext_28_3_is_stationary_5;
  reg        [15:0]   io_in_c_bypass_regNext_29_0_data_5;
  reg                 io_in_c_bypass_regNext_29_0_is_stationary_5;
  reg        [15:0]   io_in_c_bypass_regNext_29_1_data_5;
  reg                 io_in_c_bypass_regNext_29_1_is_stationary_5;
  reg        [15:0]   io_in_c_bypass_regNext_29_2_data_5;
  reg                 io_in_c_bypass_regNext_29_2_is_stationary_5;
  reg        [15:0]   io_in_c_bypass_regNext_29_3_data_5;
  reg                 io_in_c_bypass_regNext_29_3_is_stationary_5;
  reg        [15:0]   io_in_c_bypass_regNext_30_0_data_5;
  reg                 io_in_c_bypass_regNext_30_0_is_stationary_5;
  reg        [15:0]   io_in_c_bypass_regNext_30_1_data_5;
  reg                 io_in_c_bypass_regNext_30_1_is_stationary_5;
  reg        [15:0]   io_in_c_bypass_regNext_30_2_data_5;
  reg                 io_in_c_bypass_regNext_30_2_is_stationary_5;
  reg        [15:0]   io_in_c_bypass_regNext_30_3_data_5;
  reg                 io_in_c_bypass_regNext_30_3_is_stationary_5;
  reg        [15:0]   io_in_c_bypass_regNext_31_0_data_5;
  reg                 io_in_c_bypass_regNext_31_0_is_stationary_5;
  reg        [15:0]   io_in_c_bypass_regNext_31_1_data_5;
  reg                 io_in_c_bypass_regNext_31_1_is_stationary_5;
  reg        [15:0]   io_in_c_bypass_regNext_31_2_data_5;
  reg                 io_in_c_bypass_regNext_31_2_is_stationary_5;
  reg        [15:0]   io_in_c_bypass_regNext_31_3_data_5;
  reg                 io_in_c_bypass_regNext_31_3_is_stationary_5;
  reg        [15:0]   io_in_c_bypass_regNext_0_0_data_6;
  reg                 io_in_c_bypass_regNext_0_0_is_stationary_6;
  reg        [15:0]   io_in_c_bypass_regNext_0_1_data_6;
  reg                 io_in_c_bypass_regNext_0_1_is_stationary_6;
  reg        [15:0]   io_in_c_bypass_regNext_0_2_data_6;
  reg                 io_in_c_bypass_regNext_0_2_is_stationary_6;
  reg        [15:0]   io_in_c_bypass_regNext_0_3_data_6;
  reg                 io_in_c_bypass_regNext_0_3_is_stationary_6;
  reg        [15:0]   io_in_c_bypass_regNext_1_0_data_6;
  reg                 io_in_c_bypass_regNext_1_0_is_stationary_6;
  reg        [15:0]   io_in_c_bypass_regNext_1_1_data_6;
  reg                 io_in_c_bypass_regNext_1_1_is_stationary_6;
  reg        [15:0]   io_in_c_bypass_regNext_1_2_data_6;
  reg                 io_in_c_bypass_regNext_1_2_is_stationary_6;
  reg        [15:0]   io_in_c_bypass_regNext_1_3_data_6;
  reg                 io_in_c_bypass_regNext_1_3_is_stationary_6;
  reg        [15:0]   io_in_c_bypass_regNext_2_0_data_6;
  reg                 io_in_c_bypass_regNext_2_0_is_stationary_6;
  reg        [15:0]   io_in_c_bypass_regNext_2_1_data_6;
  reg                 io_in_c_bypass_regNext_2_1_is_stationary_6;
  reg        [15:0]   io_in_c_bypass_regNext_2_2_data_6;
  reg                 io_in_c_bypass_regNext_2_2_is_stationary_6;
  reg        [15:0]   io_in_c_bypass_regNext_2_3_data_6;
  reg                 io_in_c_bypass_regNext_2_3_is_stationary_6;
  reg        [15:0]   io_in_c_bypass_regNext_3_0_data_6;
  reg                 io_in_c_bypass_regNext_3_0_is_stationary_6;
  reg        [15:0]   io_in_c_bypass_regNext_3_1_data_6;
  reg                 io_in_c_bypass_regNext_3_1_is_stationary_6;
  reg        [15:0]   io_in_c_bypass_regNext_3_2_data_6;
  reg                 io_in_c_bypass_regNext_3_2_is_stationary_6;
  reg        [15:0]   io_in_c_bypass_regNext_3_3_data_6;
  reg                 io_in_c_bypass_regNext_3_3_is_stationary_6;
  reg        [15:0]   io_in_c_bypass_regNext_4_0_data_6;
  reg                 io_in_c_bypass_regNext_4_0_is_stationary_6;
  reg        [15:0]   io_in_c_bypass_regNext_4_1_data_6;
  reg                 io_in_c_bypass_regNext_4_1_is_stationary_6;
  reg        [15:0]   io_in_c_bypass_regNext_4_2_data_6;
  reg                 io_in_c_bypass_regNext_4_2_is_stationary_6;
  reg        [15:0]   io_in_c_bypass_regNext_4_3_data_6;
  reg                 io_in_c_bypass_regNext_4_3_is_stationary_6;
  reg        [15:0]   io_in_c_bypass_regNext_5_0_data_6;
  reg                 io_in_c_bypass_regNext_5_0_is_stationary_6;
  reg        [15:0]   io_in_c_bypass_regNext_5_1_data_6;
  reg                 io_in_c_bypass_regNext_5_1_is_stationary_6;
  reg        [15:0]   io_in_c_bypass_regNext_5_2_data_6;
  reg                 io_in_c_bypass_regNext_5_2_is_stationary_6;
  reg        [15:0]   io_in_c_bypass_regNext_5_3_data_6;
  reg                 io_in_c_bypass_regNext_5_3_is_stationary_6;
  reg        [15:0]   io_in_c_bypass_regNext_6_0_data_6;
  reg                 io_in_c_bypass_regNext_6_0_is_stationary_6;
  reg        [15:0]   io_in_c_bypass_regNext_6_1_data_6;
  reg                 io_in_c_bypass_regNext_6_1_is_stationary_6;
  reg        [15:0]   io_in_c_bypass_regNext_6_2_data_6;
  reg                 io_in_c_bypass_regNext_6_2_is_stationary_6;
  reg        [15:0]   io_in_c_bypass_regNext_6_3_data_6;
  reg                 io_in_c_bypass_regNext_6_3_is_stationary_6;
  reg        [15:0]   io_in_c_bypass_regNext_7_0_data_6;
  reg                 io_in_c_bypass_regNext_7_0_is_stationary_6;
  reg        [15:0]   io_in_c_bypass_regNext_7_1_data_6;
  reg                 io_in_c_bypass_regNext_7_1_is_stationary_6;
  reg        [15:0]   io_in_c_bypass_regNext_7_2_data_6;
  reg                 io_in_c_bypass_regNext_7_2_is_stationary_6;
  reg        [15:0]   io_in_c_bypass_regNext_7_3_data_6;
  reg                 io_in_c_bypass_regNext_7_3_is_stationary_6;
  reg        [15:0]   io_in_c_bypass_regNext_8_0_data_6;
  reg                 io_in_c_bypass_regNext_8_0_is_stationary_6;
  reg        [15:0]   io_in_c_bypass_regNext_8_1_data_6;
  reg                 io_in_c_bypass_regNext_8_1_is_stationary_6;
  reg        [15:0]   io_in_c_bypass_regNext_8_2_data_6;
  reg                 io_in_c_bypass_regNext_8_2_is_stationary_6;
  reg        [15:0]   io_in_c_bypass_regNext_8_3_data_6;
  reg                 io_in_c_bypass_regNext_8_3_is_stationary_6;
  reg        [15:0]   io_in_c_bypass_regNext_9_0_data_6;
  reg                 io_in_c_bypass_regNext_9_0_is_stationary_6;
  reg        [15:0]   io_in_c_bypass_regNext_9_1_data_6;
  reg                 io_in_c_bypass_regNext_9_1_is_stationary_6;
  reg        [15:0]   io_in_c_bypass_regNext_9_2_data_6;
  reg                 io_in_c_bypass_regNext_9_2_is_stationary_6;
  reg        [15:0]   io_in_c_bypass_regNext_9_3_data_6;
  reg                 io_in_c_bypass_regNext_9_3_is_stationary_6;
  reg        [15:0]   io_in_c_bypass_regNext_10_0_data_6;
  reg                 io_in_c_bypass_regNext_10_0_is_stationary_6;
  reg        [15:0]   io_in_c_bypass_regNext_10_1_data_6;
  reg                 io_in_c_bypass_regNext_10_1_is_stationary_6;
  reg        [15:0]   io_in_c_bypass_regNext_10_2_data_6;
  reg                 io_in_c_bypass_regNext_10_2_is_stationary_6;
  reg        [15:0]   io_in_c_bypass_regNext_10_3_data_6;
  reg                 io_in_c_bypass_regNext_10_3_is_stationary_6;
  reg        [15:0]   io_in_c_bypass_regNext_11_0_data_6;
  reg                 io_in_c_bypass_regNext_11_0_is_stationary_6;
  reg        [15:0]   io_in_c_bypass_regNext_11_1_data_6;
  reg                 io_in_c_bypass_regNext_11_1_is_stationary_6;
  reg        [15:0]   io_in_c_bypass_regNext_11_2_data_6;
  reg                 io_in_c_bypass_regNext_11_2_is_stationary_6;
  reg        [15:0]   io_in_c_bypass_regNext_11_3_data_6;
  reg                 io_in_c_bypass_regNext_11_3_is_stationary_6;
  reg        [15:0]   io_in_c_bypass_regNext_12_0_data_6;
  reg                 io_in_c_bypass_regNext_12_0_is_stationary_6;
  reg        [15:0]   io_in_c_bypass_regNext_12_1_data_6;
  reg                 io_in_c_bypass_regNext_12_1_is_stationary_6;
  reg        [15:0]   io_in_c_bypass_regNext_12_2_data_6;
  reg                 io_in_c_bypass_regNext_12_2_is_stationary_6;
  reg        [15:0]   io_in_c_bypass_regNext_12_3_data_6;
  reg                 io_in_c_bypass_regNext_12_3_is_stationary_6;
  reg        [15:0]   io_in_c_bypass_regNext_13_0_data_6;
  reg                 io_in_c_bypass_regNext_13_0_is_stationary_6;
  reg        [15:0]   io_in_c_bypass_regNext_13_1_data_6;
  reg                 io_in_c_bypass_regNext_13_1_is_stationary_6;
  reg        [15:0]   io_in_c_bypass_regNext_13_2_data_6;
  reg                 io_in_c_bypass_regNext_13_2_is_stationary_6;
  reg        [15:0]   io_in_c_bypass_regNext_13_3_data_6;
  reg                 io_in_c_bypass_regNext_13_3_is_stationary_6;
  reg        [15:0]   io_in_c_bypass_regNext_14_0_data_6;
  reg                 io_in_c_bypass_regNext_14_0_is_stationary_6;
  reg        [15:0]   io_in_c_bypass_regNext_14_1_data_6;
  reg                 io_in_c_bypass_regNext_14_1_is_stationary_6;
  reg        [15:0]   io_in_c_bypass_regNext_14_2_data_6;
  reg                 io_in_c_bypass_regNext_14_2_is_stationary_6;
  reg        [15:0]   io_in_c_bypass_regNext_14_3_data_6;
  reg                 io_in_c_bypass_regNext_14_3_is_stationary_6;
  reg        [15:0]   io_in_c_bypass_regNext_15_0_data_6;
  reg                 io_in_c_bypass_regNext_15_0_is_stationary_6;
  reg        [15:0]   io_in_c_bypass_regNext_15_1_data_6;
  reg                 io_in_c_bypass_regNext_15_1_is_stationary_6;
  reg        [15:0]   io_in_c_bypass_regNext_15_2_data_6;
  reg                 io_in_c_bypass_regNext_15_2_is_stationary_6;
  reg        [15:0]   io_in_c_bypass_regNext_15_3_data_6;
  reg                 io_in_c_bypass_regNext_15_3_is_stationary_6;
  reg        [15:0]   io_in_c_bypass_regNext_16_0_data_6;
  reg                 io_in_c_bypass_regNext_16_0_is_stationary_6;
  reg        [15:0]   io_in_c_bypass_regNext_16_1_data_6;
  reg                 io_in_c_bypass_regNext_16_1_is_stationary_6;
  reg        [15:0]   io_in_c_bypass_regNext_16_2_data_6;
  reg                 io_in_c_bypass_regNext_16_2_is_stationary_6;
  reg        [15:0]   io_in_c_bypass_regNext_16_3_data_6;
  reg                 io_in_c_bypass_regNext_16_3_is_stationary_6;
  reg        [15:0]   io_in_c_bypass_regNext_17_0_data_6;
  reg                 io_in_c_bypass_regNext_17_0_is_stationary_6;
  reg        [15:0]   io_in_c_bypass_regNext_17_1_data_6;
  reg                 io_in_c_bypass_regNext_17_1_is_stationary_6;
  reg        [15:0]   io_in_c_bypass_regNext_17_2_data_6;
  reg                 io_in_c_bypass_regNext_17_2_is_stationary_6;
  reg        [15:0]   io_in_c_bypass_regNext_17_3_data_6;
  reg                 io_in_c_bypass_regNext_17_3_is_stationary_6;
  reg        [15:0]   io_in_c_bypass_regNext_18_0_data_6;
  reg                 io_in_c_bypass_regNext_18_0_is_stationary_6;
  reg        [15:0]   io_in_c_bypass_regNext_18_1_data_6;
  reg                 io_in_c_bypass_regNext_18_1_is_stationary_6;
  reg        [15:0]   io_in_c_bypass_regNext_18_2_data_6;
  reg                 io_in_c_bypass_regNext_18_2_is_stationary_6;
  reg        [15:0]   io_in_c_bypass_regNext_18_3_data_6;
  reg                 io_in_c_bypass_regNext_18_3_is_stationary_6;
  reg        [15:0]   io_in_c_bypass_regNext_19_0_data_6;
  reg                 io_in_c_bypass_regNext_19_0_is_stationary_6;
  reg        [15:0]   io_in_c_bypass_regNext_19_1_data_6;
  reg                 io_in_c_bypass_regNext_19_1_is_stationary_6;
  reg        [15:0]   io_in_c_bypass_regNext_19_2_data_6;
  reg                 io_in_c_bypass_regNext_19_2_is_stationary_6;
  reg        [15:0]   io_in_c_bypass_regNext_19_3_data_6;
  reg                 io_in_c_bypass_regNext_19_3_is_stationary_6;
  reg        [15:0]   io_in_c_bypass_regNext_20_0_data_6;
  reg                 io_in_c_bypass_regNext_20_0_is_stationary_6;
  reg        [15:0]   io_in_c_bypass_regNext_20_1_data_6;
  reg                 io_in_c_bypass_regNext_20_1_is_stationary_6;
  reg        [15:0]   io_in_c_bypass_regNext_20_2_data_6;
  reg                 io_in_c_bypass_regNext_20_2_is_stationary_6;
  reg        [15:0]   io_in_c_bypass_regNext_20_3_data_6;
  reg                 io_in_c_bypass_regNext_20_3_is_stationary_6;
  reg        [15:0]   io_in_c_bypass_regNext_21_0_data_6;
  reg                 io_in_c_bypass_regNext_21_0_is_stationary_6;
  reg        [15:0]   io_in_c_bypass_regNext_21_1_data_6;
  reg                 io_in_c_bypass_regNext_21_1_is_stationary_6;
  reg        [15:0]   io_in_c_bypass_regNext_21_2_data_6;
  reg                 io_in_c_bypass_regNext_21_2_is_stationary_6;
  reg        [15:0]   io_in_c_bypass_regNext_21_3_data_6;
  reg                 io_in_c_bypass_regNext_21_3_is_stationary_6;
  reg        [15:0]   io_in_c_bypass_regNext_22_0_data_6;
  reg                 io_in_c_bypass_regNext_22_0_is_stationary_6;
  reg        [15:0]   io_in_c_bypass_regNext_22_1_data_6;
  reg                 io_in_c_bypass_regNext_22_1_is_stationary_6;
  reg        [15:0]   io_in_c_bypass_regNext_22_2_data_6;
  reg                 io_in_c_bypass_regNext_22_2_is_stationary_6;
  reg        [15:0]   io_in_c_bypass_regNext_22_3_data_6;
  reg                 io_in_c_bypass_regNext_22_3_is_stationary_6;
  reg        [15:0]   io_in_c_bypass_regNext_23_0_data_6;
  reg                 io_in_c_bypass_regNext_23_0_is_stationary_6;
  reg        [15:0]   io_in_c_bypass_regNext_23_1_data_6;
  reg                 io_in_c_bypass_regNext_23_1_is_stationary_6;
  reg        [15:0]   io_in_c_bypass_regNext_23_2_data_6;
  reg                 io_in_c_bypass_regNext_23_2_is_stationary_6;
  reg        [15:0]   io_in_c_bypass_regNext_23_3_data_6;
  reg                 io_in_c_bypass_regNext_23_3_is_stationary_6;
  reg        [15:0]   io_in_c_bypass_regNext_24_0_data_6;
  reg                 io_in_c_bypass_regNext_24_0_is_stationary_6;
  reg        [15:0]   io_in_c_bypass_regNext_24_1_data_6;
  reg                 io_in_c_bypass_regNext_24_1_is_stationary_6;
  reg        [15:0]   io_in_c_bypass_regNext_24_2_data_6;
  reg                 io_in_c_bypass_regNext_24_2_is_stationary_6;
  reg        [15:0]   io_in_c_bypass_regNext_24_3_data_6;
  reg                 io_in_c_bypass_regNext_24_3_is_stationary_6;
  reg        [15:0]   io_in_c_bypass_regNext_25_0_data_6;
  reg                 io_in_c_bypass_regNext_25_0_is_stationary_6;
  reg        [15:0]   io_in_c_bypass_regNext_25_1_data_6;
  reg                 io_in_c_bypass_regNext_25_1_is_stationary_6;
  reg        [15:0]   io_in_c_bypass_regNext_25_2_data_6;
  reg                 io_in_c_bypass_regNext_25_2_is_stationary_6;
  reg        [15:0]   io_in_c_bypass_regNext_25_3_data_6;
  reg                 io_in_c_bypass_regNext_25_3_is_stationary_6;
  reg        [15:0]   io_in_c_bypass_regNext_26_0_data_6;
  reg                 io_in_c_bypass_regNext_26_0_is_stationary_6;
  reg        [15:0]   io_in_c_bypass_regNext_26_1_data_6;
  reg                 io_in_c_bypass_regNext_26_1_is_stationary_6;
  reg        [15:0]   io_in_c_bypass_regNext_26_2_data_6;
  reg                 io_in_c_bypass_regNext_26_2_is_stationary_6;
  reg        [15:0]   io_in_c_bypass_regNext_26_3_data_6;
  reg                 io_in_c_bypass_regNext_26_3_is_stationary_6;
  reg        [15:0]   io_in_c_bypass_regNext_27_0_data_6;
  reg                 io_in_c_bypass_regNext_27_0_is_stationary_6;
  reg        [15:0]   io_in_c_bypass_regNext_27_1_data_6;
  reg                 io_in_c_bypass_regNext_27_1_is_stationary_6;
  reg        [15:0]   io_in_c_bypass_regNext_27_2_data_6;
  reg                 io_in_c_bypass_regNext_27_2_is_stationary_6;
  reg        [15:0]   io_in_c_bypass_regNext_27_3_data_6;
  reg                 io_in_c_bypass_regNext_27_3_is_stationary_6;
  reg        [15:0]   io_in_c_bypass_regNext_28_0_data_6;
  reg                 io_in_c_bypass_regNext_28_0_is_stationary_6;
  reg        [15:0]   io_in_c_bypass_regNext_28_1_data_6;
  reg                 io_in_c_bypass_regNext_28_1_is_stationary_6;
  reg        [15:0]   io_in_c_bypass_regNext_28_2_data_6;
  reg                 io_in_c_bypass_regNext_28_2_is_stationary_6;
  reg        [15:0]   io_in_c_bypass_regNext_28_3_data_6;
  reg                 io_in_c_bypass_regNext_28_3_is_stationary_6;
  reg        [15:0]   io_in_c_bypass_regNext_29_0_data_6;
  reg                 io_in_c_bypass_regNext_29_0_is_stationary_6;
  reg        [15:0]   io_in_c_bypass_regNext_29_1_data_6;
  reg                 io_in_c_bypass_regNext_29_1_is_stationary_6;
  reg        [15:0]   io_in_c_bypass_regNext_29_2_data_6;
  reg                 io_in_c_bypass_regNext_29_2_is_stationary_6;
  reg        [15:0]   io_in_c_bypass_regNext_29_3_data_6;
  reg                 io_in_c_bypass_regNext_29_3_is_stationary_6;
  reg        [15:0]   io_in_c_bypass_regNext_30_0_data_6;
  reg                 io_in_c_bypass_regNext_30_0_is_stationary_6;
  reg        [15:0]   io_in_c_bypass_regNext_30_1_data_6;
  reg                 io_in_c_bypass_regNext_30_1_is_stationary_6;
  reg        [15:0]   io_in_c_bypass_regNext_30_2_data_6;
  reg                 io_in_c_bypass_regNext_30_2_is_stationary_6;
  reg        [15:0]   io_in_c_bypass_regNext_30_3_data_6;
  reg                 io_in_c_bypass_regNext_30_3_is_stationary_6;
  reg        [15:0]   io_in_c_bypass_regNext_31_0_data_6;
  reg                 io_in_c_bypass_regNext_31_0_is_stationary_6;
  reg        [15:0]   io_in_c_bypass_regNext_31_1_data_6;
  reg                 io_in_c_bypass_regNext_31_1_is_stationary_6;
  reg        [15:0]   io_in_c_bypass_regNext_31_2_data_6;
  reg                 io_in_c_bypass_regNext_31_2_is_stationary_6;
  reg        [15:0]   io_in_c_bypass_regNext_31_3_data_6;
  reg                 io_in_c_bypass_regNext_31_3_is_stationary_6;
  reg        [15:0]   io_in_c_bypass_regNext_0_0_data_7;
  reg                 io_in_c_bypass_regNext_0_0_is_stationary_7;
  reg        [15:0]   io_in_c_bypass_regNext_0_1_data_7;
  reg                 io_in_c_bypass_regNext_0_1_is_stationary_7;
  reg        [15:0]   io_in_c_bypass_regNext_0_2_data_7;
  reg                 io_in_c_bypass_regNext_0_2_is_stationary_7;
  reg        [15:0]   io_in_c_bypass_regNext_0_3_data_7;
  reg                 io_in_c_bypass_regNext_0_3_is_stationary_7;
  reg        [15:0]   io_in_c_bypass_regNext_1_0_data_7;
  reg                 io_in_c_bypass_regNext_1_0_is_stationary_7;
  reg        [15:0]   io_in_c_bypass_regNext_1_1_data_7;
  reg                 io_in_c_bypass_regNext_1_1_is_stationary_7;
  reg        [15:0]   io_in_c_bypass_regNext_1_2_data_7;
  reg                 io_in_c_bypass_regNext_1_2_is_stationary_7;
  reg        [15:0]   io_in_c_bypass_regNext_1_3_data_7;
  reg                 io_in_c_bypass_regNext_1_3_is_stationary_7;
  reg        [15:0]   io_in_c_bypass_regNext_2_0_data_7;
  reg                 io_in_c_bypass_regNext_2_0_is_stationary_7;
  reg        [15:0]   io_in_c_bypass_regNext_2_1_data_7;
  reg                 io_in_c_bypass_regNext_2_1_is_stationary_7;
  reg        [15:0]   io_in_c_bypass_regNext_2_2_data_7;
  reg                 io_in_c_bypass_regNext_2_2_is_stationary_7;
  reg        [15:0]   io_in_c_bypass_regNext_2_3_data_7;
  reg                 io_in_c_bypass_regNext_2_3_is_stationary_7;
  reg        [15:0]   io_in_c_bypass_regNext_3_0_data_7;
  reg                 io_in_c_bypass_regNext_3_0_is_stationary_7;
  reg        [15:0]   io_in_c_bypass_regNext_3_1_data_7;
  reg                 io_in_c_bypass_regNext_3_1_is_stationary_7;
  reg        [15:0]   io_in_c_bypass_regNext_3_2_data_7;
  reg                 io_in_c_bypass_regNext_3_2_is_stationary_7;
  reg        [15:0]   io_in_c_bypass_regNext_3_3_data_7;
  reg                 io_in_c_bypass_regNext_3_3_is_stationary_7;
  reg        [15:0]   io_in_c_bypass_regNext_4_0_data_7;
  reg                 io_in_c_bypass_regNext_4_0_is_stationary_7;
  reg        [15:0]   io_in_c_bypass_regNext_4_1_data_7;
  reg                 io_in_c_bypass_regNext_4_1_is_stationary_7;
  reg        [15:0]   io_in_c_bypass_regNext_4_2_data_7;
  reg                 io_in_c_bypass_regNext_4_2_is_stationary_7;
  reg        [15:0]   io_in_c_bypass_regNext_4_3_data_7;
  reg                 io_in_c_bypass_regNext_4_3_is_stationary_7;
  reg        [15:0]   io_in_c_bypass_regNext_5_0_data_7;
  reg                 io_in_c_bypass_regNext_5_0_is_stationary_7;
  reg        [15:0]   io_in_c_bypass_regNext_5_1_data_7;
  reg                 io_in_c_bypass_regNext_5_1_is_stationary_7;
  reg        [15:0]   io_in_c_bypass_regNext_5_2_data_7;
  reg                 io_in_c_bypass_regNext_5_2_is_stationary_7;
  reg        [15:0]   io_in_c_bypass_regNext_5_3_data_7;
  reg                 io_in_c_bypass_regNext_5_3_is_stationary_7;
  reg        [15:0]   io_in_c_bypass_regNext_6_0_data_7;
  reg                 io_in_c_bypass_regNext_6_0_is_stationary_7;
  reg        [15:0]   io_in_c_bypass_regNext_6_1_data_7;
  reg                 io_in_c_bypass_regNext_6_1_is_stationary_7;
  reg        [15:0]   io_in_c_bypass_regNext_6_2_data_7;
  reg                 io_in_c_bypass_regNext_6_2_is_stationary_7;
  reg        [15:0]   io_in_c_bypass_regNext_6_3_data_7;
  reg                 io_in_c_bypass_regNext_6_3_is_stationary_7;
  reg        [15:0]   io_in_c_bypass_regNext_7_0_data_7;
  reg                 io_in_c_bypass_regNext_7_0_is_stationary_7;
  reg        [15:0]   io_in_c_bypass_regNext_7_1_data_7;
  reg                 io_in_c_bypass_regNext_7_1_is_stationary_7;
  reg        [15:0]   io_in_c_bypass_regNext_7_2_data_7;
  reg                 io_in_c_bypass_regNext_7_2_is_stationary_7;
  reg        [15:0]   io_in_c_bypass_regNext_7_3_data_7;
  reg                 io_in_c_bypass_regNext_7_3_is_stationary_7;
  reg        [15:0]   io_in_c_bypass_regNext_8_0_data_7;
  reg                 io_in_c_bypass_regNext_8_0_is_stationary_7;
  reg        [15:0]   io_in_c_bypass_regNext_8_1_data_7;
  reg                 io_in_c_bypass_regNext_8_1_is_stationary_7;
  reg        [15:0]   io_in_c_bypass_regNext_8_2_data_7;
  reg                 io_in_c_bypass_regNext_8_2_is_stationary_7;
  reg        [15:0]   io_in_c_bypass_regNext_8_3_data_7;
  reg                 io_in_c_bypass_regNext_8_3_is_stationary_7;
  reg        [15:0]   io_in_c_bypass_regNext_9_0_data_7;
  reg                 io_in_c_bypass_regNext_9_0_is_stationary_7;
  reg        [15:0]   io_in_c_bypass_regNext_9_1_data_7;
  reg                 io_in_c_bypass_regNext_9_1_is_stationary_7;
  reg        [15:0]   io_in_c_bypass_regNext_9_2_data_7;
  reg                 io_in_c_bypass_regNext_9_2_is_stationary_7;
  reg        [15:0]   io_in_c_bypass_regNext_9_3_data_7;
  reg                 io_in_c_bypass_regNext_9_3_is_stationary_7;
  reg        [15:0]   io_in_c_bypass_regNext_10_0_data_7;
  reg                 io_in_c_bypass_regNext_10_0_is_stationary_7;
  reg        [15:0]   io_in_c_bypass_regNext_10_1_data_7;
  reg                 io_in_c_bypass_regNext_10_1_is_stationary_7;
  reg        [15:0]   io_in_c_bypass_regNext_10_2_data_7;
  reg                 io_in_c_bypass_regNext_10_2_is_stationary_7;
  reg        [15:0]   io_in_c_bypass_regNext_10_3_data_7;
  reg                 io_in_c_bypass_regNext_10_3_is_stationary_7;
  reg        [15:0]   io_in_c_bypass_regNext_11_0_data_7;
  reg                 io_in_c_bypass_regNext_11_0_is_stationary_7;
  reg        [15:0]   io_in_c_bypass_regNext_11_1_data_7;
  reg                 io_in_c_bypass_regNext_11_1_is_stationary_7;
  reg        [15:0]   io_in_c_bypass_regNext_11_2_data_7;
  reg                 io_in_c_bypass_regNext_11_2_is_stationary_7;
  reg        [15:0]   io_in_c_bypass_regNext_11_3_data_7;
  reg                 io_in_c_bypass_regNext_11_3_is_stationary_7;
  reg        [15:0]   io_in_c_bypass_regNext_12_0_data_7;
  reg                 io_in_c_bypass_regNext_12_0_is_stationary_7;
  reg        [15:0]   io_in_c_bypass_regNext_12_1_data_7;
  reg                 io_in_c_bypass_regNext_12_1_is_stationary_7;
  reg        [15:0]   io_in_c_bypass_regNext_12_2_data_7;
  reg                 io_in_c_bypass_regNext_12_2_is_stationary_7;
  reg        [15:0]   io_in_c_bypass_regNext_12_3_data_7;
  reg                 io_in_c_bypass_regNext_12_3_is_stationary_7;
  reg        [15:0]   io_in_c_bypass_regNext_13_0_data_7;
  reg                 io_in_c_bypass_regNext_13_0_is_stationary_7;
  reg        [15:0]   io_in_c_bypass_regNext_13_1_data_7;
  reg                 io_in_c_bypass_regNext_13_1_is_stationary_7;
  reg        [15:0]   io_in_c_bypass_regNext_13_2_data_7;
  reg                 io_in_c_bypass_regNext_13_2_is_stationary_7;
  reg        [15:0]   io_in_c_bypass_regNext_13_3_data_7;
  reg                 io_in_c_bypass_regNext_13_3_is_stationary_7;
  reg        [15:0]   io_in_c_bypass_regNext_14_0_data_7;
  reg                 io_in_c_bypass_regNext_14_0_is_stationary_7;
  reg        [15:0]   io_in_c_bypass_regNext_14_1_data_7;
  reg                 io_in_c_bypass_regNext_14_1_is_stationary_7;
  reg        [15:0]   io_in_c_bypass_regNext_14_2_data_7;
  reg                 io_in_c_bypass_regNext_14_2_is_stationary_7;
  reg        [15:0]   io_in_c_bypass_regNext_14_3_data_7;
  reg                 io_in_c_bypass_regNext_14_3_is_stationary_7;
  reg        [15:0]   io_in_c_bypass_regNext_15_0_data_7;
  reg                 io_in_c_bypass_regNext_15_0_is_stationary_7;
  reg        [15:0]   io_in_c_bypass_regNext_15_1_data_7;
  reg                 io_in_c_bypass_regNext_15_1_is_stationary_7;
  reg        [15:0]   io_in_c_bypass_regNext_15_2_data_7;
  reg                 io_in_c_bypass_regNext_15_2_is_stationary_7;
  reg        [15:0]   io_in_c_bypass_regNext_15_3_data_7;
  reg                 io_in_c_bypass_regNext_15_3_is_stationary_7;
  reg        [15:0]   io_in_c_bypass_regNext_16_0_data_7;
  reg                 io_in_c_bypass_regNext_16_0_is_stationary_7;
  reg        [15:0]   io_in_c_bypass_regNext_16_1_data_7;
  reg                 io_in_c_bypass_regNext_16_1_is_stationary_7;
  reg        [15:0]   io_in_c_bypass_regNext_16_2_data_7;
  reg                 io_in_c_bypass_regNext_16_2_is_stationary_7;
  reg        [15:0]   io_in_c_bypass_regNext_16_3_data_7;
  reg                 io_in_c_bypass_regNext_16_3_is_stationary_7;
  reg        [15:0]   io_in_c_bypass_regNext_17_0_data_7;
  reg                 io_in_c_bypass_regNext_17_0_is_stationary_7;
  reg        [15:0]   io_in_c_bypass_regNext_17_1_data_7;
  reg                 io_in_c_bypass_regNext_17_1_is_stationary_7;
  reg        [15:0]   io_in_c_bypass_regNext_17_2_data_7;
  reg                 io_in_c_bypass_regNext_17_2_is_stationary_7;
  reg        [15:0]   io_in_c_bypass_regNext_17_3_data_7;
  reg                 io_in_c_bypass_regNext_17_3_is_stationary_7;
  reg        [15:0]   io_in_c_bypass_regNext_18_0_data_7;
  reg                 io_in_c_bypass_regNext_18_0_is_stationary_7;
  reg        [15:0]   io_in_c_bypass_regNext_18_1_data_7;
  reg                 io_in_c_bypass_regNext_18_1_is_stationary_7;
  reg        [15:0]   io_in_c_bypass_regNext_18_2_data_7;
  reg                 io_in_c_bypass_regNext_18_2_is_stationary_7;
  reg        [15:0]   io_in_c_bypass_regNext_18_3_data_7;
  reg                 io_in_c_bypass_regNext_18_3_is_stationary_7;
  reg        [15:0]   io_in_c_bypass_regNext_19_0_data_7;
  reg                 io_in_c_bypass_regNext_19_0_is_stationary_7;
  reg        [15:0]   io_in_c_bypass_regNext_19_1_data_7;
  reg                 io_in_c_bypass_regNext_19_1_is_stationary_7;
  reg        [15:0]   io_in_c_bypass_regNext_19_2_data_7;
  reg                 io_in_c_bypass_regNext_19_2_is_stationary_7;
  reg        [15:0]   io_in_c_bypass_regNext_19_3_data_7;
  reg                 io_in_c_bypass_regNext_19_3_is_stationary_7;
  reg        [15:0]   io_in_c_bypass_regNext_20_0_data_7;
  reg                 io_in_c_bypass_regNext_20_0_is_stationary_7;
  reg        [15:0]   io_in_c_bypass_regNext_20_1_data_7;
  reg                 io_in_c_bypass_regNext_20_1_is_stationary_7;
  reg        [15:0]   io_in_c_bypass_regNext_20_2_data_7;
  reg                 io_in_c_bypass_regNext_20_2_is_stationary_7;
  reg        [15:0]   io_in_c_bypass_regNext_20_3_data_7;
  reg                 io_in_c_bypass_regNext_20_3_is_stationary_7;
  reg        [15:0]   io_in_c_bypass_regNext_21_0_data_7;
  reg                 io_in_c_bypass_regNext_21_0_is_stationary_7;
  reg        [15:0]   io_in_c_bypass_regNext_21_1_data_7;
  reg                 io_in_c_bypass_regNext_21_1_is_stationary_7;
  reg        [15:0]   io_in_c_bypass_regNext_21_2_data_7;
  reg                 io_in_c_bypass_regNext_21_2_is_stationary_7;
  reg        [15:0]   io_in_c_bypass_regNext_21_3_data_7;
  reg                 io_in_c_bypass_regNext_21_3_is_stationary_7;
  reg        [15:0]   io_in_c_bypass_regNext_22_0_data_7;
  reg                 io_in_c_bypass_regNext_22_0_is_stationary_7;
  reg        [15:0]   io_in_c_bypass_regNext_22_1_data_7;
  reg                 io_in_c_bypass_regNext_22_1_is_stationary_7;
  reg        [15:0]   io_in_c_bypass_regNext_22_2_data_7;
  reg                 io_in_c_bypass_regNext_22_2_is_stationary_7;
  reg        [15:0]   io_in_c_bypass_regNext_22_3_data_7;
  reg                 io_in_c_bypass_regNext_22_3_is_stationary_7;
  reg        [15:0]   io_in_c_bypass_regNext_23_0_data_7;
  reg                 io_in_c_bypass_regNext_23_0_is_stationary_7;
  reg        [15:0]   io_in_c_bypass_regNext_23_1_data_7;
  reg                 io_in_c_bypass_regNext_23_1_is_stationary_7;
  reg        [15:0]   io_in_c_bypass_regNext_23_2_data_7;
  reg                 io_in_c_bypass_regNext_23_2_is_stationary_7;
  reg        [15:0]   io_in_c_bypass_regNext_23_3_data_7;
  reg                 io_in_c_bypass_regNext_23_3_is_stationary_7;
  reg        [15:0]   io_in_c_bypass_regNext_24_0_data_7;
  reg                 io_in_c_bypass_regNext_24_0_is_stationary_7;
  reg        [15:0]   io_in_c_bypass_regNext_24_1_data_7;
  reg                 io_in_c_bypass_regNext_24_1_is_stationary_7;
  reg        [15:0]   io_in_c_bypass_regNext_24_2_data_7;
  reg                 io_in_c_bypass_regNext_24_2_is_stationary_7;
  reg        [15:0]   io_in_c_bypass_regNext_24_3_data_7;
  reg                 io_in_c_bypass_regNext_24_3_is_stationary_7;
  reg        [15:0]   io_in_c_bypass_regNext_25_0_data_7;
  reg                 io_in_c_bypass_regNext_25_0_is_stationary_7;
  reg        [15:0]   io_in_c_bypass_regNext_25_1_data_7;
  reg                 io_in_c_bypass_regNext_25_1_is_stationary_7;
  reg        [15:0]   io_in_c_bypass_regNext_25_2_data_7;
  reg                 io_in_c_bypass_regNext_25_2_is_stationary_7;
  reg        [15:0]   io_in_c_bypass_regNext_25_3_data_7;
  reg                 io_in_c_bypass_regNext_25_3_is_stationary_7;
  reg        [15:0]   io_in_c_bypass_regNext_26_0_data_7;
  reg                 io_in_c_bypass_regNext_26_0_is_stationary_7;
  reg        [15:0]   io_in_c_bypass_regNext_26_1_data_7;
  reg                 io_in_c_bypass_regNext_26_1_is_stationary_7;
  reg        [15:0]   io_in_c_bypass_regNext_26_2_data_7;
  reg                 io_in_c_bypass_regNext_26_2_is_stationary_7;
  reg        [15:0]   io_in_c_bypass_regNext_26_3_data_7;
  reg                 io_in_c_bypass_regNext_26_3_is_stationary_7;
  reg        [15:0]   io_in_c_bypass_regNext_27_0_data_7;
  reg                 io_in_c_bypass_regNext_27_0_is_stationary_7;
  reg        [15:0]   io_in_c_bypass_regNext_27_1_data_7;
  reg                 io_in_c_bypass_regNext_27_1_is_stationary_7;
  reg        [15:0]   io_in_c_bypass_regNext_27_2_data_7;
  reg                 io_in_c_bypass_regNext_27_2_is_stationary_7;
  reg        [15:0]   io_in_c_bypass_regNext_27_3_data_7;
  reg                 io_in_c_bypass_regNext_27_3_is_stationary_7;
  reg        [15:0]   io_in_c_bypass_regNext_28_0_data_7;
  reg                 io_in_c_bypass_regNext_28_0_is_stationary_7;
  reg        [15:0]   io_in_c_bypass_regNext_28_1_data_7;
  reg                 io_in_c_bypass_regNext_28_1_is_stationary_7;
  reg        [15:0]   io_in_c_bypass_regNext_28_2_data_7;
  reg                 io_in_c_bypass_regNext_28_2_is_stationary_7;
  reg        [15:0]   io_in_c_bypass_regNext_28_3_data_7;
  reg                 io_in_c_bypass_regNext_28_3_is_stationary_7;
  reg        [15:0]   io_in_c_bypass_regNext_29_0_data_7;
  reg                 io_in_c_bypass_regNext_29_0_is_stationary_7;
  reg        [15:0]   io_in_c_bypass_regNext_29_1_data_7;
  reg                 io_in_c_bypass_regNext_29_1_is_stationary_7;
  reg        [15:0]   io_in_c_bypass_regNext_29_2_data_7;
  reg                 io_in_c_bypass_regNext_29_2_is_stationary_7;
  reg        [15:0]   io_in_c_bypass_regNext_29_3_data_7;
  reg                 io_in_c_bypass_regNext_29_3_is_stationary_7;
  reg        [15:0]   io_in_c_bypass_regNext_30_0_data_7;
  reg                 io_in_c_bypass_regNext_30_0_is_stationary_7;
  reg        [15:0]   io_in_c_bypass_regNext_30_1_data_7;
  reg                 io_in_c_bypass_regNext_30_1_is_stationary_7;
  reg        [15:0]   io_in_c_bypass_regNext_30_2_data_7;
  reg                 io_in_c_bypass_regNext_30_2_is_stationary_7;
  reg        [15:0]   io_in_c_bypass_regNext_30_3_data_7;
  reg                 io_in_c_bypass_regNext_30_3_is_stationary_7;
  reg        [15:0]   io_in_c_bypass_regNext_31_0_data_7;
  reg                 io_in_c_bypass_regNext_31_0_is_stationary_7;
  reg        [15:0]   io_in_c_bypass_regNext_31_1_data_7;
  reg                 io_in_c_bypass_regNext_31_1_is_stationary_7;
  reg        [15:0]   io_in_c_bypass_regNext_31_2_data_7;
  reg                 io_in_c_bypass_regNext_31_2_is_stationary_7;
  reg        [15:0]   io_in_c_bypass_regNext_31_3_data_7;
  reg                 io_in_c_bypass_regNext_31_3_is_stationary_7;
  reg        [15:0]   io_in_c_bypass_regNext_0_0_data_8;
  reg                 io_in_c_bypass_regNext_0_0_is_stationary_8;
  reg        [15:0]   io_in_c_bypass_regNext_0_1_data_8;
  reg                 io_in_c_bypass_regNext_0_1_is_stationary_8;
  reg        [15:0]   io_in_c_bypass_regNext_0_2_data_8;
  reg                 io_in_c_bypass_regNext_0_2_is_stationary_8;
  reg        [15:0]   io_in_c_bypass_regNext_0_3_data_8;
  reg                 io_in_c_bypass_regNext_0_3_is_stationary_8;
  reg        [15:0]   io_in_c_bypass_regNext_1_0_data_8;
  reg                 io_in_c_bypass_regNext_1_0_is_stationary_8;
  reg        [15:0]   io_in_c_bypass_regNext_1_1_data_8;
  reg                 io_in_c_bypass_regNext_1_1_is_stationary_8;
  reg        [15:0]   io_in_c_bypass_regNext_1_2_data_8;
  reg                 io_in_c_bypass_regNext_1_2_is_stationary_8;
  reg        [15:0]   io_in_c_bypass_regNext_1_3_data_8;
  reg                 io_in_c_bypass_regNext_1_3_is_stationary_8;
  reg        [15:0]   io_in_c_bypass_regNext_2_0_data_8;
  reg                 io_in_c_bypass_regNext_2_0_is_stationary_8;
  reg        [15:0]   io_in_c_bypass_regNext_2_1_data_8;
  reg                 io_in_c_bypass_regNext_2_1_is_stationary_8;
  reg        [15:0]   io_in_c_bypass_regNext_2_2_data_8;
  reg                 io_in_c_bypass_regNext_2_2_is_stationary_8;
  reg        [15:0]   io_in_c_bypass_regNext_2_3_data_8;
  reg                 io_in_c_bypass_regNext_2_3_is_stationary_8;
  reg        [15:0]   io_in_c_bypass_regNext_3_0_data_8;
  reg                 io_in_c_bypass_regNext_3_0_is_stationary_8;
  reg        [15:0]   io_in_c_bypass_regNext_3_1_data_8;
  reg                 io_in_c_bypass_regNext_3_1_is_stationary_8;
  reg        [15:0]   io_in_c_bypass_regNext_3_2_data_8;
  reg                 io_in_c_bypass_regNext_3_2_is_stationary_8;
  reg        [15:0]   io_in_c_bypass_regNext_3_3_data_8;
  reg                 io_in_c_bypass_regNext_3_3_is_stationary_8;
  reg        [15:0]   io_in_c_bypass_regNext_4_0_data_8;
  reg                 io_in_c_bypass_regNext_4_0_is_stationary_8;
  reg        [15:0]   io_in_c_bypass_regNext_4_1_data_8;
  reg                 io_in_c_bypass_regNext_4_1_is_stationary_8;
  reg        [15:0]   io_in_c_bypass_regNext_4_2_data_8;
  reg                 io_in_c_bypass_regNext_4_2_is_stationary_8;
  reg        [15:0]   io_in_c_bypass_regNext_4_3_data_8;
  reg                 io_in_c_bypass_regNext_4_3_is_stationary_8;
  reg        [15:0]   io_in_c_bypass_regNext_5_0_data_8;
  reg                 io_in_c_bypass_regNext_5_0_is_stationary_8;
  reg        [15:0]   io_in_c_bypass_regNext_5_1_data_8;
  reg                 io_in_c_bypass_regNext_5_1_is_stationary_8;
  reg        [15:0]   io_in_c_bypass_regNext_5_2_data_8;
  reg                 io_in_c_bypass_regNext_5_2_is_stationary_8;
  reg        [15:0]   io_in_c_bypass_regNext_5_3_data_8;
  reg                 io_in_c_bypass_regNext_5_3_is_stationary_8;
  reg        [15:0]   io_in_c_bypass_regNext_6_0_data_8;
  reg                 io_in_c_bypass_regNext_6_0_is_stationary_8;
  reg        [15:0]   io_in_c_bypass_regNext_6_1_data_8;
  reg                 io_in_c_bypass_regNext_6_1_is_stationary_8;
  reg        [15:0]   io_in_c_bypass_regNext_6_2_data_8;
  reg                 io_in_c_bypass_regNext_6_2_is_stationary_8;
  reg        [15:0]   io_in_c_bypass_regNext_6_3_data_8;
  reg                 io_in_c_bypass_regNext_6_3_is_stationary_8;
  reg        [15:0]   io_in_c_bypass_regNext_7_0_data_8;
  reg                 io_in_c_bypass_regNext_7_0_is_stationary_8;
  reg        [15:0]   io_in_c_bypass_regNext_7_1_data_8;
  reg                 io_in_c_bypass_regNext_7_1_is_stationary_8;
  reg        [15:0]   io_in_c_bypass_regNext_7_2_data_8;
  reg                 io_in_c_bypass_regNext_7_2_is_stationary_8;
  reg        [15:0]   io_in_c_bypass_regNext_7_3_data_8;
  reg                 io_in_c_bypass_regNext_7_3_is_stationary_8;
  reg        [15:0]   io_in_c_bypass_regNext_8_0_data_8;
  reg                 io_in_c_bypass_regNext_8_0_is_stationary_8;
  reg        [15:0]   io_in_c_bypass_regNext_8_1_data_8;
  reg                 io_in_c_bypass_regNext_8_1_is_stationary_8;
  reg        [15:0]   io_in_c_bypass_regNext_8_2_data_8;
  reg                 io_in_c_bypass_regNext_8_2_is_stationary_8;
  reg        [15:0]   io_in_c_bypass_regNext_8_3_data_8;
  reg                 io_in_c_bypass_regNext_8_3_is_stationary_8;
  reg        [15:0]   io_in_c_bypass_regNext_9_0_data_8;
  reg                 io_in_c_bypass_regNext_9_0_is_stationary_8;
  reg        [15:0]   io_in_c_bypass_regNext_9_1_data_8;
  reg                 io_in_c_bypass_regNext_9_1_is_stationary_8;
  reg        [15:0]   io_in_c_bypass_regNext_9_2_data_8;
  reg                 io_in_c_bypass_regNext_9_2_is_stationary_8;
  reg        [15:0]   io_in_c_bypass_regNext_9_3_data_8;
  reg                 io_in_c_bypass_regNext_9_3_is_stationary_8;
  reg        [15:0]   io_in_c_bypass_regNext_10_0_data_8;
  reg                 io_in_c_bypass_regNext_10_0_is_stationary_8;
  reg        [15:0]   io_in_c_bypass_regNext_10_1_data_8;
  reg                 io_in_c_bypass_regNext_10_1_is_stationary_8;
  reg        [15:0]   io_in_c_bypass_regNext_10_2_data_8;
  reg                 io_in_c_bypass_regNext_10_2_is_stationary_8;
  reg        [15:0]   io_in_c_bypass_regNext_10_3_data_8;
  reg                 io_in_c_bypass_regNext_10_3_is_stationary_8;
  reg        [15:0]   io_in_c_bypass_regNext_11_0_data_8;
  reg                 io_in_c_bypass_regNext_11_0_is_stationary_8;
  reg        [15:0]   io_in_c_bypass_regNext_11_1_data_8;
  reg                 io_in_c_bypass_regNext_11_1_is_stationary_8;
  reg        [15:0]   io_in_c_bypass_regNext_11_2_data_8;
  reg                 io_in_c_bypass_regNext_11_2_is_stationary_8;
  reg        [15:0]   io_in_c_bypass_regNext_11_3_data_8;
  reg                 io_in_c_bypass_regNext_11_3_is_stationary_8;
  reg        [15:0]   io_in_c_bypass_regNext_12_0_data_8;
  reg                 io_in_c_bypass_regNext_12_0_is_stationary_8;
  reg        [15:0]   io_in_c_bypass_regNext_12_1_data_8;
  reg                 io_in_c_bypass_regNext_12_1_is_stationary_8;
  reg        [15:0]   io_in_c_bypass_regNext_12_2_data_8;
  reg                 io_in_c_bypass_regNext_12_2_is_stationary_8;
  reg        [15:0]   io_in_c_bypass_regNext_12_3_data_8;
  reg                 io_in_c_bypass_regNext_12_3_is_stationary_8;
  reg        [15:0]   io_in_c_bypass_regNext_13_0_data_8;
  reg                 io_in_c_bypass_regNext_13_0_is_stationary_8;
  reg        [15:0]   io_in_c_bypass_regNext_13_1_data_8;
  reg                 io_in_c_bypass_regNext_13_1_is_stationary_8;
  reg        [15:0]   io_in_c_bypass_regNext_13_2_data_8;
  reg                 io_in_c_bypass_regNext_13_2_is_stationary_8;
  reg        [15:0]   io_in_c_bypass_regNext_13_3_data_8;
  reg                 io_in_c_bypass_regNext_13_3_is_stationary_8;
  reg        [15:0]   io_in_c_bypass_regNext_14_0_data_8;
  reg                 io_in_c_bypass_regNext_14_0_is_stationary_8;
  reg        [15:0]   io_in_c_bypass_regNext_14_1_data_8;
  reg                 io_in_c_bypass_regNext_14_1_is_stationary_8;
  reg        [15:0]   io_in_c_bypass_regNext_14_2_data_8;
  reg                 io_in_c_bypass_regNext_14_2_is_stationary_8;
  reg        [15:0]   io_in_c_bypass_regNext_14_3_data_8;
  reg                 io_in_c_bypass_regNext_14_3_is_stationary_8;
  reg        [15:0]   io_in_c_bypass_regNext_15_0_data_8;
  reg                 io_in_c_bypass_regNext_15_0_is_stationary_8;
  reg        [15:0]   io_in_c_bypass_regNext_15_1_data_8;
  reg                 io_in_c_bypass_regNext_15_1_is_stationary_8;
  reg        [15:0]   io_in_c_bypass_regNext_15_2_data_8;
  reg                 io_in_c_bypass_regNext_15_2_is_stationary_8;
  reg        [15:0]   io_in_c_bypass_regNext_15_3_data_8;
  reg                 io_in_c_bypass_regNext_15_3_is_stationary_8;
  reg        [15:0]   io_in_c_bypass_regNext_16_0_data_8;
  reg                 io_in_c_bypass_regNext_16_0_is_stationary_8;
  reg        [15:0]   io_in_c_bypass_regNext_16_1_data_8;
  reg                 io_in_c_bypass_regNext_16_1_is_stationary_8;
  reg        [15:0]   io_in_c_bypass_regNext_16_2_data_8;
  reg                 io_in_c_bypass_regNext_16_2_is_stationary_8;
  reg        [15:0]   io_in_c_bypass_regNext_16_3_data_8;
  reg                 io_in_c_bypass_regNext_16_3_is_stationary_8;
  reg        [15:0]   io_in_c_bypass_regNext_17_0_data_8;
  reg                 io_in_c_bypass_regNext_17_0_is_stationary_8;
  reg        [15:0]   io_in_c_bypass_regNext_17_1_data_8;
  reg                 io_in_c_bypass_regNext_17_1_is_stationary_8;
  reg        [15:0]   io_in_c_bypass_regNext_17_2_data_8;
  reg                 io_in_c_bypass_regNext_17_2_is_stationary_8;
  reg        [15:0]   io_in_c_bypass_regNext_17_3_data_8;
  reg                 io_in_c_bypass_regNext_17_3_is_stationary_8;
  reg        [15:0]   io_in_c_bypass_regNext_18_0_data_8;
  reg                 io_in_c_bypass_regNext_18_0_is_stationary_8;
  reg        [15:0]   io_in_c_bypass_regNext_18_1_data_8;
  reg                 io_in_c_bypass_regNext_18_1_is_stationary_8;
  reg        [15:0]   io_in_c_bypass_regNext_18_2_data_8;
  reg                 io_in_c_bypass_regNext_18_2_is_stationary_8;
  reg        [15:0]   io_in_c_bypass_regNext_18_3_data_8;
  reg                 io_in_c_bypass_regNext_18_3_is_stationary_8;
  reg        [15:0]   io_in_c_bypass_regNext_19_0_data_8;
  reg                 io_in_c_bypass_regNext_19_0_is_stationary_8;
  reg        [15:0]   io_in_c_bypass_regNext_19_1_data_8;
  reg                 io_in_c_bypass_regNext_19_1_is_stationary_8;
  reg        [15:0]   io_in_c_bypass_regNext_19_2_data_8;
  reg                 io_in_c_bypass_regNext_19_2_is_stationary_8;
  reg        [15:0]   io_in_c_bypass_regNext_19_3_data_8;
  reg                 io_in_c_bypass_regNext_19_3_is_stationary_8;
  reg        [15:0]   io_in_c_bypass_regNext_20_0_data_8;
  reg                 io_in_c_bypass_regNext_20_0_is_stationary_8;
  reg        [15:0]   io_in_c_bypass_regNext_20_1_data_8;
  reg                 io_in_c_bypass_regNext_20_1_is_stationary_8;
  reg        [15:0]   io_in_c_bypass_regNext_20_2_data_8;
  reg                 io_in_c_bypass_regNext_20_2_is_stationary_8;
  reg        [15:0]   io_in_c_bypass_regNext_20_3_data_8;
  reg                 io_in_c_bypass_regNext_20_3_is_stationary_8;
  reg        [15:0]   io_in_c_bypass_regNext_21_0_data_8;
  reg                 io_in_c_bypass_regNext_21_0_is_stationary_8;
  reg        [15:0]   io_in_c_bypass_regNext_21_1_data_8;
  reg                 io_in_c_bypass_regNext_21_1_is_stationary_8;
  reg        [15:0]   io_in_c_bypass_regNext_21_2_data_8;
  reg                 io_in_c_bypass_regNext_21_2_is_stationary_8;
  reg        [15:0]   io_in_c_bypass_regNext_21_3_data_8;
  reg                 io_in_c_bypass_regNext_21_3_is_stationary_8;
  reg        [15:0]   io_in_c_bypass_regNext_22_0_data_8;
  reg                 io_in_c_bypass_regNext_22_0_is_stationary_8;
  reg        [15:0]   io_in_c_bypass_regNext_22_1_data_8;
  reg                 io_in_c_bypass_regNext_22_1_is_stationary_8;
  reg        [15:0]   io_in_c_bypass_regNext_22_2_data_8;
  reg                 io_in_c_bypass_regNext_22_2_is_stationary_8;
  reg        [15:0]   io_in_c_bypass_regNext_22_3_data_8;
  reg                 io_in_c_bypass_regNext_22_3_is_stationary_8;
  reg        [15:0]   io_in_c_bypass_regNext_23_0_data_8;
  reg                 io_in_c_bypass_regNext_23_0_is_stationary_8;
  reg        [15:0]   io_in_c_bypass_regNext_23_1_data_8;
  reg                 io_in_c_bypass_regNext_23_1_is_stationary_8;
  reg        [15:0]   io_in_c_bypass_regNext_23_2_data_8;
  reg                 io_in_c_bypass_regNext_23_2_is_stationary_8;
  reg        [15:0]   io_in_c_bypass_regNext_23_3_data_8;
  reg                 io_in_c_bypass_regNext_23_3_is_stationary_8;
  reg        [15:0]   io_in_c_bypass_regNext_24_0_data_8;
  reg                 io_in_c_bypass_regNext_24_0_is_stationary_8;
  reg        [15:0]   io_in_c_bypass_regNext_24_1_data_8;
  reg                 io_in_c_bypass_regNext_24_1_is_stationary_8;
  reg        [15:0]   io_in_c_bypass_regNext_24_2_data_8;
  reg                 io_in_c_bypass_regNext_24_2_is_stationary_8;
  reg        [15:0]   io_in_c_bypass_regNext_24_3_data_8;
  reg                 io_in_c_bypass_regNext_24_3_is_stationary_8;
  reg        [15:0]   io_in_c_bypass_regNext_25_0_data_8;
  reg                 io_in_c_bypass_regNext_25_0_is_stationary_8;
  reg        [15:0]   io_in_c_bypass_regNext_25_1_data_8;
  reg                 io_in_c_bypass_regNext_25_1_is_stationary_8;
  reg        [15:0]   io_in_c_bypass_regNext_25_2_data_8;
  reg                 io_in_c_bypass_regNext_25_2_is_stationary_8;
  reg        [15:0]   io_in_c_bypass_regNext_25_3_data_8;
  reg                 io_in_c_bypass_regNext_25_3_is_stationary_8;
  reg        [15:0]   io_in_c_bypass_regNext_26_0_data_8;
  reg                 io_in_c_bypass_regNext_26_0_is_stationary_8;
  reg        [15:0]   io_in_c_bypass_regNext_26_1_data_8;
  reg                 io_in_c_bypass_regNext_26_1_is_stationary_8;
  reg        [15:0]   io_in_c_bypass_regNext_26_2_data_8;
  reg                 io_in_c_bypass_regNext_26_2_is_stationary_8;
  reg        [15:0]   io_in_c_bypass_regNext_26_3_data_8;
  reg                 io_in_c_bypass_regNext_26_3_is_stationary_8;
  reg        [15:0]   io_in_c_bypass_regNext_27_0_data_8;
  reg                 io_in_c_bypass_regNext_27_0_is_stationary_8;
  reg        [15:0]   io_in_c_bypass_regNext_27_1_data_8;
  reg                 io_in_c_bypass_regNext_27_1_is_stationary_8;
  reg        [15:0]   io_in_c_bypass_regNext_27_2_data_8;
  reg                 io_in_c_bypass_regNext_27_2_is_stationary_8;
  reg        [15:0]   io_in_c_bypass_regNext_27_3_data_8;
  reg                 io_in_c_bypass_regNext_27_3_is_stationary_8;
  reg        [15:0]   io_in_c_bypass_regNext_28_0_data_8;
  reg                 io_in_c_bypass_regNext_28_0_is_stationary_8;
  reg        [15:0]   io_in_c_bypass_regNext_28_1_data_8;
  reg                 io_in_c_bypass_regNext_28_1_is_stationary_8;
  reg        [15:0]   io_in_c_bypass_regNext_28_2_data_8;
  reg                 io_in_c_bypass_regNext_28_2_is_stationary_8;
  reg        [15:0]   io_in_c_bypass_regNext_28_3_data_8;
  reg                 io_in_c_bypass_regNext_28_3_is_stationary_8;
  reg        [15:0]   io_in_c_bypass_regNext_29_0_data_8;
  reg                 io_in_c_bypass_regNext_29_0_is_stationary_8;
  reg        [15:0]   io_in_c_bypass_regNext_29_1_data_8;
  reg                 io_in_c_bypass_regNext_29_1_is_stationary_8;
  reg        [15:0]   io_in_c_bypass_regNext_29_2_data_8;
  reg                 io_in_c_bypass_regNext_29_2_is_stationary_8;
  reg        [15:0]   io_in_c_bypass_regNext_29_3_data_8;
  reg                 io_in_c_bypass_regNext_29_3_is_stationary_8;
  reg        [15:0]   io_in_c_bypass_regNext_30_0_data_8;
  reg                 io_in_c_bypass_regNext_30_0_is_stationary_8;
  reg        [15:0]   io_in_c_bypass_regNext_30_1_data_8;
  reg                 io_in_c_bypass_regNext_30_1_is_stationary_8;
  reg        [15:0]   io_in_c_bypass_regNext_30_2_data_8;
  reg                 io_in_c_bypass_regNext_30_2_is_stationary_8;
  reg        [15:0]   io_in_c_bypass_regNext_30_3_data_8;
  reg                 io_in_c_bypass_regNext_30_3_is_stationary_8;
  reg        [15:0]   io_in_c_bypass_regNext_31_0_data_8;
  reg                 io_in_c_bypass_regNext_31_0_is_stationary_8;
  reg        [15:0]   io_in_c_bypass_regNext_31_1_data_8;
  reg                 io_in_c_bypass_regNext_31_1_is_stationary_8;
  reg        [15:0]   io_in_c_bypass_regNext_31_2_data_8;
  reg                 io_in_c_bypass_regNext_31_2_is_stationary_8;
  reg        [15:0]   io_in_c_bypass_regNext_31_3_data_8;
  reg                 io_in_c_bypass_regNext_31_3_is_stationary_8;
  reg        [15:0]   io_in_c_bypass_regNext_0_0_data_9;
  reg                 io_in_c_bypass_regNext_0_0_is_stationary_9;
  reg        [15:0]   io_in_c_bypass_regNext_0_1_data_9;
  reg                 io_in_c_bypass_regNext_0_1_is_stationary_9;
  reg        [15:0]   io_in_c_bypass_regNext_0_2_data_9;
  reg                 io_in_c_bypass_regNext_0_2_is_stationary_9;
  reg        [15:0]   io_in_c_bypass_regNext_0_3_data_9;
  reg                 io_in_c_bypass_regNext_0_3_is_stationary_9;
  reg        [15:0]   io_in_c_bypass_regNext_1_0_data_9;
  reg                 io_in_c_bypass_regNext_1_0_is_stationary_9;
  reg        [15:0]   io_in_c_bypass_regNext_1_1_data_9;
  reg                 io_in_c_bypass_regNext_1_1_is_stationary_9;
  reg        [15:0]   io_in_c_bypass_regNext_1_2_data_9;
  reg                 io_in_c_bypass_regNext_1_2_is_stationary_9;
  reg        [15:0]   io_in_c_bypass_regNext_1_3_data_9;
  reg                 io_in_c_bypass_regNext_1_3_is_stationary_9;
  reg        [15:0]   io_in_c_bypass_regNext_2_0_data_9;
  reg                 io_in_c_bypass_regNext_2_0_is_stationary_9;
  reg        [15:0]   io_in_c_bypass_regNext_2_1_data_9;
  reg                 io_in_c_bypass_regNext_2_1_is_stationary_9;
  reg        [15:0]   io_in_c_bypass_regNext_2_2_data_9;
  reg                 io_in_c_bypass_regNext_2_2_is_stationary_9;
  reg        [15:0]   io_in_c_bypass_regNext_2_3_data_9;
  reg                 io_in_c_bypass_regNext_2_3_is_stationary_9;
  reg        [15:0]   io_in_c_bypass_regNext_3_0_data_9;
  reg                 io_in_c_bypass_regNext_3_0_is_stationary_9;
  reg        [15:0]   io_in_c_bypass_regNext_3_1_data_9;
  reg                 io_in_c_bypass_regNext_3_1_is_stationary_9;
  reg        [15:0]   io_in_c_bypass_regNext_3_2_data_9;
  reg                 io_in_c_bypass_regNext_3_2_is_stationary_9;
  reg        [15:0]   io_in_c_bypass_regNext_3_3_data_9;
  reg                 io_in_c_bypass_regNext_3_3_is_stationary_9;
  reg        [15:0]   io_in_c_bypass_regNext_4_0_data_9;
  reg                 io_in_c_bypass_regNext_4_0_is_stationary_9;
  reg        [15:0]   io_in_c_bypass_regNext_4_1_data_9;
  reg                 io_in_c_bypass_regNext_4_1_is_stationary_9;
  reg        [15:0]   io_in_c_bypass_regNext_4_2_data_9;
  reg                 io_in_c_bypass_regNext_4_2_is_stationary_9;
  reg        [15:0]   io_in_c_bypass_regNext_4_3_data_9;
  reg                 io_in_c_bypass_regNext_4_3_is_stationary_9;
  reg        [15:0]   io_in_c_bypass_regNext_5_0_data_9;
  reg                 io_in_c_bypass_regNext_5_0_is_stationary_9;
  reg        [15:0]   io_in_c_bypass_regNext_5_1_data_9;
  reg                 io_in_c_bypass_regNext_5_1_is_stationary_9;
  reg        [15:0]   io_in_c_bypass_regNext_5_2_data_9;
  reg                 io_in_c_bypass_regNext_5_2_is_stationary_9;
  reg        [15:0]   io_in_c_bypass_regNext_5_3_data_9;
  reg                 io_in_c_bypass_regNext_5_3_is_stationary_9;
  reg        [15:0]   io_in_c_bypass_regNext_6_0_data_9;
  reg                 io_in_c_bypass_regNext_6_0_is_stationary_9;
  reg        [15:0]   io_in_c_bypass_regNext_6_1_data_9;
  reg                 io_in_c_bypass_regNext_6_1_is_stationary_9;
  reg        [15:0]   io_in_c_bypass_regNext_6_2_data_9;
  reg                 io_in_c_bypass_regNext_6_2_is_stationary_9;
  reg        [15:0]   io_in_c_bypass_regNext_6_3_data_9;
  reg                 io_in_c_bypass_regNext_6_3_is_stationary_9;
  reg        [15:0]   io_in_c_bypass_regNext_7_0_data_9;
  reg                 io_in_c_bypass_regNext_7_0_is_stationary_9;
  reg        [15:0]   io_in_c_bypass_regNext_7_1_data_9;
  reg                 io_in_c_bypass_regNext_7_1_is_stationary_9;
  reg        [15:0]   io_in_c_bypass_regNext_7_2_data_9;
  reg                 io_in_c_bypass_regNext_7_2_is_stationary_9;
  reg        [15:0]   io_in_c_bypass_regNext_7_3_data_9;
  reg                 io_in_c_bypass_regNext_7_3_is_stationary_9;
  reg        [15:0]   io_in_c_bypass_regNext_8_0_data_9;
  reg                 io_in_c_bypass_regNext_8_0_is_stationary_9;
  reg        [15:0]   io_in_c_bypass_regNext_8_1_data_9;
  reg                 io_in_c_bypass_regNext_8_1_is_stationary_9;
  reg        [15:0]   io_in_c_bypass_regNext_8_2_data_9;
  reg                 io_in_c_bypass_regNext_8_2_is_stationary_9;
  reg        [15:0]   io_in_c_bypass_regNext_8_3_data_9;
  reg                 io_in_c_bypass_regNext_8_3_is_stationary_9;
  reg        [15:0]   io_in_c_bypass_regNext_9_0_data_9;
  reg                 io_in_c_bypass_regNext_9_0_is_stationary_9;
  reg        [15:0]   io_in_c_bypass_regNext_9_1_data_9;
  reg                 io_in_c_bypass_regNext_9_1_is_stationary_9;
  reg        [15:0]   io_in_c_bypass_regNext_9_2_data_9;
  reg                 io_in_c_bypass_regNext_9_2_is_stationary_9;
  reg        [15:0]   io_in_c_bypass_regNext_9_3_data_9;
  reg                 io_in_c_bypass_regNext_9_3_is_stationary_9;
  reg        [15:0]   io_in_c_bypass_regNext_10_0_data_9;
  reg                 io_in_c_bypass_regNext_10_0_is_stationary_9;
  reg        [15:0]   io_in_c_bypass_regNext_10_1_data_9;
  reg                 io_in_c_bypass_regNext_10_1_is_stationary_9;
  reg        [15:0]   io_in_c_bypass_regNext_10_2_data_9;
  reg                 io_in_c_bypass_regNext_10_2_is_stationary_9;
  reg        [15:0]   io_in_c_bypass_regNext_10_3_data_9;
  reg                 io_in_c_bypass_regNext_10_3_is_stationary_9;
  reg        [15:0]   io_in_c_bypass_regNext_11_0_data_9;
  reg                 io_in_c_bypass_regNext_11_0_is_stationary_9;
  reg        [15:0]   io_in_c_bypass_regNext_11_1_data_9;
  reg                 io_in_c_bypass_regNext_11_1_is_stationary_9;
  reg        [15:0]   io_in_c_bypass_regNext_11_2_data_9;
  reg                 io_in_c_bypass_regNext_11_2_is_stationary_9;
  reg        [15:0]   io_in_c_bypass_regNext_11_3_data_9;
  reg                 io_in_c_bypass_regNext_11_3_is_stationary_9;
  reg        [15:0]   io_in_c_bypass_regNext_12_0_data_9;
  reg                 io_in_c_bypass_regNext_12_0_is_stationary_9;
  reg        [15:0]   io_in_c_bypass_regNext_12_1_data_9;
  reg                 io_in_c_bypass_regNext_12_1_is_stationary_9;
  reg        [15:0]   io_in_c_bypass_regNext_12_2_data_9;
  reg                 io_in_c_bypass_regNext_12_2_is_stationary_9;
  reg        [15:0]   io_in_c_bypass_regNext_12_3_data_9;
  reg                 io_in_c_bypass_regNext_12_3_is_stationary_9;
  reg        [15:0]   io_in_c_bypass_regNext_13_0_data_9;
  reg                 io_in_c_bypass_regNext_13_0_is_stationary_9;
  reg        [15:0]   io_in_c_bypass_regNext_13_1_data_9;
  reg                 io_in_c_bypass_regNext_13_1_is_stationary_9;
  reg        [15:0]   io_in_c_bypass_regNext_13_2_data_9;
  reg                 io_in_c_bypass_regNext_13_2_is_stationary_9;
  reg        [15:0]   io_in_c_bypass_regNext_13_3_data_9;
  reg                 io_in_c_bypass_regNext_13_3_is_stationary_9;
  reg        [15:0]   io_in_c_bypass_regNext_14_0_data_9;
  reg                 io_in_c_bypass_regNext_14_0_is_stationary_9;
  reg        [15:0]   io_in_c_bypass_regNext_14_1_data_9;
  reg                 io_in_c_bypass_regNext_14_1_is_stationary_9;
  reg        [15:0]   io_in_c_bypass_regNext_14_2_data_9;
  reg                 io_in_c_bypass_regNext_14_2_is_stationary_9;
  reg        [15:0]   io_in_c_bypass_regNext_14_3_data_9;
  reg                 io_in_c_bypass_regNext_14_3_is_stationary_9;
  reg        [15:0]   io_in_c_bypass_regNext_15_0_data_9;
  reg                 io_in_c_bypass_regNext_15_0_is_stationary_9;
  reg        [15:0]   io_in_c_bypass_regNext_15_1_data_9;
  reg                 io_in_c_bypass_regNext_15_1_is_stationary_9;
  reg        [15:0]   io_in_c_bypass_regNext_15_2_data_9;
  reg                 io_in_c_bypass_regNext_15_2_is_stationary_9;
  reg        [15:0]   io_in_c_bypass_regNext_15_3_data_9;
  reg                 io_in_c_bypass_regNext_15_3_is_stationary_9;
  reg        [15:0]   io_in_c_bypass_regNext_16_0_data_9;
  reg                 io_in_c_bypass_regNext_16_0_is_stationary_9;
  reg        [15:0]   io_in_c_bypass_regNext_16_1_data_9;
  reg                 io_in_c_bypass_regNext_16_1_is_stationary_9;
  reg        [15:0]   io_in_c_bypass_regNext_16_2_data_9;
  reg                 io_in_c_bypass_regNext_16_2_is_stationary_9;
  reg        [15:0]   io_in_c_bypass_regNext_16_3_data_9;
  reg                 io_in_c_bypass_regNext_16_3_is_stationary_9;
  reg        [15:0]   io_in_c_bypass_regNext_17_0_data_9;
  reg                 io_in_c_bypass_regNext_17_0_is_stationary_9;
  reg        [15:0]   io_in_c_bypass_regNext_17_1_data_9;
  reg                 io_in_c_bypass_regNext_17_1_is_stationary_9;
  reg        [15:0]   io_in_c_bypass_regNext_17_2_data_9;
  reg                 io_in_c_bypass_regNext_17_2_is_stationary_9;
  reg        [15:0]   io_in_c_bypass_regNext_17_3_data_9;
  reg                 io_in_c_bypass_regNext_17_3_is_stationary_9;
  reg        [15:0]   io_in_c_bypass_regNext_18_0_data_9;
  reg                 io_in_c_bypass_regNext_18_0_is_stationary_9;
  reg        [15:0]   io_in_c_bypass_regNext_18_1_data_9;
  reg                 io_in_c_bypass_regNext_18_1_is_stationary_9;
  reg        [15:0]   io_in_c_bypass_regNext_18_2_data_9;
  reg                 io_in_c_bypass_regNext_18_2_is_stationary_9;
  reg        [15:0]   io_in_c_bypass_regNext_18_3_data_9;
  reg                 io_in_c_bypass_regNext_18_3_is_stationary_9;
  reg        [15:0]   io_in_c_bypass_regNext_19_0_data_9;
  reg                 io_in_c_bypass_regNext_19_0_is_stationary_9;
  reg        [15:0]   io_in_c_bypass_regNext_19_1_data_9;
  reg                 io_in_c_bypass_regNext_19_1_is_stationary_9;
  reg        [15:0]   io_in_c_bypass_regNext_19_2_data_9;
  reg                 io_in_c_bypass_regNext_19_2_is_stationary_9;
  reg        [15:0]   io_in_c_bypass_regNext_19_3_data_9;
  reg                 io_in_c_bypass_regNext_19_3_is_stationary_9;
  reg        [15:0]   io_in_c_bypass_regNext_20_0_data_9;
  reg                 io_in_c_bypass_regNext_20_0_is_stationary_9;
  reg        [15:0]   io_in_c_bypass_regNext_20_1_data_9;
  reg                 io_in_c_bypass_regNext_20_1_is_stationary_9;
  reg        [15:0]   io_in_c_bypass_regNext_20_2_data_9;
  reg                 io_in_c_bypass_regNext_20_2_is_stationary_9;
  reg        [15:0]   io_in_c_bypass_regNext_20_3_data_9;
  reg                 io_in_c_bypass_regNext_20_3_is_stationary_9;
  reg        [15:0]   io_in_c_bypass_regNext_21_0_data_9;
  reg                 io_in_c_bypass_regNext_21_0_is_stationary_9;
  reg        [15:0]   io_in_c_bypass_regNext_21_1_data_9;
  reg                 io_in_c_bypass_regNext_21_1_is_stationary_9;
  reg        [15:0]   io_in_c_bypass_regNext_21_2_data_9;
  reg                 io_in_c_bypass_regNext_21_2_is_stationary_9;
  reg        [15:0]   io_in_c_bypass_regNext_21_3_data_9;
  reg                 io_in_c_bypass_regNext_21_3_is_stationary_9;
  reg        [15:0]   io_in_c_bypass_regNext_22_0_data_9;
  reg                 io_in_c_bypass_regNext_22_0_is_stationary_9;
  reg        [15:0]   io_in_c_bypass_regNext_22_1_data_9;
  reg                 io_in_c_bypass_regNext_22_1_is_stationary_9;
  reg        [15:0]   io_in_c_bypass_regNext_22_2_data_9;
  reg                 io_in_c_bypass_regNext_22_2_is_stationary_9;
  reg        [15:0]   io_in_c_bypass_regNext_22_3_data_9;
  reg                 io_in_c_bypass_regNext_22_3_is_stationary_9;
  reg        [15:0]   io_in_c_bypass_regNext_23_0_data_9;
  reg                 io_in_c_bypass_regNext_23_0_is_stationary_9;
  reg        [15:0]   io_in_c_bypass_regNext_23_1_data_9;
  reg                 io_in_c_bypass_regNext_23_1_is_stationary_9;
  reg        [15:0]   io_in_c_bypass_regNext_23_2_data_9;
  reg                 io_in_c_bypass_regNext_23_2_is_stationary_9;
  reg        [15:0]   io_in_c_bypass_regNext_23_3_data_9;
  reg                 io_in_c_bypass_regNext_23_3_is_stationary_9;
  reg        [15:0]   io_in_c_bypass_regNext_24_0_data_9;
  reg                 io_in_c_bypass_regNext_24_0_is_stationary_9;
  reg        [15:0]   io_in_c_bypass_regNext_24_1_data_9;
  reg                 io_in_c_bypass_regNext_24_1_is_stationary_9;
  reg        [15:0]   io_in_c_bypass_regNext_24_2_data_9;
  reg                 io_in_c_bypass_regNext_24_2_is_stationary_9;
  reg        [15:0]   io_in_c_bypass_regNext_24_3_data_9;
  reg                 io_in_c_bypass_regNext_24_3_is_stationary_9;
  reg        [15:0]   io_in_c_bypass_regNext_25_0_data_9;
  reg                 io_in_c_bypass_regNext_25_0_is_stationary_9;
  reg        [15:0]   io_in_c_bypass_regNext_25_1_data_9;
  reg                 io_in_c_bypass_regNext_25_1_is_stationary_9;
  reg        [15:0]   io_in_c_bypass_regNext_25_2_data_9;
  reg                 io_in_c_bypass_regNext_25_2_is_stationary_9;
  reg        [15:0]   io_in_c_bypass_regNext_25_3_data_9;
  reg                 io_in_c_bypass_regNext_25_3_is_stationary_9;
  reg        [15:0]   io_in_c_bypass_regNext_26_0_data_9;
  reg                 io_in_c_bypass_regNext_26_0_is_stationary_9;
  reg        [15:0]   io_in_c_bypass_regNext_26_1_data_9;
  reg                 io_in_c_bypass_regNext_26_1_is_stationary_9;
  reg        [15:0]   io_in_c_bypass_regNext_26_2_data_9;
  reg                 io_in_c_bypass_regNext_26_2_is_stationary_9;
  reg        [15:0]   io_in_c_bypass_regNext_26_3_data_9;
  reg                 io_in_c_bypass_regNext_26_3_is_stationary_9;
  reg        [15:0]   io_in_c_bypass_regNext_27_0_data_9;
  reg                 io_in_c_bypass_regNext_27_0_is_stationary_9;
  reg        [15:0]   io_in_c_bypass_regNext_27_1_data_9;
  reg                 io_in_c_bypass_regNext_27_1_is_stationary_9;
  reg        [15:0]   io_in_c_bypass_regNext_27_2_data_9;
  reg                 io_in_c_bypass_regNext_27_2_is_stationary_9;
  reg        [15:0]   io_in_c_bypass_regNext_27_3_data_9;
  reg                 io_in_c_bypass_regNext_27_3_is_stationary_9;
  reg        [15:0]   io_in_c_bypass_regNext_28_0_data_9;
  reg                 io_in_c_bypass_regNext_28_0_is_stationary_9;
  reg        [15:0]   io_in_c_bypass_regNext_28_1_data_9;
  reg                 io_in_c_bypass_regNext_28_1_is_stationary_9;
  reg        [15:0]   io_in_c_bypass_regNext_28_2_data_9;
  reg                 io_in_c_bypass_regNext_28_2_is_stationary_9;
  reg        [15:0]   io_in_c_bypass_regNext_28_3_data_9;
  reg                 io_in_c_bypass_regNext_28_3_is_stationary_9;
  reg        [15:0]   io_in_c_bypass_regNext_29_0_data_9;
  reg                 io_in_c_bypass_regNext_29_0_is_stationary_9;
  reg        [15:0]   io_in_c_bypass_regNext_29_1_data_9;
  reg                 io_in_c_bypass_regNext_29_1_is_stationary_9;
  reg        [15:0]   io_in_c_bypass_regNext_29_2_data_9;
  reg                 io_in_c_bypass_regNext_29_2_is_stationary_9;
  reg        [15:0]   io_in_c_bypass_regNext_29_3_data_9;
  reg                 io_in_c_bypass_regNext_29_3_is_stationary_9;
  reg        [15:0]   io_in_c_bypass_regNext_30_0_data_9;
  reg                 io_in_c_bypass_regNext_30_0_is_stationary_9;
  reg        [15:0]   io_in_c_bypass_regNext_30_1_data_9;
  reg                 io_in_c_bypass_regNext_30_1_is_stationary_9;
  reg        [15:0]   io_in_c_bypass_regNext_30_2_data_9;
  reg                 io_in_c_bypass_regNext_30_2_is_stationary_9;
  reg        [15:0]   io_in_c_bypass_regNext_30_3_data_9;
  reg                 io_in_c_bypass_regNext_30_3_is_stationary_9;
  reg        [15:0]   io_in_c_bypass_regNext_31_0_data_9;
  reg                 io_in_c_bypass_regNext_31_0_is_stationary_9;
  reg        [15:0]   io_in_c_bypass_regNext_31_1_data_9;
  reg                 io_in_c_bypass_regNext_31_1_is_stationary_9;
  reg        [15:0]   io_in_c_bypass_regNext_31_2_data_9;
  reg                 io_in_c_bypass_regNext_31_2_is_stationary_9;
  reg        [15:0]   io_in_c_bypass_regNext_31_3_data_9;
  reg                 io_in_c_bypass_regNext_31_3_is_stationary_9;
  reg        [15:0]   io_in_c_bypass_regNext_0_0_data_10;
  reg                 io_in_c_bypass_regNext_0_0_is_stationary_10;
  reg        [15:0]   io_in_c_bypass_regNext_0_1_data_10;
  reg                 io_in_c_bypass_regNext_0_1_is_stationary_10;
  reg        [15:0]   io_in_c_bypass_regNext_0_2_data_10;
  reg                 io_in_c_bypass_regNext_0_2_is_stationary_10;
  reg        [15:0]   io_in_c_bypass_regNext_0_3_data_10;
  reg                 io_in_c_bypass_regNext_0_3_is_stationary_10;
  reg        [15:0]   io_in_c_bypass_regNext_1_0_data_10;
  reg                 io_in_c_bypass_regNext_1_0_is_stationary_10;
  reg        [15:0]   io_in_c_bypass_regNext_1_1_data_10;
  reg                 io_in_c_bypass_regNext_1_1_is_stationary_10;
  reg        [15:0]   io_in_c_bypass_regNext_1_2_data_10;
  reg                 io_in_c_bypass_regNext_1_2_is_stationary_10;
  reg        [15:0]   io_in_c_bypass_regNext_1_3_data_10;
  reg                 io_in_c_bypass_regNext_1_3_is_stationary_10;
  reg        [15:0]   io_in_c_bypass_regNext_2_0_data_10;
  reg                 io_in_c_bypass_regNext_2_0_is_stationary_10;
  reg        [15:0]   io_in_c_bypass_regNext_2_1_data_10;
  reg                 io_in_c_bypass_regNext_2_1_is_stationary_10;
  reg        [15:0]   io_in_c_bypass_regNext_2_2_data_10;
  reg                 io_in_c_bypass_regNext_2_2_is_stationary_10;
  reg        [15:0]   io_in_c_bypass_regNext_2_3_data_10;
  reg                 io_in_c_bypass_regNext_2_3_is_stationary_10;
  reg        [15:0]   io_in_c_bypass_regNext_3_0_data_10;
  reg                 io_in_c_bypass_regNext_3_0_is_stationary_10;
  reg        [15:0]   io_in_c_bypass_regNext_3_1_data_10;
  reg                 io_in_c_bypass_regNext_3_1_is_stationary_10;
  reg        [15:0]   io_in_c_bypass_regNext_3_2_data_10;
  reg                 io_in_c_bypass_regNext_3_2_is_stationary_10;
  reg        [15:0]   io_in_c_bypass_regNext_3_3_data_10;
  reg                 io_in_c_bypass_regNext_3_3_is_stationary_10;
  reg        [15:0]   io_in_c_bypass_regNext_4_0_data_10;
  reg                 io_in_c_bypass_regNext_4_0_is_stationary_10;
  reg        [15:0]   io_in_c_bypass_regNext_4_1_data_10;
  reg                 io_in_c_bypass_regNext_4_1_is_stationary_10;
  reg        [15:0]   io_in_c_bypass_regNext_4_2_data_10;
  reg                 io_in_c_bypass_regNext_4_2_is_stationary_10;
  reg        [15:0]   io_in_c_bypass_regNext_4_3_data_10;
  reg                 io_in_c_bypass_regNext_4_3_is_stationary_10;
  reg        [15:0]   io_in_c_bypass_regNext_5_0_data_10;
  reg                 io_in_c_bypass_regNext_5_0_is_stationary_10;
  reg        [15:0]   io_in_c_bypass_regNext_5_1_data_10;
  reg                 io_in_c_bypass_regNext_5_1_is_stationary_10;
  reg        [15:0]   io_in_c_bypass_regNext_5_2_data_10;
  reg                 io_in_c_bypass_regNext_5_2_is_stationary_10;
  reg        [15:0]   io_in_c_bypass_regNext_5_3_data_10;
  reg                 io_in_c_bypass_regNext_5_3_is_stationary_10;
  reg        [15:0]   io_in_c_bypass_regNext_6_0_data_10;
  reg                 io_in_c_bypass_regNext_6_0_is_stationary_10;
  reg        [15:0]   io_in_c_bypass_regNext_6_1_data_10;
  reg                 io_in_c_bypass_regNext_6_1_is_stationary_10;
  reg        [15:0]   io_in_c_bypass_regNext_6_2_data_10;
  reg                 io_in_c_bypass_regNext_6_2_is_stationary_10;
  reg        [15:0]   io_in_c_bypass_regNext_6_3_data_10;
  reg                 io_in_c_bypass_regNext_6_3_is_stationary_10;
  reg        [15:0]   io_in_c_bypass_regNext_7_0_data_10;
  reg                 io_in_c_bypass_regNext_7_0_is_stationary_10;
  reg        [15:0]   io_in_c_bypass_regNext_7_1_data_10;
  reg                 io_in_c_bypass_regNext_7_1_is_stationary_10;
  reg        [15:0]   io_in_c_bypass_regNext_7_2_data_10;
  reg                 io_in_c_bypass_regNext_7_2_is_stationary_10;
  reg        [15:0]   io_in_c_bypass_regNext_7_3_data_10;
  reg                 io_in_c_bypass_regNext_7_3_is_stationary_10;
  reg        [15:0]   io_in_c_bypass_regNext_8_0_data_10;
  reg                 io_in_c_bypass_regNext_8_0_is_stationary_10;
  reg        [15:0]   io_in_c_bypass_regNext_8_1_data_10;
  reg                 io_in_c_bypass_regNext_8_1_is_stationary_10;
  reg        [15:0]   io_in_c_bypass_regNext_8_2_data_10;
  reg                 io_in_c_bypass_regNext_8_2_is_stationary_10;
  reg        [15:0]   io_in_c_bypass_regNext_8_3_data_10;
  reg                 io_in_c_bypass_regNext_8_3_is_stationary_10;
  reg        [15:0]   io_in_c_bypass_regNext_9_0_data_10;
  reg                 io_in_c_bypass_regNext_9_0_is_stationary_10;
  reg        [15:0]   io_in_c_bypass_regNext_9_1_data_10;
  reg                 io_in_c_bypass_regNext_9_1_is_stationary_10;
  reg        [15:0]   io_in_c_bypass_regNext_9_2_data_10;
  reg                 io_in_c_bypass_regNext_9_2_is_stationary_10;
  reg        [15:0]   io_in_c_bypass_regNext_9_3_data_10;
  reg                 io_in_c_bypass_regNext_9_3_is_stationary_10;
  reg        [15:0]   io_in_c_bypass_regNext_10_0_data_10;
  reg                 io_in_c_bypass_regNext_10_0_is_stationary_10;
  reg        [15:0]   io_in_c_bypass_regNext_10_1_data_10;
  reg                 io_in_c_bypass_regNext_10_1_is_stationary_10;
  reg        [15:0]   io_in_c_bypass_regNext_10_2_data_10;
  reg                 io_in_c_bypass_regNext_10_2_is_stationary_10;
  reg        [15:0]   io_in_c_bypass_regNext_10_3_data_10;
  reg                 io_in_c_bypass_regNext_10_3_is_stationary_10;
  reg        [15:0]   io_in_c_bypass_regNext_11_0_data_10;
  reg                 io_in_c_bypass_regNext_11_0_is_stationary_10;
  reg        [15:0]   io_in_c_bypass_regNext_11_1_data_10;
  reg                 io_in_c_bypass_regNext_11_1_is_stationary_10;
  reg        [15:0]   io_in_c_bypass_regNext_11_2_data_10;
  reg                 io_in_c_bypass_regNext_11_2_is_stationary_10;
  reg        [15:0]   io_in_c_bypass_regNext_11_3_data_10;
  reg                 io_in_c_bypass_regNext_11_3_is_stationary_10;
  reg        [15:0]   io_in_c_bypass_regNext_12_0_data_10;
  reg                 io_in_c_bypass_regNext_12_0_is_stationary_10;
  reg        [15:0]   io_in_c_bypass_regNext_12_1_data_10;
  reg                 io_in_c_bypass_regNext_12_1_is_stationary_10;
  reg        [15:0]   io_in_c_bypass_regNext_12_2_data_10;
  reg                 io_in_c_bypass_regNext_12_2_is_stationary_10;
  reg        [15:0]   io_in_c_bypass_regNext_12_3_data_10;
  reg                 io_in_c_bypass_regNext_12_3_is_stationary_10;
  reg        [15:0]   io_in_c_bypass_regNext_13_0_data_10;
  reg                 io_in_c_bypass_regNext_13_0_is_stationary_10;
  reg        [15:0]   io_in_c_bypass_regNext_13_1_data_10;
  reg                 io_in_c_bypass_regNext_13_1_is_stationary_10;
  reg        [15:0]   io_in_c_bypass_regNext_13_2_data_10;
  reg                 io_in_c_bypass_regNext_13_2_is_stationary_10;
  reg        [15:0]   io_in_c_bypass_regNext_13_3_data_10;
  reg                 io_in_c_bypass_regNext_13_3_is_stationary_10;
  reg        [15:0]   io_in_c_bypass_regNext_14_0_data_10;
  reg                 io_in_c_bypass_regNext_14_0_is_stationary_10;
  reg        [15:0]   io_in_c_bypass_regNext_14_1_data_10;
  reg                 io_in_c_bypass_regNext_14_1_is_stationary_10;
  reg        [15:0]   io_in_c_bypass_regNext_14_2_data_10;
  reg                 io_in_c_bypass_regNext_14_2_is_stationary_10;
  reg        [15:0]   io_in_c_bypass_regNext_14_3_data_10;
  reg                 io_in_c_bypass_regNext_14_3_is_stationary_10;
  reg        [15:0]   io_in_c_bypass_regNext_15_0_data_10;
  reg                 io_in_c_bypass_regNext_15_0_is_stationary_10;
  reg        [15:0]   io_in_c_bypass_regNext_15_1_data_10;
  reg                 io_in_c_bypass_regNext_15_1_is_stationary_10;
  reg        [15:0]   io_in_c_bypass_regNext_15_2_data_10;
  reg                 io_in_c_bypass_regNext_15_2_is_stationary_10;
  reg        [15:0]   io_in_c_bypass_regNext_15_3_data_10;
  reg                 io_in_c_bypass_regNext_15_3_is_stationary_10;
  reg        [15:0]   io_in_c_bypass_regNext_16_0_data_10;
  reg                 io_in_c_bypass_regNext_16_0_is_stationary_10;
  reg        [15:0]   io_in_c_bypass_regNext_16_1_data_10;
  reg                 io_in_c_bypass_regNext_16_1_is_stationary_10;
  reg        [15:0]   io_in_c_bypass_regNext_16_2_data_10;
  reg                 io_in_c_bypass_regNext_16_2_is_stationary_10;
  reg        [15:0]   io_in_c_bypass_regNext_16_3_data_10;
  reg                 io_in_c_bypass_regNext_16_3_is_stationary_10;
  reg        [15:0]   io_in_c_bypass_regNext_17_0_data_10;
  reg                 io_in_c_bypass_regNext_17_0_is_stationary_10;
  reg        [15:0]   io_in_c_bypass_regNext_17_1_data_10;
  reg                 io_in_c_bypass_regNext_17_1_is_stationary_10;
  reg        [15:0]   io_in_c_bypass_regNext_17_2_data_10;
  reg                 io_in_c_bypass_regNext_17_2_is_stationary_10;
  reg        [15:0]   io_in_c_bypass_regNext_17_3_data_10;
  reg                 io_in_c_bypass_regNext_17_3_is_stationary_10;
  reg        [15:0]   io_in_c_bypass_regNext_18_0_data_10;
  reg                 io_in_c_bypass_regNext_18_0_is_stationary_10;
  reg        [15:0]   io_in_c_bypass_regNext_18_1_data_10;
  reg                 io_in_c_bypass_regNext_18_1_is_stationary_10;
  reg        [15:0]   io_in_c_bypass_regNext_18_2_data_10;
  reg                 io_in_c_bypass_regNext_18_2_is_stationary_10;
  reg        [15:0]   io_in_c_bypass_regNext_18_3_data_10;
  reg                 io_in_c_bypass_regNext_18_3_is_stationary_10;
  reg        [15:0]   io_in_c_bypass_regNext_19_0_data_10;
  reg                 io_in_c_bypass_regNext_19_0_is_stationary_10;
  reg        [15:0]   io_in_c_bypass_regNext_19_1_data_10;
  reg                 io_in_c_bypass_regNext_19_1_is_stationary_10;
  reg        [15:0]   io_in_c_bypass_regNext_19_2_data_10;
  reg                 io_in_c_bypass_regNext_19_2_is_stationary_10;
  reg        [15:0]   io_in_c_bypass_regNext_19_3_data_10;
  reg                 io_in_c_bypass_regNext_19_3_is_stationary_10;
  reg        [15:0]   io_in_c_bypass_regNext_20_0_data_10;
  reg                 io_in_c_bypass_regNext_20_0_is_stationary_10;
  reg        [15:0]   io_in_c_bypass_regNext_20_1_data_10;
  reg                 io_in_c_bypass_regNext_20_1_is_stationary_10;
  reg        [15:0]   io_in_c_bypass_regNext_20_2_data_10;
  reg                 io_in_c_bypass_regNext_20_2_is_stationary_10;
  reg        [15:0]   io_in_c_bypass_regNext_20_3_data_10;
  reg                 io_in_c_bypass_regNext_20_3_is_stationary_10;
  reg        [15:0]   io_in_c_bypass_regNext_21_0_data_10;
  reg                 io_in_c_bypass_regNext_21_0_is_stationary_10;
  reg        [15:0]   io_in_c_bypass_regNext_21_1_data_10;
  reg                 io_in_c_bypass_regNext_21_1_is_stationary_10;
  reg        [15:0]   io_in_c_bypass_regNext_21_2_data_10;
  reg                 io_in_c_bypass_regNext_21_2_is_stationary_10;
  reg        [15:0]   io_in_c_bypass_regNext_21_3_data_10;
  reg                 io_in_c_bypass_regNext_21_3_is_stationary_10;
  reg        [15:0]   io_in_c_bypass_regNext_22_0_data_10;
  reg                 io_in_c_bypass_regNext_22_0_is_stationary_10;
  reg        [15:0]   io_in_c_bypass_regNext_22_1_data_10;
  reg                 io_in_c_bypass_regNext_22_1_is_stationary_10;
  reg        [15:0]   io_in_c_bypass_regNext_22_2_data_10;
  reg                 io_in_c_bypass_regNext_22_2_is_stationary_10;
  reg        [15:0]   io_in_c_bypass_regNext_22_3_data_10;
  reg                 io_in_c_bypass_regNext_22_3_is_stationary_10;
  reg        [15:0]   io_in_c_bypass_regNext_23_0_data_10;
  reg                 io_in_c_bypass_regNext_23_0_is_stationary_10;
  reg        [15:0]   io_in_c_bypass_regNext_23_1_data_10;
  reg                 io_in_c_bypass_regNext_23_1_is_stationary_10;
  reg        [15:0]   io_in_c_bypass_regNext_23_2_data_10;
  reg                 io_in_c_bypass_regNext_23_2_is_stationary_10;
  reg        [15:0]   io_in_c_bypass_regNext_23_3_data_10;
  reg                 io_in_c_bypass_regNext_23_3_is_stationary_10;
  reg        [15:0]   io_in_c_bypass_regNext_24_0_data_10;
  reg                 io_in_c_bypass_regNext_24_0_is_stationary_10;
  reg        [15:0]   io_in_c_bypass_regNext_24_1_data_10;
  reg                 io_in_c_bypass_regNext_24_1_is_stationary_10;
  reg        [15:0]   io_in_c_bypass_regNext_24_2_data_10;
  reg                 io_in_c_bypass_regNext_24_2_is_stationary_10;
  reg        [15:0]   io_in_c_bypass_regNext_24_3_data_10;
  reg                 io_in_c_bypass_regNext_24_3_is_stationary_10;
  reg        [15:0]   io_in_c_bypass_regNext_25_0_data_10;
  reg                 io_in_c_bypass_regNext_25_0_is_stationary_10;
  reg        [15:0]   io_in_c_bypass_regNext_25_1_data_10;
  reg                 io_in_c_bypass_regNext_25_1_is_stationary_10;
  reg        [15:0]   io_in_c_bypass_regNext_25_2_data_10;
  reg                 io_in_c_bypass_regNext_25_2_is_stationary_10;
  reg        [15:0]   io_in_c_bypass_regNext_25_3_data_10;
  reg                 io_in_c_bypass_regNext_25_3_is_stationary_10;
  reg        [15:0]   io_in_c_bypass_regNext_26_0_data_10;
  reg                 io_in_c_bypass_regNext_26_0_is_stationary_10;
  reg        [15:0]   io_in_c_bypass_regNext_26_1_data_10;
  reg                 io_in_c_bypass_regNext_26_1_is_stationary_10;
  reg        [15:0]   io_in_c_bypass_regNext_26_2_data_10;
  reg                 io_in_c_bypass_regNext_26_2_is_stationary_10;
  reg        [15:0]   io_in_c_bypass_regNext_26_3_data_10;
  reg                 io_in_c_bypass_regNext_26_3_is_stationary_10;
  reg        [15:0]   io_in_c_bypass_regNext_27_0_data_10;
  reg                 io_in_c_bypass_regNext_27_0_is_stationary_10;
  reg        [15:0]   io_in_c_bypass_regNext_27_1_data_10;
  reg                 io_in_c_bypass_regNext_27_1_is_stationary_10;
  reg        [15:0]   io_in_c_bypass_regNext_27_2_data_10;
  reg                 io_in_c_bypass_regNext_27_2_is_stationary_10;
  reg        [15:0]   io_in_c_bypass_regNext_27_3_data_10;
  reg                 io_in_c_bypass_regNext_27_3_is_stationary_10;
  reg        [15:0]   io_in_c_bypass_regNext_28_0_data_10;
  reg                 io_in_c_bypass_regNext_28_0_is_stationary_10;
  reg        [15:0]   io_in_c_bypass_regNext_28_1_data_10;
  reg                 io_in_c_bypass_regNext_28_1_is_stationary_10;
  reg        [15:0]   io_in_c_bypass_regNext_28_2_data_10;
  reg                 io_in_c_bypass_regNext_28_2_is_stationary_10;
  reg        [15:0]   io_in_c_bypass_regNext_28_3_data_10;
  reg                 io_in_c_bypass_regNext_28_3_is_stationary_10;
  reg        [15:0]   io_in_c_bypass_regNext_29_0_data_10;
  reg                 io_in_c_bypass_regNext_29_0_is_stationary_10;
  reg        [15:0]   io_in_c_bypass_regNext_29_1_data_10;
  reg                 io_in_c_bypass_regNext_29_1_is_stationary_10;
  reg        [15:0]   io_in_c_bypass_regNext_29_2_data_10;
  reg                 io_in_c_bypass_regNext_29_2_is_stationary_10;
  reg        [15:0]   io_in_c_bypass_regNext_29_3_data_10;
  reg                 io_in_c_bypass_regNext_29_3_is_stationary_10;
  reg        [15:0]   io_in_c_bypass_regNext_30_0_data_10;
  reg                 io_in_c_bypass_regNext_30_0_is_stationary_10;
  reg        [15:0]   io_in_c_bypass_regNext_30_1_data_10;
  reg                 io_in_c_bypass_regNext_30_1_is_stationary_10;
  reg        [15:0]   io_in_c_bypass_regNext_30_2_data_10;
  reg                 io_in_c_bypass_regNext_30_2_is_stationary_10;
  reg        [15:0]   io_in_c_bypass_regNext_30_3_data_10;
  reg                 io_in_c_bypass_regNext_30_3_is_stationary_10;
  reg        [15:0]   io_in_c_bypass_regNext_31_0_data_10;
  reg                 io_in_c_bypass_regNext_31_0_is_stationary_10;
  reg        [15:0]   io_in_c_bypass_regNext_31_1_data_10;
  reg                 io_in_c_bypass_regNext_31_1_is_stationary_10;
  reg        [15:0]   io_in_c_bypass_regNext_31_2_data_10;
  reg                 io_in_c_bypass_regNext_31_2_is_stationary_10;
  reg        [15:0]   io_in_c_bypass_regNext_31_3_data_10;
  reg                 io_in_c_bypass_regNext_31_3_is_stationary_10;
  reg        [15:0]   io_in_c_bypass_regNext_0_0_data_11;
  reg                 io_in_c_bypass_regNext_0_0_is_stationary_11;
  reg        [15:0]   io_in_c_bypass_regNext_0_1_data_11;
  reg                 io_in_c_bypass_regNext_0_1_is_stationary_11;
  reg        [15:0]   io_in_c_bypass_regNext_0_2_data_11;
  reg                 io_in_c_bypass_regNext_0_2_is_stationary_11;
  reg        [15:0]   io_in_c_bypass_regNext_0_3_data_11;
  reg                 io_in_c_bypass_regNext_0_3_is_stationary_11;
  reg        [15:0]   io_in_c_bypass_regNext_1_0_data_11;
  reg                 io_in_c_bypass_regNext_1_0_is_stationary_11;
  reg        [15:0]   io_in_c_bypass_regNext_1_1_data_11;
  reg                 io_in_c_bypass_regNext_1_1_is_stationary_11;
  reg        [15:0]   io_in_c_bypass_regNext_1_2_data_11;
  reg                 io_in_c_bypass_regNext_1_2_is_stationary_11;
  reg        [15:0]   io_in_c_bypass_regNext_1_3_data_11;
  reg                 io_in_c_bypass_regNext_1_3_is_stationary_11;
  reg        [15:0]   io_in_c_bypass_regNext_2_0_data_11;
  reg                 io_in_c_bypass_regNext_2_0_is_stationary_11;
  reg        [15:0]   io_in_c_bypass_regNext_2_1_data_11;
  reg                 io_in_c_bypass_regNext_2_1_is_stationary_11;
  reg        [15:0]   io_in_c_bypass_regNext_2_2_data_11;
  reg                 io_in_c_bypass_regNext_2_2_is_stationary_11;
  reg        [15:0]   io_in_c_bypass_regNext_2_3_data_11;
  reg                 io_in_c_bypass_regNext_2_3_is_stationary_11;
  reg        [15:0]   io_in_c_bypass_regNext_3_0_data_11;
  reg                 io_in_c_bypass_regNext_3_0_is_stationary_11;
  reg        [15:0]   io_in_c_bypass_regNext_3_1_data_11;
  reg                 io_in_c_bypass_regNext_3_1_is_stationary_11;
  reg        [15:0]   io_in_c_bypass_regNext_3_2_data_11;
  reg                 io_in_c_bypass_regNext_3_2_is_stationary_11;
  reg        [15:0]   io_in_c_bypass_regNext_3_3_data_11;
  reg                 io_in_c_bypass_regNext_3_3_is_stationary_11;
  reg        [15:0]   io_in_c_bypass_regNext_4_0_data_11;
  reg                 io_in_c_bypass_regNext_4_0_is_stationary_11;
  reg        [15:0]   io_in_c_bypass_regNext_4_1_data_11;
  reg                 io_in_c_bypass_regNext_4_1_is_stationary_11;
  reg        [15:0]   io_in_c_bypass_regNext_4_2_data_11;
  reg                 io_in_c_bypass_regNext_4_2_is_stationary_11;
  reg        [15:0]   io_in_c_bypass_regNext_4_3_data_11;
  reg                 io_in_c_bypass_regNext_4_3_is_stationary_11;
  reg        [15:0]   io_in_c_bypass_regNext_5_0_data_11;
  reg                 io_in_c_bypass_regNext_5_0_is_stationary_11;
  reg        [15:0]   io_in_c_bypass_regNext_5_1_data_11;
  reg                 io_in_c_bypass_regNext_5_1_is_stationary_11;
  reg        [15:0]   io_in_c_bypass_regNext_5_2_data_11;
  reg                 io_in_c_bypass_regNext_5_2_is_stationary_11;
  reg        [15:0]   io_in_c_bypass_regNext_5_3_data_11;
  reg                 io_in_c_bypass_regNext_5_3_is_stationary_11;
  reg        [15:0]   io_in_c_bypass_regNext_6_0_data_11;
  reg                 io_in_c_bypass_regNext_6_0_is_stationary_11;
  reg        [15:0]   io_in_c_bypass_regNext_6_1_data_11;
  reg                 io_in_c_bypass_regNext_6_1_is_stationary_11;
  reg        [15:0]   io_in_c_bypass_regNext_6_2_data_11;
  reg                 io_in_c_bypass_regNext_6_2_is_stationary_11;
  reg        [15:0]   io_in_c_bypass_regNext_6_3_data_11;
  reg                 io_in_c_bypass_regNext_6_3_is_stationary_11;
  reg        [15:0]   io_in_c_bypass_regNext_7_0_data_11;
  reg                 io_in_c_bypass_regNext_7_0_is_stationary_11;
  reg        [15:0]   io_in_c_bypass_regNext_7_1_data_11;
  reg                 io_in_c_bypass_regNext_7_1_is_stationary_11;
  reg        [15:0]   io_in_c_bypass_regNext_7_2_data_11;
  reg                 io_in_c_bypass_regNext_7_2_is_stationary_11;
  reg        [15:0]   io_in_c_bypass_regNext_7_3_data_11;
  reg                 io_in_c_bypass_regNext_7_3_is_stationary_11;
  reg        [15:0]   io_in_c_bypass_regNext_8_0_data_11;
  reg                 io_in_c_bypass_regNext_8_0_is_stationary_11;
  reg        [15:0]   io_in_c_bypass_regNext_8_1_data_11;
  reg                 io_in_c_bypass_regNext_8_1_is_stationary_11;
  reg        [15:0]   io_in_c_bypass_regNext_8_2_data_11;
  reg                 io_in_c_bypass_regNext_8_2_is_stationary_11;
  reg        [15:0]   io_in_c_bypass_regNext_8_3_data_11;
  reg                 io_in_c_bypass_regNext_8_3_is_stationary_11;
  reg        [15:0]   io_in_c_bypass_regNext_9_0_data_11;
  reg                 io_in_c_bypass_regNext_9_0_is_stationary_11;
  reg        [15:0]   io_in_c_bypass_regNext_9_1_data_11;
  reg                 io_in_c_bypass_regNext_9_1_is_stationary_11;
  reg        [15:0]   io_in_c_bypass_regNext_9_2_data_11;
  reg                 io_in_c_bypass_regNext_9_2_is_stationary_11;
  reg        [15:0]   io_in_c_bypass_regNext_9_3_data_11;
  reg                 io_in_c_bypass_regNext_9_3_is_stationary_11;
  reg        [15:0]   io_in_c_bypass_regNext_10_0_data_11;
  reg                 io_in_c_bypass_regNext_10_0_is_stationary_11;
  reg        [15:0]   io_in_c_bypass_regNext_10_1_data_11;
  reg                 io_in_c_bypass_regNext_10_1_is_stationary_11;
  reg        [15:0]   io_in_c_bypass_regNext_10_2_data_11;
  reg                 io_in_c_bypass_regNext_10_2_is_stationary_11;
  reg        [15:0]   io_in_c_bypass_regNext_10_3_data_11;
  reg                 io_in_c_bypass_regNext_10_3_is_stationary_11;
  reg        [15:0]   io_in_c_bypass_regNext_11_0_data_11;
  reg                 io_in_c_bypass_regNext_11_0_is_stationary_11;
  reg        [15:0]   io_in_c_bypass_regNext_11_1_data_11;
  reg                 io_in_c_bypass_regNext_11_1_is_stationary_11;
  reg        [15:0]   io_in_c_bypass_regNext_11_2_data_11;
  reg                 io_in_c_bypass_regNext_11_2_is_stationary_11;
  reg        [15:0]   io_in_c_bypass_regNext_11_3_data_11;
  reg                 io_in_c_bypass_regNext_11_3_is_stationary_11;
  reg        [15:0]   io_in_c_bypass_regNext_12_0_data_11;
  reg                 io_in_c_bypass_regNext_12_0_is_stationary_11;
  reg        [15:0]   io_in_c_bypass_regNext_12_1_data_11;
  reg                 io_in_c_bypass_regNext_12_1_is_stationary_11;
  reg        [15:0]   io_in_c_bypass_regNext_12_2_data_11;
  reg                 io_in_c_bypass_regNext_12_2_is_stationary_11;
  reg        [15:0]   io_in_c_bypass_regNext_12_3_data_11;
  reg                 io_in_c_bypass_regNext_12_3_is_stationary_11;
  reg        [15:0]   io_in_c_bypass_regNext_13_0_data_11;
  reg                 io_in_c_bypass_regNext_13_0_is_stationary_11;
  reg        [15:0]   io_in_c_bypass_regNext_13_1_data_11;
  reg                 io_in_c_bypass_regNext_13_1_is_stationary_11;
  reg        [15:0]   io_in_c_bypass_regNext_13_2_data_11;
  reg                 io_in_c_bypass_regNext_13_2_is_stationary_11;
  reg        [15:0]   io_in_c_bypass_regNext_13_3_data_11;
  reg                 io_in_c_bypass_regNext_13_3_is_stationary_11;
  reg        [15:0]   io_in_c_bypass_regNext_14_0_data_11;
  reg                 io_in_c_bypass_regNext_14_0_is_stationary_11;
  reg        [15:0]   io_in_c_bypass_regNext_14_1_data_11;
  reg                 io_in_c_bypass_regNext_14_1_is_stationary_11;
  reg        [15:0]   io_in_c_bypass_regNext_14_2_data_11;
  reg                 io_in_c_bypass_regNext_14_2_is_stationary_11;
  reg        [15:0]   io_in_c_bypass_regNext_14_3_data_11;
  reg                 io_in_c_bypass_regNext_14_3_is_stationary_11;
  reg        [15:0]   io_in_c_bypass_regNext_15_0_data_11;
  reg                 io_in_c_bypass_regNext_15_0_is_stationary_11;
  reg        [15:0]   io_in_c_bypass_regNext_15_1_data_11;
  reg                 io_in_c_bypass_regNext_15_1_is_stationary_11;
  reg        [15:0]   io_in_c_bypass_regNext_15_2_data_11;
  reg                 io_in_c_bypass_regNext_15_2_is_stationary_11;
  reg        [15:0]   io_in_c_bypass_regNext_15_3_data_11;
  reg                 io_in_c_bypass_regNext_15_3_is_stationary_11;
  reg        [15:0]   io_in_c_bypass_regNext_16_0_data_11;
  reg                 io_in_c_bypass_regNext_16_0_is_stationary_11;
  reg        [15:0]   io_in_c_bypass_regNext_16_1_data_11;
  reg                 io_in_c_bypass_regNext_16_1_is_stationary_11;
  reg        [15:0]   io_in_c_bypass_regNext_16_2_data_11;
  reg                 io_in_c_bypass_regNext_16_2_is_stationary_11;
  reg        [15:0]   io_in_c_bypass_regNext_16_3_data_11;
  reg                 io_in_c_bypass_regNext_16_3_is_stationary_11;
  reg        [15:0]   io_in_c_bypass_regNext_17_0_data_11;
  reg                 io_in_c_bypass_regNext_17_0_is_stationary_11;
  reg        [15:0]   io_in_c_bypass_regNext_17_1_data_11;
  reg                 io_in_c_bypass_regNext_17_1_is_stationary_11;
  reg        [15:0]   io_in_c_bypass_regNext_17_2_data_11;
  reg                 io_in_c_bypass_regNext_17_2_is_stationary_11;
  reg        [15:0]   io_in_c_bypass_regNext_17_3_data_11;
  reg                 io_in_c_bypass_regNext_17_3_is_stationary_11;
  reg        [15:0]   io_in_c_bypass_regNext_18_0_data_11;
  reg                 io_in_c_bypass_regNext_18_0_is_stationary_11;
  reg        [15:0]   io_in_c_bypass_regNext_18_1_data_11;
  reg                 io_in_c_bypass_regNext_18_1_is_stationary_11;
  reg        [15:0]   io_in_c_bypass_regNext_18_2_data_11;
  reg                 io_in_c_bypass_regNext_18_2_is_stationary_11;
  reg        [15:0]   io_in_c_bypass_regNext_18_3_data_11;
  reg                 io_in_c_bypass_regNext_18_3_is_stationary_11;
  reg        [15:0]   io_in_c_bypass_regNext_19_0_data_11;
  reg                 io_in_c_bypass_regNext_19_0_is_stationary_11;
  reg        [15:0]   io_in_c_bypass_regNext_19_1_data_11;
  reg                 io_in_c_bypass_regNext_19_1_is_stationary_11;
  reg        [15:0]   io_in_c_bypass_regNext_19_2_data_11;
  reg                 io_in_c_bypass_regNext_19_2_is_stationary_11;
  reg        [15:0]   io_in_c_bypass_regNext_19_3_data_11;
  reg                 io_in_c_bypass_regNext_19_3_is_stationary_11;
  reg        [15:0]   io_in_c_bypass_regNext_20_0_data_11;
  reg                 io_in_c_bypass_regNext_20_0_is_stationary_11;
  reg        [15:0]   io_in_c_bypass_regNext_20_1_data_11;
  reg                 io_in_c_bypass_regNext_20_1_is_stationary_11;
  reg        [15:0]   io_in_c_bypass_regNext_20_2_data_11;
  reg                 io_in_c_bypass_regNext_20_2_is_stationary_11;
  reg        [15:0]   io_in_c_bypass_regNext_20_3_data_11;
  reg                 io_in_c_bypass_regNext_20_3_is_stationary_11;
  reg        [15:0]   io_in_c_bypass_regNext_21_0_data_11;
  reg                 io_in_c_bypass_regNext_21_0_is_stationary_11;
  reg        [15:0]   io_in_c_bypass_regNext_21_1_data_11;
  reg                 io_in_c_bypass_regNext_21_1_is_stationary_11;
  reg        [15:0]   io_in_c_bypass_regNext_21_2_data_11;
  reg                 io_in_c_bypass_regNext_21_2_is_stationary_11;
  reg        [15:0]   io_in_c_bypass_regNext_21_3_data_11;
  reg                 io_in_c_bypass_regNext_21_3_is_stationary_11;
  reg        [15:0]   io_in_c_bypass_regNext_22_0_data_11;
  reg                 io_in_c_bypass_regNext_22_0_is_stationary_11;
  reg        [15:0]   io_in_c_bypass_regNext_22_1_data_11;
  reg                 io_in_c_bypass_regNext_22_1_is_stationary_11;
  reg        [15:0]   io_in_c_bypass_regNext_22_2_data_11;
  reg                 io_in_c_bypass_regNext_22_2_is_stationary_11;
  reg        [15:0]   io_in_c_bypass_regNext_22_3_data_11;
  reg                 io_in_c_bypass_regNext_22_3_is_stationary_11;
  reg        [15:0]   io_in_c_bypass_regNext_23_0_data_11;
  reg                 io_in_c_bypass_regNext_23_0_is_stationary_11;
  reg        [15:0]   io_in_c_bypass_regNext_23_1_data_11;
  reg                 io_in_c_bypass_regNext_23_1_is_stationary_11;
  reg        [15:0]   io_in_c_bypass_regNext_23_2_data_11;
  reg                 io_in_c_bypass_regNext_23_2_is_stationary_11;
  reg        [15:0]   io_in_c_bypass_regNext_23_3_data_11;
  reg                 io_in_c_bypass_regNext_23_3_is_stationary_11;
  reg        [15:0]   io_in_c_bypass_regNext_24_0_data_11;
  reg                 io_in_c_bypass_regNext_24_0_is_stationary_11;
  reg        [15:0]   io_in_c_bypass_regNext_24_1_data_11;
  reg                 io_in_c_bypass_regNext_24_1_is_stationary_11;
  reg        [15:0]   io_in_c_bypass_regNext_24_2_data_11;
  reg                 io_in_c_bypass_regNext_24_2_is_stationary_11;
  reg        [15:0]   io_in_c_bypass_regNext_24_3_data_11;
  reg                 io_in_c_bypass_regNext_24_3_is_stationary_11;
  reg        [15:0]   io_in_c_bypass_regNext_25_0_data_11;
  reg                 io_in_c_bypass_regNext_25_0_is_stationary_11;
  reg        [15:0]   io_in_c_bypass_regNext_25_1_data_11;
  reg                 io_in_c_bypass_regNext_25_1_is_stationary_11;
  reg        [15:0]   io_in_c_bypass_regNext_25_2_data_11;
  reg                 io_in_c_bypass_regNext_25_2_is_stationary_11;
  reg        [15:0]   io_in_c_bypass_regNext_25_3_data_11;
  reg                 io_in_c_bypass_regNext_25_3_is_stationary_11;
  reg        [15:0]   io_in_c_bypass_regNext_26_0_data_11;
  reg                 io_in_c_bypass_regNext_26_0_is_stationary_11;
  reg        [15:0]   io_in_c_bypass_regNext_26_1_data_11;
  reg                 io_in_c_bypass_regNext_26_1_is_stationary_11;
  reg        [15:0]   io_in_c_bypass_regNext_26_2_data_11;
  reg                 io_in_c_bypass_regNext_26_2_is_stationary_11;
  reg        [15:0]   io_in_c_bypass_regNext_26_3_data_11;
  reg                 io_in_c_bypass_regNext_26_3_is_stationary_11;
  reg        [15:0]   io_in_c_bypass_regNext_27_0_data_11;
  reg                 io_in_c_bypass_regNext_27_0_is_stationary_11;
  reg        [15:0]   io_in_c_bypass_regNext_27_1_data_11;
  reg                 io_in_c_bypass_regNext_27_1_is_stationary_11;
  reg        [15:0]   io_in_c_bypass_regNext_27_2_data_11;
  reg                 io_in_c_bypass_regNext_27_2_is_stationary_11;
  reg        [15:0]   io_in_c_bypass_regNext_27_3_data_11;
  reg                 io_in_c_bypass_regNext_27_3_is_stationary_11;
  reg        [15:0]   io_in_c_bypass_regNext_28_0_data_11;
  reg                 io_in_c_bypass_regNext_28_0_is_stationary_11;
  reg        [15:0]   io_in_c_bypass_regNext_28_1_data_11;
  reg                 io_in_c_bypass_regNext_28_1_is_stationary_11;
  reg        [15:0]   io_in_c_bypass_regNext_28_2_data_11;
  reg                 io_in_c_bypass_regNext_28_2_is_stationary_11;
  reg        [15:0]   io_in_c_bypass_regNext_28_3_data_11;
  reg                 io_in_c_bypass_regNext_28_3_is_stationary_11;
  reg        [15:0]   io_in_c_bypass_regNext_29_0_data_11;
  reg                 io_in_c_bypass_regNext_29_0_is_stationary_11;
  reg        [15:0]   io_in_c_bypass_regNext_29_1_data_11;
  reg                 io_in_c_bypass_regNext_29_1_is_stationary_11;
  reg        [15:0]   io_in_c_bypass_regNext_29_2_data_11;
  reg                 io_in_c_bypass_regNext_29_2_is_stationary_11;
  reg        [15:0]   io_in_c_bypass_regNext_29_3_data_11;
  reg                 io_in_c_bypass_regNext_29_3_is_stationary_11;
  reg        [15:0]   io_in_c_bypass_regNext_30_0_data_11;
  reg                 io_in_c_bypass_regNext_30_0_is_stationary_11;
  reg        [15:0]   io_in_c_bypass_regNext_30_1_data_11;
  reg                 io_in_c_bypass_regNext_30_1_is_stationary_11;
  reg        [15:0]   io_in_c_bypass_regNext_30_2_data_11;
  reg                 io_in_c_bypass_regNext_30_2_is_stationary_11;
  reg        [15:0]   io_in_c_bypass_regNext_30_3_data_11;
  reg                 io_in_c_bypass_regNext_30_3_is_stationary_11;
  reg        [15:0]   io_in_c_bypass_regNext_31_0_data_11;
  reg                 io_in_c_bypass_regNext_31_0_is_stationary_11;
  reg        [15:0]   io_in_c_bypass_regNext_31_1_data_11;
  reg                 io_in_c_bypass_regNext_31_1_is_stationary_11;
  reg        [15:0]   io_in_c_bypass_regNext_31_2_data_11;
  reg                 io_in_c_bypass_regNext_31_2_is_stationary_11;
  reg        [15:0]   io_in_c_bypass_regNext_31_3_data_11;
  reg                 io_in_c_bypass_regNext_31_3_is_stationary_11;
  reg        [15:0]   io_in_c_bypass_regNext_0_0_data_12;
  reg                 io_in_c_bypass_regNext_0_0_is_stationary_12;
  reg        [15:0]   io_in_c_bypass_regNext_0_1_data_12;
  reg                 io_in_c_bypass_regNext_0_1_is_stationary_12;
  reg        [15:0]   io_in_c_bypass_regNext_0_2_data_12;
  reg                 io_in_c_bypass_regNext_0_2_is_stationary_12;
  reg        [15:0]   io_in_c_bypass_regNext_0_3_data_12;
  reg                 io_in_c_bypass_regNext_0_3_is_stationary_12;
  reg        [15:0]   io_in_c_bypass_regNext_1_0_data_12;
  reg                 io_in_c_bypass_regNext_1_0_is_stationary_12;
  reg        [15:0]   io_in_c_bypass_regNext_1_1_data_12;
  reg                 io_in_c_bypass_regNext_1_1_is_stationary_12;
  reg        [15:0]   io_in_c_bypass_regNext_1_2_data_12;
  reg                 io_in_c_bypass_regNext_1_2_is_stationary_12;
  reg        [15:0]   io_in_c_bypass_regNext_1_3_data_12;
  reg                 io_in_c_bypass_regNext_1_3_is_stationary_12;
  reg        [15:0]   io_in_c_bypass_regNext_2_0_data_12;
  reg                 io_in_c_bypass_regNext_2_0_is_stationary_12;
  reg        [15:0]   io_in_c_bypass_regNext_2_1_data_12;
  reg                 io_in_c_bypass_regNext_2_1_is_stationary_12;
  reg        [15:0]   io_in_c_bypass_regNext_2_2_data_12;
  reg                 io_in_c_bypass_regNext_2_2_is_stationary_12;
  reg        [15:0]   io_in_c_bypass_regNext_2_3_data_12;
  reg                 io_in_c_bypass_regNext_2_3_is_stationary_12;
  reg        [15:0]   io_in_c_bypass_regNext_3_0_data_12;
  reg                 io_in_c_bypass_regNext_3_0_is_stationary_12;
  reg        [15:0]   io_in_c_bypass_regNext_3_1_data_12;
  reg                 io_in_c_bypass_regNext_3_1_is_stationary_12;
  reg        [15:0]   io_in_c_bypass_regNext_3_2_data_12;
  reg                 io_in_c_bypass_regNext_3_2_is_stationary_12;
  reg        [15:0]   io_in_c_bypass_regNext_3_3_data_12;
  reg                 io_in_c_bypass_regNext_3_3_is_stationary_12;
  reg        [15:0]   io_in_c_bypass_regNext_4_0_data_12;
  reg                 io_in_c_bypass_regNext_4_0_is_stationary_12;
  reg        [15:0]   io_in_c_bypass_regNext_4_1_data_12;
  reg                 io_in_c_bypass_regNext_4_1_is_stationary_12;
  reg        [15:0]   io_in_c_bypass_regNext_4_2_data_12;
  reg                 io_in_c_bypass_regNext_4_2_is_stationary_12;
  reg        [15:0]   io_in_c_bypass_regNext_4_3_data_12;
  reg                 io_in_c_bypass_regNext_4_3_is_stationary_12;
  reg        [15:0]   io_in_c_bypass_regNext_5_0_data_12;
  reg                 io_in_c_bypass_regNext_5_0_is_stationary_12;
  reg        [15:0]   io_in_c_bypass_regNext_5_1_data_12;
  reg                 io_in_c_bypass_regNext_5_1_is_stationary_12;
  reg        [15:0]   io_in_c_bypass_regNext_5_2_data_12;
  reg                 io_in_c_bypass_regNext_5_2_is_stationary_12;
  reg        [15:0]   io_in_c_bypass_regNext_5_3_data_12;
  reg                 io_in_c_bypass_regNext_5_3_is_stationary_12;
  reg        [15:0]   io_in_c_bypass_regNext_6_0_data_12;
  reg                 io_in_c_bypass_regNext_6_0_is_stationary_12;
  reg        [15:0]   io_in_c_bypass_regNext_6_1_data_12;
  reg                 io_in_c_bypass_regNext_6_1_is_stationary_12;
  reg        [15:0]   io_in_c_bypass_regNext_6_2_data_12;
  reg                 io_in_c_bypass_regNext_6_2_is_stationary_12;
  reg        [15:0]   io_in_c_bypass_regNext_6_3_data_12;
  reg                 io_in_c_bypass_regNext_6_3_is_stationary_12;
  reg        [15:0]   io_in_c_bypass_regNext_7_0_data_12;
  reg                 io_in_c_bypass_regNext_7_0_is_stationary_12;
  reg        [15:0]   io_in_c_bypass_regNext_7_1_data_12;
  reg                 io_in_c_bypass_regNext_7_1_is_stationary_12;
  reg        [15:0]   io_in_c_bypass_regNext_7_2_data_12;
  reg                 io_in_c_bypass_regNext_7_2_is_stationary_12;
  reg        [15:0]   io_in_c_bypass_regNext_7_3_data_12;
  reg                 io_in_c_bypass_regNext_7_3_is_stationary_12;
  reg        [15:0]   io_in_c_bypass_regNext_8_0_data_12;
  reg                 io_in_c_bypass_regNext_8_0_is_stationary_12;
  reg        [15:0]   io_in_c_bypass_regNext_8_1_data_12;
  reg                 io_in_c_bypass_regNext_8_1_is_stationary_12;
  reg        [15:0]   io_in_c_bypass_regNext_8_2_data_12;
  reg                 io_in_c_bypass_regNext_8_2_is_stationary_12;
  reg        [15:0]   io_in_c_bypass_regNext_8_3_data_12;
  reg                 io_in_c_bypass_regNext_8_3_is_stationary_12;
  reg        [15:0]   io_in_c_bypass_regNext_9_0_data_12;
  reg                 io_in_c_bypass_regNext_9_0_is_stationary_12;
  reg        [15:0]   io_in_c_bypass_regNext_9_1_data_12;
  reg                 io_in_c_bypass_regNext_9_1_is_stationary_12;
  reg        [15:0]   io_in_c_bypass_regNext_9_2_data_12;
  reg                 io_in_c_bypass_regNext_9_2_is_stationary_12;
  reg        [15:0]   io_in_c_bypass_regNext_9_3_data_12;
  reg                 io_in_c_bypass_regNext_9_3_is_stationary_12;
  reg        [15:0]   io_in_c_bypass_regNext_10_0_data_12;
  reg                 io_in_c_bypass_regNext_10_0_is_stationary_12;
  reg        [15:0]   io_in_c_bypass_regNext_10_1_data_12;
  reg                 io_in_c_bypass_regNext_10_1_is_stationary_12;
  reg        [15:0]   io_in_c_bypass_regNext_10_2_data_12;
  reg                 io_in_c_bypass_regNext_10_2_is_stationary_12;
  reg        [15:0]   io_in_c_bypass_regNext_10_3_data_12;
  reg                 io_in_c_bypass_regNext_10_3_is_stationary_12;
  reg        [15:0]   io_in_c_bypass_regNext_11_0_data_12;
  reg                 io_in_c_bypass_regNext_11_0_is_stationary_12;
  reg        [15:0]   io_in_c_bypass_regNext_11_1_data_12;
  reg                 io_in_c_bypass_regNext_11_1_is_stationary_12;
  reg        [15:0]   io_in_c_bypass_regNext_11_2_data_12;
  reg                 io_in_c_bypass_regNext_11_2_is_stationary_12;
  reg        [15:0]   io_in_c_bypass_regNext_11_3_data_12;
  reg                 io_in_c_bypass_regNext_11_3_is_stationary_12;
  reg        [15:0]   io_in_c_bypass_regNext_12_0_data_12;
  reg                 io_in_c_bypass_regNext_12_0_is_stationary_12;
  reg        [15:0]   io_in_c_bypass_regNext_12_1_data_12;
  reg                 io_in_c_bypass_regNext_12_1_is_stationary_12;
  reg        [15:0]   io_in_c_bypass_regNext_12_2_data_12;
  reg                 io_in_c_bypass_regNext_12_2_is_stationary_12;
  reg        [15:0]   io_in_c_bypass_regNext_12_3_data_12;
  reg                 io_in_c_bypass_regNext_12_3_is_stationary_12;
  reg        [15:0]   io_in_c_bypass_regNext_13_0_data_12;
  reg                 io_in_c_bypass_regNext_13_0_is_stationary_12;
  reg        [15:0]   io_in_c_bypass_regNext_13_1_data_12;
  reg                 io_in_c_bypass_regNext_13_1_is_stationary_12;
  reg        [15:0]   io_in_c_bypass_regNext_13_2_data_12;
  reg                 io_in_c_bypass_regNext_13_2_is_stationary_12;
  reg        [15:0]   io_in_c_bypass_regNext_13_3_data_12;
  reg                 io_in_c_bypass_regNext_13_3_is_stationary_12;
  reg        [15:0]   io_in_c_bypass_regNext_14_0_data_12;
  reg                 io_in_c_bypass_regNext_14_0_is_stationary_12;
  reg        [15:0]   io_in_c_bypass_regNext_14_1_data_12;
  reg                 io_in_c_bypass_regNext_14_1_is_stationary_12;
  reg        [15:0]   io_in_c_bypass_regNext_14_2_data_12;
  reg                 io_in_c_bypass_regNext_14_2_is_stationary_12;
  reg        [15:0]   io_in_c_bypass_regNext_14_3_data_12;
  reg                 io_in_c_bypass_regNext_14_3_is_stationary_12;
  reg        [15:0]   io_in_c_bypass_regNext_15_0_data_12;
  reg                 io_in_c_bypass_regNext_15_0_is_stationary_12;
  reg        [15:0]   io_in_c_bypass_regNext_15_1_data_12;
  reg                 io_in_c_bypass_regNext_15_1_is_stationary_12;
  reg        [15:0]   io_in_c_bypass_regNext_15_2_data_12;
  reg                 io_in_c_bypass_regNext_15_2_is_stationary_12;
  reg        [15:0]   io_in_c_bypass_regNext_15_3_data_12;
  reg                 io_in_c_bypass_regNext_15_3_is_stationary_12;
  reg        [15:0]   io_in_c_bypass_regNext_16_0_data_12;
  reg                 io_in_c_bypass_regNext_16_0_is_stationary_12;
  reg        [15:0]   io_in_c_bypass_regNext_16_1_data_12;
  reg                 io_in_c_bypass_regNext_16_1_is_stationary_12;
  reg        [15:0]   io_in_c_bypass_regNext_16_2_data_12;
  reg                 io_in_c_bypass_regNext_16_2_is_stationary_12;
  reg        [15:0]   io_in_c_bypass_regNext_16_3_data_12;
  reg                 io_in_c_bypass_regNext_16_3_is_stationary_12;
  reg        [15:0]   io_in_c_bypass_regNext_17_0_data_12;
  reg                 io_in_c_bypass_regNext_17_0_is_stationary_12;
  reg        [15:0]   io_in_c_bypass_regNext_17_1_data_12;
  reg                 io_in_c_bypass_regNext_17_1_is_stationary_12;
  reg        [15:0]   io_in_c_bypass_regNext_17_2_data_12;
  reg                 io_in_c_bypass_regNext_17_2_is_stationary_12;
  reg        [15:0]   io_in_c_bypass_regNext_17_3_data_12;
  reg                 io_in_c_bypass_regNext_17_3_is_stationary_12;
  reg        [15:0]   io_in_c_bypass_regNext_18_0_data_12;
  reg                 io_in_c_bypass_regNext_18_0_is_stationary_12;
  reg        [15:0]   io_in_c_bypass_regNext_18_1_data_12;
  reg                 io_in_c_bypass_regNext_18_1_is_stationary_12;
  reg        [15:0]   io_in_c_bypass_regNext_18_2_data_12;
  reg                 io_in_c_bypass_regNext_18_2_is_stationary_12;
  reg        [15:0]   io_in_c_bypass_regNext_18_3_data_12;
  reg                 io_in_c_bypass_regNext_18_3_is_stationary_12;
  reg        [15:0]   io_in_c_bypass_regNext_19_0_data_12;
  reg                 io_in_c_bypass_regNext_19_0_is_stationary_12;
  reg        [15:0]   io_in_c_bypass_regNext_19_1_data_12;
  reg                 io_in_c_bypass_regNext_19_1_is_stationary_12;
  reg        [15:0]   io_in_c_bypass_regNext_19_2_data_12;
  reg                 io_in_c_bypass_regNext_19_2_is_stationary_12;
  reg        [15:0]   io_in_c_bypass_regNext_19_3_data_12;
  reg                 io_in_c_bypass_regNext_19_3_is_stationary_12;
  reg        [15:0]   io_in_c_bypass_regNext_20_0_data_12;
  reg                 io_in_c_bypass_regNext_20_0_is_stationary_12;
  reg        [15:0]   io_in_c_bypass_regNext_20_1_data_12;
  reg                 io_in_c_bypass_regNext_20_1_is_stationary_12;
  reg        [15:0]   io_in_c_bypass_regNext_20_2_data_12;
  reg                 io_in_c_bypass_regNext_20_2_is_stationary_12;
  reg        [15:0]   io_in_c_bypass_regNext_20_3_data_12;
  reg                 io_in_c_bypass_regNext_20_3_is_stationary_12;
  reg        [15:0]   io_in_c_bypass_regNext_21_0_data_12;
  reg                 io_in_c_bypass_regNext_21_0_is_stationary_12;
  reg        [15:0]   io_in_c_bypass_regNext_21_1_data_12;
  reg                 io_in_c_bypass_regNext_21_1_is_stationary_12;
  reg        [15:0]   io_in_c_bypass_regNext_21_2_data_12;
  reg                 io_in_c_bypass_regNext_21_2_is_stationary_12;
  reg        [15:0]   io_in_c_bypass_regNext_21_3_data_12;
  reg                 io_in_c_bypass_regNext_21_3_is_stationary_12;
  reg        [15:0]   io_in_c_bypass_regNext_22_0_data_12;
  reg                 io_in_c_bypass_regNext_22_0_is_stationary_12;
  reg        [15:0]   io_in_c_bypass_regNext_22_1_data_12;
  reg                 io_in_c_bypass_regNext_22_1_is_stationary_12;
  reg        [15:0]   io_in_c_bypass_regNext_22_2_data_12;
  reg                 io_in_c_bypass_regNext_22_2_is_stationary_12;
  reg        [15:0]   io_in_c_bypass_regNext_22_3_data_12;
  reg                 io_in_c_bypass_regNext_22_3_is_stationary_12;
  reg        [15:0]   io_in_c_bypass_regNext_23_0_data_12;
  reg                 io_in_c_bypass_regNext_23_0_is_stationary_12;
  reg        [15:0]   io_in_c_bypass_regNext_23_1_data_12;
  reg                 io_in_c_bypass_regNext_23_1_is_stationary_12;
  reg        [15:0]   io_in_c_bypass_regNext_23_2_data_12;
  reg                 io_in_c_bypass_regNext_23_2_is_stationary_12;
  reg        [15:0]   io_in_c_bypass_regNext_23_3_data_12;
  reg                 io_in_c_bypass_regNext_23_3_is_stationary_12;
  reg        [15:0]   io_in_c_bypass_regNext_24_0_data_12;
  reg                 io_in_c_bypass_regNext_24_0_is_stationary_12;
  reg        [15:0]   io_in_c_bypass_regNext_24_1_data_12;
  reg                 io_in_c_bypass_regNext_24_1_is_stationary_12;
  reg        [15:0]   io_in_c_bypass_regNext_24_2_data_12;
  reg                 io_in_c_bypass_regNext_24_2_is_stationary_12;
  reg        [15:0]   io_in_c_bypass_regNext_24_3_data_12;
  reg                 io_in_c_bypass_regNext_24_3_is_stationary_12;
  reg        [15:0]   io_in_c_bypass_regNext_25_0_data_12;
  reg                 io_in_c_bypass_regNext_25_0_is_stationary_12;
  reg        [15:0]   io_in_c_bypass_regNext_25_1_data_12;
  reg                 io_in_c_bypass_regNext_25_1_is_stationary_12;
  reg        [15:0]   io_in_c_bypass_regNext_25_2_data_12;
  reg                 io_in_c_bypass_regNext_25_2_is_stationary_12;
  reg        [15:0]   io_in_c_bypass_regNext_25_3_data_12;
  reg                 io_in_c_bypass_regNext_25_3_is_stationary_12;
  reg        [15:0]   io_in_c_bypass_regNext_26_0_data_12;
  reg                 io_in_c_bypass_regNext_26_0_is_stationary_12;
  reg        [15:0]   io_in_c_bypass_regNext_26_1_data_12;
  reg                 io_in_c_bypass_regNext_26_1_is_stationary_12;
  reg        [15:0]   io_in_c_bypass_regNext_26_2_data_12;
  reg                 io_in_c_bypass_regNext_26_2_is_stationary_12;
  reg        [15:0]   io_in_c_bypass_regNext_26_3_data_12;
  reg                 io_in_c_bypass_regNext_26_3_is_stationary_12;
  reg        [15:0]   io_in_c_bypass_regNext_27_0_data_12;
  reg                 io_in_c_bypass_regNext_27_0_is_stationary_12;
  reg        [15:0]   io_in_c_bypass_regNext_27_1_data_12;
  reg                 io_in_c_bypass_regNext_27_1_is_stationary_12;
  reg        [15:0]   io_in_c_bypass_regNext_27_2_data_12;
  reg                 io_in_c_bypass_regNext_27_2_is_stationary_12;
  reg        [15:0]   io_in_c_bypass_regNext_27_3_data_12;
  reg                 io_in_c_bypass_regNext_27_3_is_stationary_12;
  reg        [15:0]   io_in_c_bypass_regNext_28_0_data_12;
  reg                 io_in_c_bypass_regNext_28_0_is_stationary_12;
  reg        [15:0]   io_in_c_bypass_regNext_28_1_data_12;
  reg                 io_in_c_bypass_regNext_28_1_is_stationary_12;
  reg        [15:0]   io_in_c_bypass_regNext_28_2_data_12;
  reg                 io_in_c_bypass_regNext_28_2_is_stationary_12;
  reg        [15:0]   io_in_c_bypass_regNext_28_3_data_12;
  reg                 io_in_c_bypass_regNext_28_3_is_stationary_12;
  reg        [15:0]   io_in_c_bypass_regNext_29_0_data_12;
  reg                 io_in_c_bypass_regNext_29_0_is_stationary_12;
  reg        [15:0]   io_in_c_bypass_regNext_29_1_data_12;
  reg                 io_in_c_bypass_regNext_29_1_is_stationary_12;
  reg        [15:0]   io_in_c_bypass_regNext_29_2_data_12;
  reg                 io_in_c_bypass_regNext_29_2_is_stationary_12;
  reg        [15:0]   io_in_c_bypass_regNext_29_3_data_12;
  reg                 io_in_c_bypass_regNext_29_3_is_stationary_12;
  reg        [15:0]   io_in_c_bypass_regNext_30_0_data_12;
  reg                 io_in_c_bypass_regNext_30_0_is_stationary_12;
  reg        [15:0]   io_in_c_bypass_regNext_30_1_data_12;
  reg                 io_in_c_bypass_regNext_30_1_is_stationary_12;
  reg        [15:0]   io_in_c_bypass_regNext_30_2_data_12;
  reg                 io_in_c_bypass_regNext_30_2_is_stationary_12;
  reg        [15:0]   io_in_c_bypass_regNext_30_3_data_12;
  reg                 io_in_c_bypass_regNext_30_3_is_stationary_12;
  reg        [15:0]   io_in_c_bypass_regNext_31_0_data_12;
  reg                 io_in_c_bypass_regNext_31_0_is_stationary_12;
  reg        [15:0]   io_in_c_bypass_regNext_31_1_data_12;
  reg                 io_in_c_bypass_regNext_31_1_is_stationary_12;
  reg        [15:0]   io_in_c_bypass_regNext_31_2_data_12;
  reg                 io_in_c_bypass_regNext_31_2_is_stationary_12;
  reg        [15:0]   io_in_c_bypass_regNext_31_3_data_12;
  reg                 io_in_c_bypass_regNext_31_3_is_stationary_12;
  reg        [15:0]   io_in_c_bypass_regNext_0_0_data_13;
  reg                 io_in_c_bypass_regNext_0_0_is_stationary_13;
  reg        [15:0]   io_in_c_bypass_regNext_0_1_data_13;
  reg                 io_in_c_bypass_regNext_0_1_is_stationary_13;
  reg        [15:0]   io_in_c_bypass_regNext_0_2_data_13;
  reg                 io_in_c_bypass_regNext_0_2_is_stationary_13;
  reg        [15:0]   io_in_c_bypass_regNext_0_3_data_13;
  reg                 io_in_c_bypass_regNext_0_3_is_stationary_13;
  reg        [15:0]   io_in_c_bypass_regNext_1_0_data_13;
  reg                 io_in_c_bypass_regNext_1_0_is_stationary_13;
  reg        [15:0]   io_in_c_bypass_regNext_1_1_data_13;
  reg                 io_in_c_bypass_regNext_1_1_is_stationary_13;
  reg        [15:0]   io_in_c_bypass_regNext_1_2_data_13;
  reg                 io_in_c_bypass_regNext_1_2_is_stationary_13;
  reg        [15:0]   io_in_c_bypass_regNext_1_3_data_13;
  reg                 io_in_c_bypass_regNext_1_3_is_stationary_13;
  reg        [15:0]   io_in_c_bypass_regNext_2_0_data_13;
  reg                 io_in_c_bypass_regNext_2_0_is_stationary_13;
  reg        [15:0]   io_in_c_bypass_regNext_2_1_data_13;
  reg                 io_in_c_bypass_regNext_2_1_is_stationary_13;
  reg        [15:0]   io_in_c_bypass_regNext_2_2_data_13;
  reg                 io_in_c_bypass_regNext_2_2_is_stationary_13;
  reg        [15:0]   io_in_c_bypass_regNext_2_3_data_13;
  reg                 io_in_c_bypass_regNext_2_3_is_stationary_13;
  reg        [15:0]   io_in_c_bypass_regNext_3_0_data_13;
  reg                 io_in_c_bypass_regNext_3_0_is_stationary_13;
  reg        [15:0]   io_in_c_bypass_regNext_3_1_data_13;
  reg                 io_in_c_bypass_regNext_3_1_is_stationary_13;
  reg        [15:0]   io_in_c_bypass_regNext_3_2_data_13;
  reg                 io_in_c_bypass_regNext_3_2_is_stationary_13;
  reg        [15:0]   io_in_c_bypass_regNext_3_3_data_13;
  reg                 io_in_c_bypass_regNext_3_3_is_stationary_13;
  reg        [15:0]   io_in_c_bypass_regNext_4_0_data_13;
  reg                 io_in_c_bypass_regNext_4_0_is_stationary_13;
  reg        [15:0]   io_in_c_bypass_regNext_4_1_data_13;
  reg                 io_in_c_bypass_regNext_4_1_is_stationary_13;
  reg        [15:0]   io_in_c_bypass_regNext_4_2_data_13;
  reg                 io_in_c_bypass_regNext_4_2_is_stationary_13;
  reg        [15:0]   io_in_c_bypass_regNext_4_3_data_13;
  reg                 io_in_c_bypass_regNext_4_3_is_stationary_13;
  reg        [15:0]   io_in_c_bypass_regNext_5_0_data_13;
  reg                 io_in_c_bypass_regNext_5_0_is_stationary_13;
  reg        [15:0]   io_in_c_bypass_regNext_5_1_data_13;
  reg                 io_in_c_bypass_regNext_5_1_is_stationary_13;
  reg        [15:0]   io_in_c_bypass_regNext_5_2_data_13;
  reg                 io_in_c_bypass_regNext_5_2_is_stationary_13;
  reg        [15:0]   io_in_c_bypass_regNext_5_3_data_13;
  reg                 io_in_c_bypass_regNext_5_3_is_stationary_13;
  reg        [15:0]   io_in_c_bypass_regNext_6_0_data_13;
  reg                 io_in_c_bypass_regNext_6_0_is_stationary_13;
  reg        [15:0]   io_in_c_bypass_regNext_6_1_data_13;
  reg                 io_in_c_bypass_regNext_6_1_is_stationary_13;
  reg        [15:0]   io_in_c_bypass_regNext_6_2_data_13;
  reg                 io_in_c_bypass_regNext_6_2_is_stationary_13;
  reg        [15:0]   io_in_c_bypass_regNext_6_3_data_13;
  reg                 io_in_c_bypass_regNext_6_3_is_stationary_13;
  reg        [15:0]   io_in_c_bypass_regNext_7_0_data_13;
  reg                 io_in_c_bypass_regNext_7_0_is_stationary_13;
  reg        [15:0]   io_in_c_bypass_regNext_7_1_data_13;
  reg                 io_in_c_bypass_regNext_7_1_is_stationary_13;
  reg        [15:0]   io_in_c_bypass_regNext_7_2_data_13;
  reg                 io_in_c_bypass_regNext_7_2_is_stationary_13;
  reg        [15:0]   io_in_c_bypass_regNext_7_3_data_13;
  reg                 io_in_c_bypass_regNext_7_3_is_stationary_13;
  reg        [15:0]   io_in_c_bypass_regNext_8_0_data_13;
  reg                 io_in_c_bypass_regNext_8_0_is_stationary_13;
  reg        [15:0]   io_in_c_bypass_regNext_8_1_data_13;
  reg                 io_in_c_bypass_regNext_8_1_is_stationary_13;
  reg        [15:0]   io_in_c_bypass_regNext_8_2_data_13;
  reg                 io_in_c_bypass_regNext_8_2_is_stationary_13;
  reg        [15:0]   io_in_c_bypass_regNext_8_3_data_13;
  reg                 io_in_c_bypass_regNext_8_3_is_stationary_13;
  reg        [15:0]   io_in_c_bypass_regNext_9_0_data_13;
  reg                 io_in_c_bypass_regNext_9_0_is_stationary_13;
  reg        [15:0]   io_in_c_bypass_regNext_9_1_data_13;
  reg                 io_in_c_bypass_regNext_9_1_is_stationary_13;
  reg        [15:0]   io_in_c_bypass_regNext_9_2_data_13;
  reg                 io_in_c_bypass_regNext_9_2_is_stationary_13;
  reg        [15:0]   io_in_c_bypass_regNext_9_3_data_13;
  reg                 io_in_c_bypass_regNext_9_3_is_stationary_13;
  reg        [15:0]   io_in_c_bypass_regNext_10_0_data_13;
  reg                 io_in_c_bypass_regNext_10_0_is_stationary_13;
  reg        [15:0]   io_in_c_bypass_regNext_10_1_data_13;
  reg                 io_in_c_bypass_regNext_10_1_is_stationary_13;
  reg        [15:0]   io_in_c_bypass_regNext_10_2_data_13;
  reg                 io_in_c_bypass_regNext_10_2_is_stationary_13;
  reg        [15:0]   io_in_c_bypass_regNext_10_3_data_13;
  reg                 io_in_c_bypass_regNext_10_3_is_stationary_13;
  reg        [15:0]   io_in_c_bypass_regNext_11_0_data_13;
  reg                 io_in_c_bypass_regNext_11_0_is_stationary_13;
  reg        [15:0]   io_in_c_bypass_regNext_11_1_data_13;
  reg                 io_in_c_bypass_regNext_11_1_is_stationary_13;
  reg        [15:0]   io_in_c_bypass_regNext_11_2_data_13;
  reg                 io_in_c_bypass_regNext_11_2_is_stationary_13;
  reg        [15:0]   io_in_c_bypass_regNext_11_3_data_13;
  reg                 io_in_c_bypass_regNext_11_3_is_stationary_13;
  reg        [15:0]   io_in_c_bypass_regNext_12_0_data_13;
  reg                 io_in_c_bypass_regNext_12_0_is_stationary_13;
  reg        [15:0]   io_in_c_bypass_regNext_12_1_data_13;
  reg                 io_in_c_bypass_regNext_12_1_is_stationary_13;
  reg        [15:0]   io_in_c_bypass_regNext_12_2_data_13;
  reg                 io_in_c_bypass_regNext_12_2_is_stationary_13;
  reg        [15:0]   io_in_c_bypass_regNext_12_3_data_13;
  reg                 io_in_c_bypass_regNext_12_3_is_stationary_13;
  reg        [15:0]   io_in_c_bypass_regNext_13_0_data_13;
  reg                 io_in_c_bypass_regNext_13_0_is_stationary_13;
  reg        [15:0]   io_in_c_bypass_regNext_13_1_data_13;
  reg                 io_in_c_bypass_regNext_13_1_is_stationary_13;
  reg        [15:0]   io_in_c_bypass_regNext_13_2_data_13;
  reg                 io_in_c_bypass_regNext_13_2_is_stationary_13;
  reg        [15:0]   io_in_c_bypass_regNext_13_3_data_13;
  reg                 io_in_c_bypass_regNext_13_3_is_stationary_13;
  reg        [15:0]   io_in_c_bypass_regNext_14_0_data_13;
  reg                 io_in_c_bypass_regNext_14_0_is_stationary_13;
  reg        [15:0]   io_in_c_bypass_regNext_14_1_data_13;
  reg                 io_in_c_bypass_regNext_14_1_is_stationary_13;
  reg        [15:0]   io_in_c_bypass_regNext_14_2_data_13;
  reg                 io_in_c_bypass_regNext_14_2_is_stationary_13;
  reg        [15:0]   io_in_c_bypass_regNext_14_3_data_13;
  reg                 io_in_c_bypass_regNext_14_3_is_stationary_13;
  reg        [15:0]   io_in_c_bypass_regNext_15_0_data_13;
  reg                 io_in_c_bypass_regNext_15_0_is_stationary_13;
  reg        [15:0]   io_in_c_bypass_regNext_15_1_data_13;
  reg                 io_in_c_bypass_regNext_15_1_is_stationary_13;
  reg        [15:0]   io_in_c_bypass_regNext_15_2_data_13;
  reg                 io_in_c_bypass_regNext_15_2_is_stationary_13;
  reg        [15:0]   io_in_c_bypass_regNext_15_3_data_13;
  reg                 io_in_c_bypass_regNext_15_3_is_stationary_13;
  reg        [15:0]   io_in_c_bypass_regNext_16_0_data_13;
  reg                 io_in_c_bypass_regNext_16_0_is_stationary_13;
  reg        [15:0]   io_in_c_bypass_regNext_16_1_data_13;
  reg                 io_in_c_bypass_regNext_16_1_is_stationary_13;
  reg        [15:0]   io_in_c_bypass_regNext_16_2_data_13;
  reg                 io_in_c_bypass_regNext_16_2_is_stationary_13;
  reg        [15:0]   io_in_c_bypass_regNext_16_3_data_13;
  reg                 io_in_c_bypass_regNext_16_3_is_stationary_13;
  reg        [15:0]   io_in_c_bypass_regNext_17_0_data_13;
  reg                 io_in_c_bypass_regNext_17_0_is_stationary_13;
  reg        [15:0]   io_in_c_bypass_regNext_17_1_data_13;
  reg                 io_in_c_bypass_regNext_17_1_is_stationary_13;
  reg        [15:0]   io_in_c_bypass_regNext_17_2_data_13;
  reg                 io_in_c_bypass_regNext_17_2_is_stationary_13;
  reg        [15:0]   io_in_c_bypass_regNext_17_3_data_13;
  reg                 io_in_c_bypass_regNext_17_3_is_stationary_13;
  reg        [15:0]   io_in_c_bypass_regNext_18_0_data_13;
  reg                 io_in_c_bypass_regNext_18_0_is_stationary_13;
  reg        [15:0]   io_in_c_bypass_regNext_18_1_data_13;
  reg                 io_in_c_bypass_regNext_18_1_is_stationary_13;
  reg        [15:0]   io_in_c_bypass_regNext_18_2_data_13;
  reg                 io_in_c_bypass_regNext_18_2_is_stationary_13;
  reg        [15:0]   io_in_c_bypass_regNext_18_3_data_13;
  reg                 io_in_c_bypass_regNext_18_3_is_stationary_13;
  reg        [15:0]   io_in_c_bypass_regNext_19_0_data_13;
  reg                 io_in_c_bypass_regNext_19_0_is_stationary_13;
  reg        [15:0]   io_in_c_bypass_regNext_19_1_data_13;
  reg                 io_in_c_bypass_regNext_19_1_is_stationary_13;
  reg        [15:0]   io_in_c_bypass_regNext_19_2_data_13;
  reg                 io_in_c_bypass_regNext_19_2_is_stationary_13;
  reg        [15:0]   io_in_c_bypass_regNext_19_3_data_13;
  reg                 io_in_c_bypass_regNext_19_3_is_stationary_13;
  reg        [15:0]   io_in_c_bypass_regNext_20_0_data_13;
  reg                 io_in_c_bypass_regNext_20_0_is_stationary_13;
  reg        [15:0]   io_in_c_bypass_regNext_20_1_data_13;
  reg                 io_in_c_bypass_regNext_20_1_is_stationary_13;
  reg        [15:0]   io_in_c_bypass_regNext_20_2_data_13;
  reg                 io_in_c_bypass_regNext_20_2_is_stationary_13;
  reg        [15:0]   io_in_c_bypass_regNext_20_3_data_13;
  reg                 io_in_c_bypass_regNext_20_3_is_stationary_13;
  reg        [15:0]   io_in_c_bypass_regNext_21_0_data_13;
  reg                 io_in_c_bypass_regNext_21_0_is_stationary_13;
  reg        [15:0]   io_in_c_bypass_regNext_21_1_data_13;
  reg                 io_in_c_bypass_regNext_21_1_is_stationary_13;
  reg        [15:0]   io_in_c_bypass_regNext_21_2_data_13;
  reg                 io_in_c_bypass_regNext_21_2_is_stationary_13;
  reg        [15:0]   io_in_c_bypass_regNext_21_3_data_13;
  reg                 io_in_c_bypass_regNext_21_3_is_stationary_13;
  reg        [15:0]   io_in_c_bypass_regNext_22_0_data_13;
  reg                 io_in_c_bypass_regNext_22_0_is_stationary_13;
  reg        [15:0]   io_in_c_bypass_regNext_22_1_data_13;
  reg                 io_in_c_bypass_regNext_22_1_is_stationary_13;
  reg        [15:0]   io_in_c_bypass_regNext_22_2_data_13;
  reg                 io_in_c_bypass_regNext_22_2_is_stationary_13;
  reg        [15:0]   io_in_c_bypass_regNext_22_3_data_13;
  reg                 io_in_c_bypass_regNext_22_3_is_stationary_13;
  reg        [15:0]   io_in_c_bypass_regNext_23_0_data_13;
  reg                 io_in_c_bypass_regNext_23_0_is_stationary_13;
  reg        [15:0]   io_in_c_bypass_regNext_23_1_data_13;
  reg                 io_in_c_bypass_regNext_23_1_is_stationary_13;
  reg        [15:0]   io_in_c_bypass_regNext_23_2_data_13;
  reg                 io_in_c_bypass_regNext_23_2_is_stationary_13;
  reg        [15:0]   io_in_c_bypass_regNext_23_3_data_13;
  reg                 io_in_c_bypass_regNext_23_3_is_stationary_13;
  reg        [15:0]   io_in_c_bypass_regNext_24_0_data_13;
  reg                 io_in_c_bypass_regNext_24_0_is_stationary_13;
  reg        [15:0]   io_in_c_bypass_regNext_24_1_data_13;
  reg                 io_in_c_bypass_regNext_24_1_is_stationary_13;
  reg        [15:0]   io_in_c_bypass_regNext_24_2_data_13;
  reg                 io_in_c_bypass_regNext_24_2_is_stationary_13;
  reg        [15:0]   io_in_c_bypass_regNext_24_3_data_13;
  reg                 io_in_c_bypass_regNext_24_3_is_stationary_13;
  reg        [15:0]   io_in_c_bypass_regNext_25_0_data_13;
  reg                 io_in_c_bypass_regNext_25_0_is_stationary_13;
  reg        [15:0]   io_in_c_bypass_regNext_25_1_data_13;
  reg                 io_in_c_bypass_regNext_25_1_is_stationary_13;
  reg        [15:0]   io_in_c_bypass_regNext_25_2_data_13;
  reg                 io_in_c_bypass_regNext_25_2_is_stationary_13;
  reg        [15:0]   io_in_c_bypass_regNext_25_3_data_13;
  reg                 io_in_c_bypass_regNext_25_3_is_stationary_13;
  reg        [15:0]   io_in_c_bypass_regNext_26_0_data_13;
  reg                 io_in_c_bypass_regNext_26_0_is_stationary_13;
  reg        [15:0]   io_in_c_bypass_regNext_26_1_data_13;
  reg                 io_in_c_bypass_regNext_26_1_is_stationary_13;
  reg        [15:0]   io_in_c_bypass_regNext_26_2_data_13;
  reg                 io_in_c_bypass_regNext_26_2_is_stationary_13;
  reg        [15:0]   io_in_c_bypass_regNext_26_3_data_13;
  reg                 io_in_c_bypass_regNext_26_3_is_stationary_13;
  reg        [15:0]   io_in_c_bypass_regNext_27_0_data_13;
  reg                 io_in_c_bypass_regNext_27_0_is_stationary_13;
  reg        [15:0]   io_in_c_bypass_regNext_27_1_data_13;
  reg                 io_in_c_bypass_regNext_27_1_is_stationary_13;
  reg        [15:0]   io_in_c_bypass_regNext_27_2_data_13;
  reg                 io_in_c_bypass_regNext_27_2_is_stationary_13;
  reg        [15:0]   io_in_c_bypass_regNext_27_3_data_13;
  reg                 io_in_c_bypass_regNext_27_3_is_stationary_13;
  reg        [15:0]   io_in_c_bypass_regNext_28_0_data_13;
  reg                 io_in_c_bypass_regNext_28_0_is_stationary_13;
  reg        [15:0]   io_in_c_bypass_regNext_28_1_data_13;
  reg                 io_in_c_bypass_regNext_28_1_is_stationary_13;
  reg        [15:0]   io_in_c_bypass_regNext_28_2_data_13;
  reg                 io_in_c_bypass_regNext_28_2_is_stationary_13;
  reg        [15:0]   io_in_c_bypass_regNext_28_3_data_13;
  reg                 io_in_c_bypass_regNext_28_3_is_stationary_13;
  reg        [15:0]   io_in_c_bypass_regNext_29_0_data_13;
  reg                 io_in_c_bypass_regNext_29_0_is_stationary_13;
  reg        [15:0]   io_in_c_bypass_regNext_29_1_data_13;
  reg                 io_in_c_bypass_regNext_29_1_is_stationary_13;
  reg        [15:0]   io_in_c_bypass_regNext_29_2_data_13;
  reg                 io_in_c_bypass_regNext_29_2_is_stationary_13;
  reg        [15:0]   io_in_c_bypass_regNext_29_3_data_13;
  reg                 io_in_c_bypass_regNext_29_3_is_stationary_13;
  reg        [15:0]   io_in_c_bypass_regNext_30_0_data_13;
  reg                 io_in_c_bypass_regNext_30_0_is_stationary_13;
  reg        [15:0]   io_in_c_bypass_regNext_30_1_data_13;
  reg                 io_in_c_bypass_regNext_30_1_is_stationary_13;
  reg        [15:0]   io_in_c_bypass_regNext_30_2_data_13;
  reg                 io_in_c_bypass_regNext_30_2_is_stationary_13;
  reg        [15:0]   io_in_c_bypass_regNext_30_3_data_13;
  reg                 io_in_c_bypass_regNext_30_3_is_stationary_13;
  reg        [15:0]   io_in_c_bypass_regNext_31_0_data_13;
  reg                 io_in_c_bypass_regNext_31_0_is_stationary_13;
  reg        [15:0]   io_in_c_bypass_regNext_31_1_data_13;
  reg                 io_in_c_bypass_regNext_31_1_is_stationary_13;
  reg        [15:0]   io_in_c_bypass_regNext_31_2_data_13;
  reg                 io_in_c_bypass_regNext_31_2_is_stationary_13;
  reg        [15:0]   io_in_c_bypass_regNext_31_3_data_13;
  reg                 io_in_c_bypass_regNext_31_3_is_stationary_13;
  reg        [15:0]   io_in_c_bypass_regNext_0_0_data_14;
  reg                 io_in_c_bypass_regNext_0_0_is_stationary_14;
  reg        [15:0]   io_in_c_bypass_regNext_0_1_data_14;
  reg                 io_in_c_bypass_regNext_0_1_is_stationary_14;
  reg        [15:0]   io_in_c_bypass_regNext_0_2_data_14;
  reg                 io_in_c_bypass_regNext_0_2_is_stationary_14;
  reg        [15:0]   io_in_c_bypass_regNext_0_3_data_14;
  reg                 io_in_c_bypass_regNext_0_3_is_stationary_14;
  reg        [15:0]   io_in_c_bypass_regNext_1_0_data_14;
  reg                 io_in_c_bypass_regNext_1_0_is_stationary_14;
  reg        [15:0]   io_in_c_bypass_regNext_1_1_data_14;
  reg                 io_in_c_bypass_regNext_1_1_is_stationary_14;
  reg        [15:0]   io_in_c_bypass_regNext_1_2_data_14;
  reg                 io_in_c_bypass_regNext_1_2_is_stationary_14;
  reg        [15:0]   io_in_c_bypass_regNext_1_3_data_14;
  reg                 io_in_c_bypass_regNext_1_3_is_stationary_14;
  reg        [15:0]   io_in_c_bypass_regNext_2_0_data_14;
  reg                 io_in_c_bypass_regNext_2_0_is_stationary_14;
  reg        [15:0]   io_in_c_bypass_regNext_2_1_data_14;
  reg                 io_in_c_bypass_regNext_2_1_is_stationary_14;
  reg        [15:0]   io_in_c_bypass_regNext_2_2_data_14;
  reg                 io_in_c_bypass_regNext_2_2_is_stationary_14;
  reg        [15:0]   io_in_c_bypass_regNext_2_3_data_14;
  reg                 io_in_c_bypass_regNext_2_3_is_stationary_14;
  reg        [15:0]   io_in_c_bypass_regNext_3_0_data_14;
  reg                 io_in_c_bypass_regNext_3_0_is_stationary_14;
  reg        [15:0]   io_in_c_bypass_regNext_3_1_data_14;
  reg                 io_in_c_bypass_regNext_3_1_is_stationary_14;
  reg        [15:0]   io_in_c_bypass_regNext_3_2_data_14;
  reg                 io_in_c_bypass_regNext_3_2_is_stationary_14;
  reg        [15:0]   io_in_c_bypass_regNext_3_3_data_14;
  reg                 io_in_c_bypass_regNext_3_3_is_stationary_14;
  reg        [15:0]   io_in_c_bypass_regNext_4_0_data_14;
  reg                 io_in_c_bypass_regNext_4_0_is_stationary_14;
  reg        [15:0]   io_in_c_bypass_regNext_4_1_data_14;
  reg                 io_in_c_bypass_regNext_4_1_is_stationary_14;
  reg        [15:0]   io_in_c_bypass_regNext_4_2_data_14;
  reg                 io_in_c_bypass_regNext_4_2_is_stationary_14;
  reg        [15:0]   io_in_c_bypass_regNext_4_3_data_14;
  reg                 io_in_c_bypass_regNext_4_3_is_stationary_14;
  reg        [15:0]   io_in_c_bypass_regNext_5_0_data_14;
  reg                 io_in_c_bypass_regNext_5_0_is_stationary_14;
  reg        [15:0]   io_in_c_bypass_regNext_5_1_data_14;
  reg                 io_in_c_bypass_regNext_5_1_is_stationary_14;
  reg        [15:0]   io_in_c_bypass_regNext_5_2_data_14;
  reg                 io_in_c_bypass_regNext_5_2_is_stationary_14;
  reg        [15:0]   io_in_c_bypass_regNext_5_3_data_14;
  reg                 io_in_c_bypass_regNext_5_3_is_stationary_14;
  reg        [15:0]   io_in_c_bypass_regNext_6_0_data_14;
  reg                 io_in_c_bypass_regNext_6_0_is_stationary_14;
  reg        [15:0]   io_in_c_bypass_regNext_6_1_data_14;
  reg                 io_in_c_bypass_regNext_6_1_is_stationary_14;
  reg        [15:0]   io_in_c_bypass_regNext_6_2_data_14;
  reg                 io_in_c_bypass_regNext_6_2_is_stationary_14;
  reg        [15:0]   io_in_c_bypass_regNext_6_3_data_14;
  reg                 io_in_c_bypass_regNext_6_3_is_stationary_14;
  reg        [15:0]   io_in_c_bypass_regNext_7_0_data_14;
  reg                 io_in_c_bypass_regNext_7_0_is_stationary_14;
  reg        [15:0]   io_in_c_bypass_regNext_7_1_data_14;
  reg                 io_in_c_bypass_regNext_7_1_is_stationary_14;
  reg        [15:0]   io_in_c_bypass_regNext_7_2_data_14;
  reg                 io_in_c_bypass_regNext_7_2_is_stationary_14;
  reg        [15:0]   io_in_c_bypass_regNext_7_3_data_14;
  reg                 io_in_c_bypass_regNext_7_3_is_stationary_14;
  reg        [15:0]   io_in_c_bypass_regNext_8_0_data_14;
  reg                 io_in_c_bypass_regNext_8_0_is_stationary_14;
  reg        [15:0]   io_in_c_bypass_regNext_8_1_data_14;
  reg                 io_in_c_bypass_regNext_8_1_is_stationary_14;
  reg        [15:0]   io_in_c_bypass_regNext_8_2_data_14;
  reg                 io_in_c_bypass_regNext_8_2_is_stationary_14;
  reg        [15:0]   io_in_c_bypass_regNext_8_3_data_14;
  reg                 io_in_c_bypass_regNext_8_3_is_stationary_14;
  reg        [15:0]   io_in_c_bypass_regNext_9_0_data_14;
  reg                 io_in_c_bypass_regNext_9_0_is_stationary_14;
  reg        [15:0]   io_in_c_bypass_regNext_9_1_data_14;
  reg                 io_in_c_bypass_regNext_9_1_is_stationary_14;
  reg        [15:0]   io_in_c_bypass_regNext_9_2_data_14;
  reg                 io_in_c_bypass_regNext_9_2_is_stationary_14;
  reg        [15:0]   io_in_c_bypass_regNext_9_3_data_14;
  reg                 io_in_c_bypass_regNext_9_3_is_stationary_14;
  reg        [15:0]   io_in_c_bypass_regNext_10_0_data_14;
  reg                 io_in_c_bypass_regNext_10_0_is_stationary_14;
  reg        [15:0]   io_in_c_bypass_regNext_10_1_data_14;
  reg                 io_in_c_bypass_regNext_10_1_is_stationary_14;
  reg        [15:0]   io_in_c_bypass_regNext_10_2_data_14;
  reg                 io_in_c_bypass_regNext_10_2_is_stationary_14;
  reg        [15:0]   io_in_c_bypass_regNext_10_3_data_14;
  reg                 io_in_c_bypass_regNext_10_3_is_stationary_14;
  reg        [15:0]   io_in_c_bypass_regNext_11_0_data_14;
  reg                 io_in_c_bypass_regNext_11_0_is_stationary_14;
  reg        [15:0]   io_in_c_bypass_regNext_11_1_data_14;
  reg                 io_in_c_bypass_regNext_11_1_is_stationary_14;
  reg        [15:0]   io_in_c_bypass_regNext_11_2_data_14;
  reg                 io_in_c_bypass_regNext_11_2_is_stationary_14;
  reg        [15:0]   io_in_c_bypass_regNext_11_3_data_14;
  reg                 io_in_c_bypass_regNext_11_3_is_stationary_14;
  reg        [15:0]   io_in_c_bypass_regNext_12_0_data_14;
  reg                 io_in_c_bypass_regNext_12_0_is_stationary_14;
  reg        [15:0]   io_in_c_bypass_regNext_12_1_data_14;
  reg                 io_in_c_bypass_regNext_12_1_is_stationary_14;
  reg        [15:0]   io_in_c_bypass_regNext_12_2_data_14;
  reg                 io_in_c_bypass_regNext_12_2_is_stationary_14;
  reg        [15:0]   io_in_c_bypass_regNext_12_3_data_14;
  reg                 io_in_c_bypass_regNext_12_3_is_stationary_14;
  reg        [15:0]   io_in_c_bypass_regNext_13_0_data_14;
  reg                 io_in_c_bypass_regNext_13_0_is_stationary_14;
  reg        [15:0]   io_in_c_bypass_regNext_13_1_data_14;
  reg                 io_in_c_bypass_regNext_13_1_is_stationary_14;
  reg        [15:0]   io_in_c_bypass_regNext_13_2_data_14;
  reg                 io_in_c_bypass_regNext_13_2_is_stationary_14;
  reg        [15:0]   io_in_c_bypass_regNext_13_3_data_14;
  reg                 io_in_c_bypass_regNext_13_3_is_stationary_14;
  reg        [15:0]   io_in_c_bypass_regNext_14_0_data_14;
  reg                 io_in_c_bypass_regNext_14_0_is_stationary_14;
  reg        [15:0]   io_in_c_bypass_regNext_14_1_data_14;
  reg                 io_in_c_bypass_regNext_14_1_is_stationary_14;
  reg        [15:0]   io_in_c_bypass_regNext_14_2_data_14;
  reg                 io_in_c_bypass_regNext_14_2_is_stationary_14;
  reg        [15:0]   io_in_c_bypass_regNext_14_3_data_14;
  reg                 io_in_c_bypass_regNext_14_3_is_stationary_14;
  reg        [15:0]   io_in_c_bypass_regNext_15_0_data_14;
  reg                 io_in_c_bypass_regNext_15_0_is_stationary_14;
  reg        [15:0]   io_in_c_bypass_regNext_15_1_data_14;
  reg                 io_in_c_bypass_regNext_15_1_is_stationary_14;
  reg        [15:0]   io_in_c_bypass_regNext_15_2_data_14;
  reg                 io_in_c_bypass_regNext_15_2_is_stationary_14;
  reg        [15:0]   io_in_c_bypass_regNext_15_3_data_14;
  reg                 io_in_c_bypass_regNext_15_3_is_stationary_14;
  reg        [15:0]   io_in_c_bypass_regNext_16_0_data_14;
  reg                 io_in_c_bypass_regNext_16_0_is_stationary_14;
  reg        [15:0]   io_in_c_bypass_regNext_16_1_data_14;
  reg                 io_in_c_bypass_regNext_16_1_is_stationary_14;
  reg        [15:0]   io_in_c_bypass_regNext_16_2_data_14;
  reg                 io_in_c_bypass_regNext_16_2_is_stationary_14;
  reg        [15:0]   io_in_c_bypass_regNext_16_3_data_14;
  reg                 io_in_c_bypass_regNext_16_3_is_stationary_14;
  reg        [15:0]   io_in_c_bypass_regNext_17_0_data_14;
  reg                 io_in_c_bypass_regNext_17_0_is_stationary_14;
  reg        [15:0]   io_in_c_bypass_regNext_17_1_data_14;
  reg                 io_in_c_bypass_regNext_17_1_is_stationary_14;
  reg        [15:0]   io_in_c_bypass_regNext_17_2_data_14;
  reg                 io_in_c_bypass_regNext_17_2_is_stationary_14;
  reg        [15:0]   io_in_c_bypass_regNext_17_3_data_14;
  reg                 io_in_c_bypass_regNext_17_3_is_stationary_14;
  reg        [15:0]   io_in_c_bypass_regNext_18_0_data_14;
  reg                 io_in_c_bypass_regNext_18_0_is_stationary_14;
  reg        [15:0]   io_in_c_bypass_regNext_18_1_data_14;
  reg                 io_in_c_bypass_regNext_18_1_is_stationary_14;
  reg        [15:0]   io_in_c_bypass_regNext_18_2_data_14;
  reg                 io_in_c_bypass_regNext_18_2_is_stationary_14;
  reg        [15:0]   io_in_c_bypass_regNext_18_3_data_14;
  reg                 io_in_c_bypass_regNext_18_3_is_stationary_14;
  reg        [15:0]   io_in_c_bypass_regNext_19_0_data_14;
  reg                 io_in_c_bypass_regNext_19_0_is_stationary_14;
  reg        [15:0]   io_in_c_bypass_regNext_19_1_data_14;
  reg                 io_in_c_bypass_regNext_19_1_is_stationary_14;
  reg        [15:0]   io_in_c_bypass_regNext_19_2_data_14;
  reg                 io_in_c_bypass_regNext_19_2_is_stationary_14;
  reg        [15:0]   io_in_c_bypass_regNext_19_3_data_14;
  reg                 io_in_c_bypass_regNext_19_3_is_stationary_14;
  reg        [15:0]   io_in_c_bypass_regNext_20_0_data_14;
  reg                 io_in_c_bypass_regNext_20_0_is_stationary_14;
  reg        [15:0]   io_in_c_bypass_regNext_20_1_data_14;
  reg                 io_in_c_bypass_regNext_20_1_is_stationary_14;
  reg        [15:0]   io_in_c_bypass_regNext_20_2_data_14;
  reg                 io_in_c_bypass_regNext_20_2_is_stationary_14;
  reg        [15:0]   io_in_c_bypass_regNext_20_3_data_14;
  reg                 io_in_c_bypass_regNext_20_3_is_stationary_14;
  reg        [15:0]   io_in_c_bypass_regNext_21_0_data_14;
  reg                 io_in_c_bypass_regNext_21_0_is_stationary_14;
  reg        [15:0]   io_in_c_bypass_regNext_21_1_data_14;
  reg                 io_in_c_bypass_regNext_21_1_is_stationary_14;
  reg        [15:0]   io_in_c_bypass_regNext_21_2_data_14;
  reg                 io_in_c_bypass_regNext_21_2_is_stationary_14;
  reg        [15:0]   io_in_c_bypass_regNext_21_3_data_14;
  reg                 io_in_c_bypass_regNext_21_3_is_stationary_14;
  reg        [15:0]   io_in_c_bypass_regNext_22_0_data_14;
  reg                 io_in_c_bypass_regNext_22_0_is_stationary_14;
  reg        [15:0]   io_in_c_bypass_regNext_22_1_data_14;
  reg                 io_in_c_bypass_regNext_22_1_is_stationary_14;
  reg        [15:0]   io_in_c_bypass_regNext_22_2_data_14;
  reg                 io_in_c_bypass_regNext_22_2_is_stationary_14;
  reg        [15:0]   io_in_c_bypass_regNext_22_3_data_14;
  reg                 io_in_c_bypass_regNext_22_3_is_stationary_14;
  reg        [15:0]   io_in_c_bypass_regNext_23_0_data_14;
  reg                 io_in_c_bypass_regNext_23_0_is_stationary_14;
  reg        [15:0]   io_in_c_bypass_regNext_23_1_data_14;
  reg                 io_in_c_bypass_regNext_23_1_is_stationary_14;
  reg        [15:0]   io_in_c_bypass_regNext_23_2_data_14;
  reg                 io_in_c_bypass_regNext_23_2_is_stationary_14;
  reg        [15:0]   io_in_c_bypass_regNext_23_3_data_14;
  reg                 io_in_c_bypass_regNext_23_3_is_stationary_14;
  reg        [15:0]   io_in_c_bypass_regNext_24_0_data_14;
  reg                 io_in_c_bypass_regNext_24_0_is_stationary_14;
  reg        [15:0]   io_in_c_bypass_regNext_24_1_data_14;
  reg                 io_in_c_bypass_regNext_24_1_is_stationary_14;
  reg        [15:0]   io_in_c_bypass_regNext_24_2_data_14;
  reg                 io_in_c_bypass_regNext_24_2_is_stationary_14;
  reg        [15:0]   io_in_c_bypass_regNext_24_3_data_14;
  reg                 io_in_c_bypass_regNext_24_3_is_stationary_14;
  reg        [15:0]   io_in_c_bypass_regNext_25_0_data_14;
  reg                 io_in_c_bypass_regNext_25_0_is_stationary_14;
  reg        [15:0]   io_in_c_bypass_regNext_25_1_data_14;
  reg                 io_in_c_bypass_regNext_25_1_is_stationary_14;
  reg        [15:0]   io_in_c_bypass_regNext_25_2_data_14;
  reg                 io_in_c_bypass_regNext_25_2_is_stationary_14;
  reg        [15:0]   io_in_c_bypass_regNext_25_3_data_14;
  reg                 io_in_c_bypass_regNext_25_3_is_stationary_14;
  reg        [15:0]   io_in_c_bypass_regNext_26_0_data_14;
  reg                 io_in_c_bypass_regNext_26_0_is_stationary_14;
  reg        [15:0]   io_in_c_bypass_regNext_26_1_data_14;
  reg                 io_in_c_bypass_regNext_26_1_is_stationary_14;
  reg        [15:0]   io_in_c_bypass_regNext_26_2_data_14;
  reg                 io_in_c_bypass_regNext_26_2_is_stationary_14;
  reg        [15:0]   io_in_c_bypass_regNext_26_3_data_14;
  reg                 io_in_c_bypass_regNext_26_3_is_stationary_14;
  reg        [15:0]   io_in_c_bypass_regNext_27_0_data_14;
  reg                 io_in_c_bypass_regNext_27_0_is_stationary_14;
  reg        [15:0]   io_in_c_bypass_regNext_27_1_data_14;
  reg                 io_in_c_bypass_regNext_27_1_is_stationary_14;
  reg        [15:0]   io_in_c_bypass_regNext_27_2_data_14;
  reg                 io_in_c_bypass_regNext_27_2_is_stationary_14;
  reg        [15:0]   io_in_c_bypass_regNext_27_3_data_14;
  reg                 io_in_c_bypass_regNext_27_3_is_stationary_14;
  reg        [15:0]   io_in_c_bypass_regNext_28_0_data_14;
  reg                 io_in_c_bypass_regNext_28_0_is_stationary_14;
  reg        [15:0]   io_in_c_bypass_regNext_28_1_data_14;
  reg                 io_in_c_bypass_regNext_28_1_is_stationary_14;
  reg        [15:0]   io_in_c_bypass_regNext_28_2_data_14;
  reg                 io_in_c_bypass_regNext_28_2_is_stationary_14;
  reg        [15:0]   io_in_c_bypass_regNext_28_3_data_14;
  reg                 io_in_c_bypass_regNext_28_3_is_stationary_14;
  reg        [15:0]   io_in_c_bypass_regNext_29_0_data_14;
  reg                 io_in_c_bypass_regNext_29_0_is_stationary_14;
  reg        [15:0]   io_in_c_bypass_regNext_29_1_data_14;
  reg                 io_in_c_bypass_regNext_29_1_is_stationary_14;
  reg        [15:0]   io_in_c_bypass_regNext_29_2_data_14;
  reg                 io_in_c_bypass_regNext_29_2_is_stationary_14;
  reg        [15:0]   io_in_c_bypass_regNext_29_3_data_14;
  reg                 io_in_c_bypass_regNext_29_3_is_stationary_14;
  reg        [15:0]   io_in_c_bypass_regNext_30_0_data_14;
  reg                 io_in_c_bypass_regNext_30_0_is_stationary_14;
  reg        [15:0]   io_in_c_bypass_regNext_30_1_data_14;
  reg                 io_in_c_bypass_regNext_30_1_is_stationary_14;
  reg        [15:0]   io_in_c_bypass_regNext_30_2_data_14;
  reg                 io_in_c_bypass_regNext_30_2_is_stationary_14;
  reg        [15:0]   io_in_c_bypass_regNext_30_3_data_14;
  reg                 io_in_c_bypass_regNext_30_3_is_stationary_14;
  reg        [15:0]   io_in_c_bypass_regNext_31_0_data_14;
  reg                 io_in_c_bypass_regNext_31_0_is_stationary_14;
  reg        [15:0]   io_in_c_bypass_regNext_31_1_data_14;
  reg                 io_in_c_bypass_regNext_31_1_is_stationary_14;
  reg        [15:0]   io_in_c_bypass_regNext_31_2_data_14;
  reg                 io_in_c_bypass_regNext_31_2_is_stationary_14;
  reg        [15:0]   io_in_c_bypass_regNext_31_3_data_14;
  reg                 io_in_c_bypass_regNext_31_3_is_stationary_14;
  reg        [15:0]   io_in_c_bypass_regNext_0_0_data_15;
  reg                 io_in_c_bypass_regNext_0_0_is_stationary_15;
  reg        [15:0]   io_in_c_bypass_regNext_0_1_data_15;
  reg                 io_in_c_bypass_regNext_0_1_is_stationary_15;
  reg        [15:0]   io_in_c_bypass_regNext_0_2_data_15;
  reg                 io_in_c_bypass_regNext_0_2_is_stationary_15;
  reg        [15:0]   io_in_c_bypass_regNext_0_3_data_15;
  reg                 io_in_c_bypass_regNext_0_3_is_stationary_15;
  reg        [15:0]   io_in_c_bypass_regNext_1_0_data_15;
  reg                 io_in_c_bypass_regNext_1_0_is_stationary_15;
  reg        [15:0]   io_in_c_bypass_regNext_1_1_data_15;
  reg                 io_in_c_bypass_regNext_1_1_is_stationary_15;
  reg        [15:0]   io_in_c_bypass_regNext_1_2_data_15;
  reg                 io_in_c_bypass_regNext_1_2_is_stationary_15;
  reg        [15:0]   io_in_c_bypass_regNext_1_3_data_15;
  reg                 io_in_c_bypass_regNext_1_3_is_stationary_15;
  reg        [15:0]   io_in_c_bypass_regNext_2_0_data_15;
  reg                 io_in_c_bypass_regNext_2_0_is_stationary_15;
  reg        [15:0]   io_in_c_bypass_regNext_2_1_data_15;
  reg                 io_in_c_bypass_regNext_2_1_is_stationary_15;
  reg        [15:0]   io_in_c_bypass_regNext_2_2_data_15;
  reg                 io_in_c_bypass_regNext_2_2_is_stationary_15;
  reg        [15:0]   io_in_c_bypass_regNext_2_3_data_15;
  reg                 io_in_c_bypass_regNext_2_3_is_stationary_15;
  reg        [15:0]   io_in_c_bypass_regNext_3_0_data_15;
  reg                 io_in_c_bypass_regNext_3_0_is_stationary_15;
  reg        [15:0]   io_in_c_bypass_regNext_3_1_data_15;
  reg                 io_in_c_bypass_regNext_3_1_is_stationary_15;
  reg        [15:0]   io_in_c_bypass_regNext_3_2_data_15;
  reg                 io_in_c_bypass_regNext_3_2_is_stationary_15;
  reg        [15:0]   io_in_c_bypass_regNext_3_3_data_15;
  reg                 io_in_c_bypass_regNext_3_3_is_stationary_15;
  reg        [15:0]   io_in_c_bypass_regNext_4_0_data_15;
  reg                 io_in_c_bypass_regNext_4_0_is_stationary_15;
  reg        [15:0]   io_in_c_bypass_regNext_4_1_data_15;
  reg                 io_in_c_bypass_regNext_4_1_is_stationary_15;
  reg        [15:0]   io_in_c_bypass_regNext_4_2_data_15;
  reg                 io_in_c_bypass_regNext_4_2_is_stationary_15;
  reg        [15:0]   io_in_c_bypass_regNext_4_3_data_15;
  reg                 io_in_c_bypass_regNext_4_3_is_stationary_15;
  reg        [15:0]   io_in_c_bypass_regNext_5_0_data_15;
  reg                 io_in_c_bypass_regNext_5_0_is_stationary_15;
  reg        [15:0]   io_in_c_bypass_regNext_5_1_data_15;
  reg                 io_in_c_bypass_regNext_5_1_is_stationary_15;
  reg        [15:0]   io_in_c_bypass_regNext_5_2_data_15;
  reg                 io_in_c_bypass_regNext_5_2_is_stationary_15;
  reg        [15:0]   io_in_c_bypass_regNext_5_3_data_15;
  reg                 io_in_c_bypass_regNext_5_3_is_stationary_15;
  reg        [15:0]   io_in_c_bypass_regNext_6_0_data_15;
  reg                 io_in_c_bypass_regNext_6_0_is_stationary_15;
  reg        [15:0]   io_in_c_bypass_regNext_6_1_data_15;
  reg                 io_in_c_bypass_regNext_6_1_is_stationary_15;
  reg        [15:0]   io_in_c_bypass_regNext_6_2_data_15;
  reg                 io_in_c_bypass_regNext_6_2_is_stationary_15;
  reg        [15:0]   io_in_c_bypass_regNext_6_3_data_15;
  reg                 io_in_c_bypass_regNext_6_3_is_stationary_15;
  reg        [15:0]   io_in_c_bypass_regNext_7_0_data_15;
  reg                 io_in_c_bypass_regNext_7_0_is_stationary_15;
  reg        [15:0]   io_in_c_bypass_regNext_7_1_data_15;
  reg                 io_in_c_bypass_regNext_7_1_is_stationary_15;
  reg        [15:0]   io_in_c_bypass_regNext_7_2_data_15;
  reg                 io_in_c_bypass_regNext_7_2_is_stationary_15;
  reg        [15:0]   io_in_c_bypass_regNext_7_3_data_15;
  reg                 io_in_c_bypass_regNext_7_3_is_stationary_15;
  reg        [15:0]   io_in_c_bypass_regNext_8_0_data_15;
  reg                 io_in_c_bypass_regNext_8_0_is_stationary_15;
  reg        [15:0]   io_in_c_bypass_regNext_8_1_data_15;
  reg                 io_in_c_bypass_regNext_8_1_is_stationary_15;
  reg        [15:0]   io_in_c_bypass_regNext_8_2_data_15;
  reg                 io_in_c_bypass_regNext_8_2_is_stationary_15;
  reg        [15:0]   io_in_c_bypass_regNext_8_3_data_15;
  reg                 io_in_c_bypass_regNext_8_3_is_stationary_15;
  reg        [15:0]   io_in_c_bypass_regNext_9_0_data_15;
  reg                 io_in_c_bypass_regNext_9_0_is_stationary_15;
  reg        [15:0]   io_in_c_bypass_regNext_9_1_data_15;
  reg                 io_in_c_bypass_regNext_9_1_is_stationary_15;
  reg        [15:0]   io_in_c_bypass_regNext_9_2_data_15;
  reg                 io_in_c_bypass_regNext_9_2_is_stationary_15;
  reg        [15:0]   io_in_c_bypass_regNext_9_3_data_15;
  reg                 io_in_c_bypass_regNext_9_3_is_stationary_15;
  reg        [15:0]   io_in_c_bypass_regNext_10_0_data_15;
  reg                 io_in_c_bypass_regNext_10_0_is_stationary_15;
  reg        [15:0]   io_in_c_bypass_regNext_10_1_data_15;
  reg                 io_in_c_bypass_regNext_10_1_is_stationary_15;
  reg        [15:0]   io_in_c_bypass_regNext_10_2_data_15;
  reg                 io_in_c_bypass_regNext_10_2_is_stationary_15;
  reg        [15:0]   io_in_c_bypass_regNext_10_3_data_15;
  reg                 io_in_c_bypass_regNext_10_3_is_stationary_15;
  reg        [15:0]   io_in_c_bypass_regNext_11_0_data_15;
  reg                 io_in_c_bypass_regNext_11_0_is_stationary_15;
  reg        [15:0]   io_in_c_bypass_regNext_11_1_data_15;
  reg                 io_in_c_bypass_regNext_11_1_is_stationary_15;
  reg        [15:0]   io_in_c_bypass_regNext_11_2_data_15;
  reg                 io_in_c_bypass_regNext_11_2_is_stationary_15;
  reg        [15:0]   io_in_c_bypass_regNext_11_3_data_15;
  reg                 io_in_c_bypass_regNext_11_3_is_stationary_15;
  reg        [15:0]   io_in_c_bypass_regNext_12_0_data_15;
  reg                 io_in_c_bypass_regNext_12_0_is_stationary_15;
  reg        [15:0]   io_in_c_bypass_regNext_12_1_data_15;
  reg                 io_in_c_bypass_regNext_12_1_is_stationary_15;
  reg        [15:0]   io_in_c_bypass_regNext_12_2_data_15;
  reg                 io_in_c_bypass_regNext_12_2_is_stationary_15;
  reg        [15:0]   io_in_c_bypass_regNext_12_3_data_15;
  reg                 io_in_c_bypass_regNext_12_3_is_stationary_15;
  reg        [15:0]   io_in_c_bypass_regNext_13_0_data_15;
  reg                 io_in_c_bypass_regNext_13_0_is_stationary_15;
  reg        [15:0]   io_in_c_bypass_regNext_13_1_data_15;
  reg                 io_in_c_bypass_regNext_13_1_is_stationary_15;
  reg        [15:0]   io_in_c_bypass_regNext_13_2_data_15;
  reg                 io_in_c_bypass_regNext_13_2_is_stationary_15;
  reg        [15:0]   io_in_c_bypass_regNext_13_3_data_15;
  reg                 io_in_c_bypass_regNext_13_3_is_stationary_15;
  reg        [15:0]   io_in_c_bypass_regNext_14_0_data_15;
  reg                 io_in_c_bypass_regNext_14_0_is_stationary_15;
  reg        [15:0]   io_in_c_bypass_regNext_14_1_data_15;
  reg                 io_in_c_bypass_regNext_14_1_is_stationary_15;
  reg        [15:0]   io_in_c_bypass_regNext_14_2_data_15;
  reg                 io_in_c_bypass_regNext_14_2_is_stationary_15;
  reg        [15:0]   io_in_c_bypass_regNext_14_3_data_15;
  reg                 io_in_c_bypass_regNext_14_3_is_stationary_15;
  reg        [15:0]   io_in_c_bypass_regNext_15_0_data_15;
  reg                 io_in_c_bypass_regNext_15_0_is_stationary_15;
  reg        [15:0]   io_in_c_bypass_regNext_15_1_data_15;
  reg                 io_in_c_bypass_regNext_15_1_is_stationary_15;
  reg        [15:0]   io_in_c_bypass_regNext_15_2_data_15;
  reg                 io_in_c_bypass_regNext_15_2_is_stationary_15;
  reg        [15:0]   io_in_c_bypass_regNext_15_3_data_15;
  reg                 io_in_c_bypass_regNext_15_3_is_stationary_15;
  reg        [15:0]   io_in_c_bypass_regNext_16_0_data_15;
  reg                 io_in_c_bypass_regNext_16_0_is_stationary_15;
  reg        [15:0]   io_in_c_bypass_regNext_16_1_data_15;
  reg                 io_in_c_bypass_regNext_16_1_is_stationary_15;
  reg        [15:0]   io_in_c_bypass_regNext_16_2_data_15;
  reg                 io_in_c_bypass_regNext_16_2_is_stationary_15;
  reg        [15:0]   io_in_c_bypass_regNext_16_3_data_15;
  reg                 io_in_c_bypass_regNext_16_3_is_stationary_15;
  reg        [15:0]   io_in_c_bypass_regNext_17_0_data_15;
  reg                 io_in_c_bypass_regNext_17_0_is_stationary_15;
  reg        [15:0]   io_in_c_bypass_regNext_17_1_data_15;
  reg                 io_in_c_bypass_regNext_17_1_is_stationary_15;
  reg        [15:0]   io_in_c_bypass_regNext_17_2_data_15;
  reg                 io_in_c_bypass_regNext_17_2_is_stationary_15;
  reg        [15:0]   io_in_c_bypass_regNext_17_3_data_15;
  reg                 io_in_c_bypass_regNext_17_3_is_stationary_15;
  reg        [15:0]   io_in_c_bypass_regNext_18_0_data_15;
  reg                 io_in_c_bypass_regNext_18_0_is_stationary_15;
  reg        [15:0]   io_in_c_bypass_regNext_18_1_data_15;
  reg                 io_in_c_bypass_regNext_18_1_is_stationary_15;
  reg        [15:0]   io_in_c_bypass_regNext_18_2_data_15;
  reg                 io_in_c_bypass_regNext_18_2_is_stationary_15;
  reg        [15:0]   io_in_c_bypass_regNext_18_3_data_15;
  reg                 io_in_c_bypass_regNext_18_3_is_stationary_15;
  reg        [15:0]   io_in_c_bypass_regNext_19_0_data_15;
  reg                 io_in_c_bypass_regNext_19_0_is_stationary_15;
  reg        [15:0]   io_in_c_bypass_regNext_19_1_data_15;
  reg                 io_in_c_bypass_regNext_19_1_is_stationary_15;
  reg        [15:0]   io_in_c_bypass_regNext_19_2_data_15;
  reg                 io_in_c_bypass_regNext_19_2_is_stationary_15;
  reg        [15:0]   io_in_c_bypass_regNext_19_3_data_15;
  reg                 io_in_c_bypass_regNext_19_3_is_stationary_15;
  reg        [15:0]   io_in_c_bypass_regNext_20_0_data_15;
  reg                 io_in_c_bypass_regNext_20_0_is_stationary_15;
  reg        [15:0]   io_in_c_bypass_regNext_20_1_data_15;
  reg                 io_in_c_bypass_regNext_20_1_is_stationary_15;
  reg        [15:0]   io_in_c_bypass_regNext_20_2_data_15;
  reg                 io_in_c_bypass_regNext_20_2_is_stationary_15;
  reg        [15:0]   io_in_c_bypass_regNext_20_3_data_15;
  reg                 io_in_c_bypass_regNext_20_3_is_stationary_15;
  reg        [15:0]   io_in_c_bypass_regNext_21_0_data_15;
  reg                 io_in_c_bypass_regNext_21_0_is_stationary_15;
  reg        [15:0]   io_in_c_bypass_regNext_21_1_data_15;
  reg                 io_in_c_bypass_regNext_21_1_is_stationary_15;
  reg        [15:0]   io_in_c_bypass_regNext_21_2_data_15;
  reg                 io_in_c_bypass_regNext_21_2_is_stationary_15;
  reg        [15:0]   io_in_c_bypass_regNext_21_3_data_15;
  reg                 io_in_c_bypass_regNext_21_3_is_stationary_15;
  reg        [15:0]   io_in_c_bypass_regNext_22_0_data_15;
  reg                 io_in_c_bypass_regNext_22_0_is_stationary_15;
  reg        [15:0]   io_in_c_bypass_regNext_22_1_data_15;
  reg                 io_in_c_bypass_regNext_22_1_is_stationary_15;
  reg        [15:0]   io_in_c_bypass_regNext_22_2_data_15;
  reg                 io_in_c_bypass_regNext_22_2_is_stationary_15;
  reg        [15:0]   io_in_c_bypass_regNext_22_3_data_15;
  reg                 io_in_c_bypass_regNext_22_3_is_stationary_15;
  reg        [15:0]   io_in_c_bypass_regNext_23_0_data_15;
  reg                 io_in_c_bypass_regNext_23_0_is_stationary_15;
  reg        [15:0]   io_in_c_bypass_regNext_23_1_data_15;
  reg                 io_in_c_bypass_regNext_23_1_is_stationary_15;
  reg        [15:0]   io_in_c_bypass_regNext_23_2_data_15;
  reg                 io_in_c_bypass_regNext_23_2_is_stationary_15;
  reg        [15:0]   io_in_c_bypass_regNext_23_3_data_15;
  reg                 io_in_c_bypass_regNext_23_3_is_stationary_15;
  reg        [15:0]   io_in_c_bypass_regNext_24_0_data_15;
  reg                 io_in_c_bypass_regNext_24_0_is_stationary_15;
  reg        [15:0]   io_in_c_bypass_regNext_24_1_data_15;
  reg                 io_in_c_bypass_regNext_24_1_is_stationary_15;
  reg        [15:0]   io_in_c_bypass_regNext_24_2_data_15;
  reg                 io_in_c_bypass_regNext_24_2_is_stationary_15;
  reg        [15:0]   io_in_c_bypass_regNext_24_3_data_15;
  reg                 io_in_c_bypass_regNext_24_3_is_stationary_15;
  reg        [15:0]   io_in_c_bypass_regNext_25_0_data_15;
  reg                 io_in_c_bypass_regNext_25_0_is_stationary_15;
  reg        [15:0]   io_in_c_bypass_regNext_25_1_data_15;
  reg                 io_in_c_bypass_regNext_25_1_is_stationary_15;
  reg        [15:0]   io_in_c_bypass_regNext_25_2_data_15;
  reg                 io_in_c_bypass_regNext_25_2_is_stationary_15;
  reg        [15:0]   io_in_c_bypass_regNext_25_3_data_15;
  reg                 io_in_c_bypass_regNext_25_3_is_stationary_15;
  reg        [15:0]   io_in_c_bypass_regNext_26_0_data_15;
  reg                 io_in_c_bypass_regNext_26_0_is_stationary_15;
  reg        [15:0]   io_in_c_bypass_regNext_26_1_data_15;
  reg                 io_in_c_bypass_regNext_26_1_is_stationary_15;
  reg        [15:0]   io_in_c_bypass_regNext_26_2_data_15;
  reg                 io_in_c_bypass_regNext_26_2_is_stationary_15;
  reg        [15:0]   io_in_c_bypass_regNext_26_3_data_15;
  reg                 io_in_c_bypass_regNext_26_3_is_stationary_15;
  reg        [15:0]   io_in_c_bypass_regNext_27_0_data_15;
  reg                 io_in_c_bypass_regNext_27_0_is_stationary_15;
  reg        [15:0]   io_in_c_bypass_regNext_27_1_data_15;
  reg                 io_in_c_bypass_regNext_27_1_is_stationary_15;
  reg        [15:0]   io_in_c_bypass_regNext_27_2_data_15;
  reg                 io_in_c_bypass_regNext_27_2_is_stationary_15;
  reg        [15:0]   io_in_c_bypass_regNext_27_3_data_15;
  reg                 io_in_c_bypass_regNext_27_3_is_stationary_15;
  reg        [15:0]   io_in_c_bypass_regNext_28_0_data_15;
  reg                 io_in_c_bypass_regNext_28_0_is_stationary_15;
  reg        [15:0]   io_in_c_bypass_regNext_28_1_data_15;
  reg                 io_in_c_bypass_regNext_28_1_is_stationary_15;
  reg        [15:0]   io_in_c_bypass_regNext_28_2_data_15;
  reg                 io_in_c_bypass_regNext_28_2_is_stationary_15;
  reg        [15:0]   io_in_c_bypass_regNext_28_3_data_15;
  reg                 io_in_c_bypass_regNext_28_3_is_stationary_15;
  reg        [15:0]   io_in_c_bypass_regNext_29_0_data_15;
  reg                 io_in_c_bypass_regNext_29_0_is_stationary_15;
  reg        [15:0]   io_in_c_bypass_regNext_29_1_data_15;
  reg                 io_in_c_bypass_regNext_29_1_is_stationary_15;
  reg        [15:0]   io_in_c_bypass_regNext_29_2_data_15;
  reg                 io_in_c_bypass_regNext_29_2_is_stationary_15;
  reg        [15:0]   io_in_c_bypass_regNext_29_3_data_15;
  reg                 io_in_c_bypass_regNext_29_3_is_stationary_15;
  reg        [15:0]   io_in_c_bypass_regNext_30_0_data_15;
  reg                 io_in_c_bypass_regNext_30_0_is_stationary_15;
  reg        [15:0]   io_in_c_bypass_regNext_30_1_data_15;
  reg                 io_in_c_bypass_regNext_30_1_is_stationary_15;
  reg        [15:0]   io_in_c_bypass_regNext_30_2_data_15;
  reg                 io_in_c_bypass_regNext_30_2_is_stationary_15;
  reg        [15:0]   io_in_c_bypass_regNext_30_3_data_15;
  reg                 io_in_c_bypass_regNext_30_3_is_stationary_15;
  reg        [15:0]   io_in_c_bypass_regNext_31_0_data_15;
  reg                 io_in_c_bypass_regNext_31_0_is_stationary_15;
  reg        [15:0]   io_in_c_bypass_regNext_31_1_data_15;
  reg                 io_in_c_bypass_regNext_31_1_is_stationary_15;
  reg        [15:0]   io_in_c_bypass_regNext_31_2_data_15;
  reg                 io_in_c_bypass_regNext_31_2_is_stationary_15;
  reg        [15:0]   io_in_c_bypass_regNext_31_3_data_15;
  reg                 io_in_c_bypass_regNext_31_3_is_stationary_15;
  reg        [15:0]   io_in_c_bypass_regNext_0_0_data_16;
  reg                 io_in_c_bypass_regNext_0_0_is_stationary_16;
  reg        [15:0]   io_in_c_bypass_regNext_0_1_data_16;
  reg                 io_in_c_bypass_regNext_0_1_is_stationary_16;
  reg        [15:0]   io_in_c_bypass_regNext_0_2_data_16;
  reg                 io_in_c_bypass_regNext_0_2_is_stationary_16;
  reg        [15:0]   io_in_c_bypass_regNext_0_3_data_16;
  reg                 io_in_c_bypass_regNext_0_3_is_stationary_16;
  reg        [15:0]   io_in_c_bypass_regNext_1_0_data_16;
  reg                 io_in_c_bypass_regNext_1_0_is_stationary_16;
  reg        [15:0]   io_in_c_bypass_regNext_1_1_data_16;
  reg                 io_in_c_bypass_regNext_1_1_is_stationary_16;
  reg        [15:0]   io_in_c_bypass_regNext_1_2_data_16;
  reg                 io_in_c_bypass_regNext_1_2_is_stationary_16;
  reg        [15:0]   io_in_c_bypass_regNext_1_3_data_16;
  reg                 io_in_c_bypass_regNext_1_3_is_stationary_16;
  reg        [15:0]   io_in_c_bypass_regNext_2_0_data_16;
  reg                 io_in_c_bypass_regNext_2_0_is_stationary_16;
  reg        [15:0]   io_in_c_bypass_regNext_2_1_data_16;
  reg                 io_in_c_bypass_regNext_2_1_is_stationary_16;
  reg        [15:0]   io_in_c_bypass_regNext_2_2_data_16;
  reg                 io_in_c_bypass_regNext_2_2_is_stationary_16;
  reg        [15:0]   io_in_c_bypass_regNext_2_3_data_16;
  reg                 io_in_c_bypass_regNext_2_3_is_stationary_16;
  reg        [15:0]   io_in_c_bypass_regNext_3_0_data_16;
  reg                 io_in_c_bypass_regNext_3_0_is_stationary_16;
  reg        [15:0]   io_in_c_bypass_regNext_3_1_data_16;
  reg                 io_in_c_bypass_regNext_3_1_is_stationary_16;
  reg        [15:0]   io_in_c_bypass_regNext_3_2_data_16;
  reg                 io_in_c_bypass_regNext_3_2_is_stationary_16;
  reg        [15:0]   io_in_c_bypass_regNext_3_3_data_16;
  reg                 io_in_c_bypass_regNext_3_3_is_stationary_16;
  reg        [15:0]   io_in_c_bypass_regNext_4_0_data_16;
  reg                 io_in_c_bypass_regNext_4_0_is_stationary_16;
  reg        [15:0]   io_in_c_bypass_regNext_4_1_data_16;
  reg                 io_in_c_bypass_regNext_4_1_is_stationary_16;
  reg        [15:0]   io_in_c_bypass_regNext_4_2_data_16;
  reg                 io_in_c_bypass_regNext_4_2_is_stationary_16;
  reg        [15:0]   io_in_c_bypass_regNext_4_3_data_16;
  reg                 io_in_c_bypass_regNext_4_3_is_stationary_16;
  reg        [15:0]   io_in_c_bypass_regNext_5_0_data_16;
  reg                 io_in_c_bypass_regNext_5_0_is_stationary_16;
  reg        [15:0]   io_in_c_bypass_regNext_5_1_data_16;
  reg                 io_in_c_bypass_regNext_5_1_is_stationary_16;
  reg        [15:0]   io_in_c_bypass_regNext_5_2_data_16;
  reg                 io_in_c_bypass_regNext_5_2_is_stationary_16;
  reg        [15:0]   io_in_c_bypass_regNext_5_3_data_16;
  reg                 io_in_c_bypass_regNext_5_3_is_stationary_16;
  reg        [15:0]   io_in_c_bypass_regNext_6_0_data_16;
  reg                 io_in_c_bypass_regNext_6_0_is_stationary_16;
  reg        [15:0]   io_in_c_bypass_regNext_6_1_data_16;
  reg                 io_in_c_bypass_regNext_6_1_is_stationary_16;
  reg        [15:0]   io_in_c_bypass_regNext_6_2_data_16;
  reg                 io_in_c_bypass_regNext_6_2_is_stationary_16;
  reg        [15:0]   io_in_c_bypass_regNext_6_3_data_16;
  reg                 io_in_c_bypass_regNext_6_3_is_stationary_16;
  reg        [15:0]   io_in_c_bypass_regNext_7_0_data_16;
  reg                 io_in_c_bypass_regNext_7_0_is_stationary_16;
  reg        [15:0]   io_in_c_bypass_regNext_7_1_data_16;
  reg                 io_in_c_bypass_regNext_7_1_is_stationary_16;
  reg        [15:0]   io_in_c_bypass_regNext_7_2_data_16;
  reg                 io_in_c_bypass_regNext_7_2_is_stationary_16;
  reg        [15:0]   io_in_c_bypass_regNext_7_3_data_16;
  reg                 io_in_c_bypass_regNext_7_3_is_stationary_16;
  reg        [15:0]   io_in_c_bypass_regNext_8_0_data_16;
  reg                 io_in_c_bypass_regNext_8_0_is_stationary_16;
  reg        [15:0]   io_in_c_bypass_regNext_8_1_data_16;
  reg                 io_in_c_bypass_regNext_8_1_is_stationary_16;
  reg        [15:0]   io_in_c_bypass_regNext_8_2_data_16;
  reg                 io_in_c_bypass_regNext_8_2_is_stationary_16;
  reg        [15:0]   io_in_c_bypass_regNext_8_3_data_16;
  reg                 io_in_c_bypass_regNext_8_3_is_stationary_16;
  reg        [15:0]   io_in_c_bypass_regNext_9_0_data_16;
  reg                 io_in_c_bypass_regNext_9_0_is_stationary_16;
  reg        [15:0]   io_in_c_bypass_regNext_9_1_data_16;
  reg                 io_in_c_bypass_regNext_9_1_is_stationary_16;
  reg        [15:0]   io_in_c_bypass_regNext_9_2_data_16;
  reg                 io_in_c_bypass_regNext_9_2_is_stationary_16;
  reg        [15:0]   io_in_c_bypass_regNext_9_3_data_16;
  reg                 io_in_c_bypass_regNext_9_3_is_stationary_16;
  reg        [15:0]   io_in_c_bypass_regNext_10_0_data_16;
  reg                 io_in_c_bypass_regNext_10_0_is_stationary_16;
  reg        [15:0]   io_in_c_bypass_regNext_10_1_data_16;
  reg                 io_in_c_bypass_regNext_10_1_is_stationary_16;
  reg        [15:0]   io_in_c_bypass_regNext_10_2_data_16;
  reg                 io_in_c_bypass_regNext_10_2_is_stationary_16;
  reg        [15:0]   io_in_c_bypass_regNext_10_3_data_16;
  reg                 io_in_c_bypass_regNext_10_3_is_stationary_16;
  reg        [15:0]   io_in_c_bypass_regNext_11_0_data_16;
  reg                 io_in_c_bypass_regNext_11_0_is_stationary_16;
  reg        [15:0]   io_in_c_bypass_regNext_11_1_data_16;
  reg                 io_in_c_bypass_regNext_11_1_is_stationary_16;
  reg        [15:0]   io_in_c_bypass_regNext_11_2_data_16;
  reg                 io_in_c_bypass_regNext_11_2_is_stationary_16;
  reg        [15:0]   io_in_c_bypass_regNext_11_3_data_16;
  reg                 io_in_c_bypass_regNext_11_3_is_stationary_16;
  reg        [15:0]   io_in_c_bypass_regNext_12_0_data_16;
  reg                 io_in_c_bypass_regNext_12_0_is_stationary_16;
  reg        [15:0]   io_in_c_bypass_regNext_12_1_data_16;
  reg                 io_in_c_bypass_regNext_12_1_is_stationary_16;
  reg        [15:0]   io_in_c_bypass_regNext_12_2_data_16;
  reg                 io_in_c_bypass_regNext_12_2_is_stationary_16;
  reg        [15:0]   io_in_c_bypass_regNext_12_3_data_16;
  reg                 io_in_c_bypass_regNext_12_3_is_stationary_16;
  reg        [15:0]   io_in_c_bypass_regNext_13_0_data_16;
  reg                 io_in_c_bypass_regNext_13_0_is_stationary_16;
  reg        [15:0]   io_in_c_bypass_regNext_13_1_data_16;
  reg                 io_in_c_bypass_regNext_13_1_is_stationary_16;
  reg        [15:0]   io_in_c_bypass_regNext_13_2_data_16;
  reg                 io_in_c_bypass_regNext_13_2_is_stationary_16;
  reg        [15:0]   io_in_c_bypass_regNext_13_3_data_16;
  reg                 io_in_c_bypass_regNext_13_3_is_stationary_16;
  reg        [15:0]   io_in_c_bypass_regNext_14_0_data_16;
  reg                 io_in_c_bypass_regNext_14_0_is_stationary_16;
  reg        [15:0]   io_in_c_bypass_regNext_14_1_data_16;
  reg                 io_in_c_bypass_regNext_14_1_is_stationary_16;
  reg        [15:0]   io_in_c_bypass_regNext_14_2_data_16;
  reg                 io_in_c_bypass_regNext_14_2_is_stationary_16;
  reg        [15:0]   io_in_c_bypass_regNext_14_3_data_16;
  reg                 io_in_c_bypass_regNext_14_3_is_stationary_16;
  reg        [15:0]   io_in_c_bypass_regNext_15_0_data_16;
  reg                 io_in_c_bypass_regNext_15_0_is_stationary_16;
  reg        [15:0]   io_in_c_bypass_regNext_15_1_data_16;
  reg                 io_in_c_bypass_regNext_15_1_is_stationary_16;
  reg        [15:0]   io_in_c_bypass_regNext_15_2_data_16;
  reg                 io_in_c_bypass_regNext_15_2_is_stationary_16;
  reg        [15:0]   io_in_c_bypass_regNext_15_3_data_16;
  reg                 io_in_c_bypass_regNext_15_3_is_stationary_16;
  reg        [15:0]   io_in_c_bypass_regNext_16_0_data_16;
  reg                 io_in_c_bypass_regNext_16_0_is_stationary_16;
  reg        [15:0]   io_in_c_bypass_regNext_16_1_data_16;
  reg                 io_in_c_bypass_regNext_16_1_is_stationary_16;
  reg        [15:0]   io_in_c_bypass_regNext_16_2_data_16;
  reg                 io_in_c_bypass_regNext_16_2_is_stationary_16;
  reg        [15:0]   io_in_c_bypass_regNext_16_3_data_16;
  reg                 io_in_c_bypass_regNext_16_3_is_stationary_16;
  reg        [15:0]   io_in_c_bypass_regNext_17_0_data_16;
  reg                 io_in_c_bypass_regNext_17_0_is_stationary_16;
  reg        [15:0]   io_in_c_bypass_regNext_17_1_data_16;
  reg                 io_in_c_bypass_regNext_17_1_is_stationary_16;
  reg        [15:0]   io_in_c_bypass_regNext_17_2_data_16;
  reg                 io_in_c_bypass_regNext_17_2_is_stationary_16;
  reg        [15:0]   io_in_c_bypass_regNext_17_3_data_16;
  reg                 io_in_c_bypass_regNext_17_3_is_stationary_16;
  reg        [15:0]   io_in_c_bypass_regNext_18_0_data_16;
  reg                 io_in_c_bypass_regNext_18_0_is_stationary_16;
  reg        [15:0]   io_in_c_bypass_regNext_18_1_data_16;
  reg                 io_in_c_bypass_regNext_18_1_is_stationary_16;
  reg        [15:0]   io_in_c_bypass_regNext_18_2_data_16;
  reg                 io_in_c_bypass_regNext_18_2_is_stationary_16;
  reg        [15:0]   io_in_c_bypass_regNext_18_3_data_16;
  reg                 io_in_c_bypass_regNext_18_3_is_stationary_16;
  reg        [15:0]   io_in_c_bypass_regNext_19_0_data_16;
  reg                 io_in_c_bypass_regNext_19_0_is_stationary_16;
  reg        [15:0]   io_in_c_bypass_regNext_19_1_data_16;
  reg                 io_in_c_bypass_regNext_19_1_is_stationary_16;
  reg        [15:0]   io_in_c_bypass_regNext_19_2_data_16;
  reg                 io_in_c_bypass_regNext_19_2_is_stationary_16;
  reg        [15:0]   io_in_c_bypass_regNext_19_3_data_16;
  reg                 io_in_c_bypass_regNext_19_3_is_stationary_16;
  reg        [15:0]   io_in_c_bypass_regNext_20_0_data_16;
  reg                 io_in_c_bypass_regNext_20_0_is_stationary_16;
  reg        [15:0]   io_in_c_bypass_regNext_20_1_data_16;
  reg                 io_in_c_bypass_regNext_20_1_is_stationary_16;
  reg        [15:0]   io_in_c_bypass_regNext_20_2_data_16;
  reg                 io_in_c_bypass_regNext_20_2_is_stationary_16;
  reg        [15:0]   io_in_c_bypass_regNext_20_3_data_16;
  reg                 io_in_c_bypass_regNext_20_3_is_stationary_16;
  reg        [15:0]   io_in_c_bypass_regNext_21_0_data_16;
  reg                 io_in_c_bypass_regNext_21_0_is_stationary_16;
  reg        [15:0]   io_in_c_bypass_regNext_21_1_data_16;
  reg                 io_in_c_bypass_regNext_21_1_is_stationary_16;
  reg        [15:0]   io_in_c_bypass_regNext_21_2_data_16;
  reg                 io_in_c_bypass_regNext_21_2_is_stationary_16;
  reg        [15:0]   io_in_c_bypass_regNext_21_3_data_16;
  reg                 io_in_c_bypass_regNext_21_3_is_stationary_16;
  reg        [15:0]   io_in_c_bypass_regNext_22_0_data_16;
  reg                 io_in_c_bypass_regNext_22_0_is_stationary_16;
  reg        [15:0]   io_in_c_bypass_regNext_22_1_data_16;
  reg                 io_in_c_bypass_regNext_22_1_is_stationary_16;
  reg        [15:0]   io_in_c_bypass_regNext_22_2_data_16;
  reg                 io_in_c_bypass_regNext_22_2_is_stationary_16;
  reg        [15:0]   io_in_c_bypass_regNext_22_3_data_16;
  reg                 io_in_c_bypass_regNext_22_3_is_stationary_16;
  reg        [15:0]   io_in_c_bypass_regNext_23_0_data_16;
  reg                 io_in_c_bypass_regNext_23_0_is_stationary_16;
  reg        [15:0]   io_in_c_bypass_regNext_23_1_data_16;
  reg                 io_in_c_bypass_regNext_23_1_is_stationary_16;
  reg        [15:0]   io_in_c_bypass_regNext_23_2_data_16;
  reg                 io_in_c_bypass_regNext_23_2_is_stationary_16;
  reg        [15:0]   io_in_c_bypass_regNext_23_3_data_16;
  reg                 io_in_c_bypass_regNext_23_3_is_stationary_16;
  reg        [15:0]   io_in_c_bypass_regNext_24_0_data_16;
  reg                 io_in_c_bypass_regNext_24_0_is_stationary_16;
  reg        [15:0]   io_in_c_bypass_regNext_24_1_data_16;
  reg                 io_in_c_bypass_regNext_24_1_is_stationary_16;
  reg        [15:0]   io_in_c_bypass_regNext_24_2_data_16;
  reg                 io_in_c_bypass_regNext_24_2_is_stationary_16;
  reg        [15:0]   io_in_c_bypass_regNext_24_3_data_16;
  reg                 io_in_c_bypass_regNext_24_3_is_stationary_16;
  reg        [15:0]   io_in_c_bypass_regNext_25_0_data_16;
  reg                 io_in_c_bypass_regNext_25_0_is_stationary_16;
  reg        [15:0]   io_in_c_bypass_regNext_25_1_data_16;
  reg                 io_in_c_bypass_regNext_25_1_is_stationary_16;
  reg        [15:0]   io_in_c_bypass_regNext_25_2_data_16;
  reg                 io_in_c_bypass_regNext_25_2_is_stationary_16;
  reg        [15:0]   io_in_c_bypass_regNext_25_3_data_16;
  reg                 io_in_c_bypass_regNext_25_3_is_stationary_16;
  reg        [15:0]   io_in_c_bypass_regNext_26_0_data_16;
  reg                 io_in_c_bypass_regNext_26_0_is_stationary_16;
  reg        [15:0]   io_in_c_bypass_regNext_26_1_data_16;
  reg                 io_in_c_bypass_regNext_26_1_is_stationary_16;
  reg        [15:0]   io_in_c_bypass_regNext_26_2_data_16;
  reg                 io_in_c_bypass_regNext_26_2_is_stationary_16;
  reg        [15:0]   io_in_c_bypass_regNext_26_3_data_16;
  reg                 io_in_c_bypass_regNext_26_3_is_stationary_16;
  reg        [15:0]   io_in_c_bypass_regNext_27_0_data_16;
  reg                 io_in_c_bypass_regNext_27_0_is_stationary_16;
  reg        [15:0]   io_in_c_bypass_regNext_27_1_data_16;
  reg                 io_in_c_bypass_regNext_27_1_is_stationary_16;
  reg        [15:0]   io_in_c_bypass_regNext_27_2_data_16;
  reg                 io_in_c_bypass_regNext_27_2_is_stationary_16;
  reg        [15:0]   io_in_c_bypass_regNext_27_3_data_16;
  reg                 io_in_c_bypass_regNext_27_3_is_stationary_16;
  reg        [15:0]   io_in_c_bypass_regNext_28_0_data_16;
  reg                 io_in_c_bypass_regNext_28_0_is_stationary_16;
  reg        [15:0]   io_in_c_bypass_regNext_28_1_data_16;
  reg                 io_in_c_bypass_regNext_28_1_is_stationary_16;
  reg        [15:0]   io_in_c_bypass_regNext_28_2_data_16;
  reg                 io_in_c_bypass_regNext_28_2_is_stationary_16;
  reg        [15:0]   io_in_c_bypass_regNext_28_3_data_16;
  reg                 io_in_c_bypass_regNext_28_3_is_stationary_16;
  reg        [15:0]   io_in_c_bypass_regNext_29_0_data_16;
  reg                 io_in_c_bypass_regNext_29_0_is_stationary_16;
  reg        [15:0]   io_in_c_bypass_regNext_29_1_data_16;
  reg                 io_in_c_bypass_regNext_29_1_is_stationary_16;
  reg        [15:0]   io_in_c_bypass_regNext_29_2_data_16;
  reg                 io_in_c_bypass_regNext_29_2_is_stationary_16;
  reg        [15:0]   io_in_c_bypass_regNext_29_3_data_16;
  reg                 io_in_c_bypass_regNext_29_3_is_stationary_16;
  reg        [15:0]   io_in_c_bypass_regNext_30_0_data_16;
  reg                 io_in_c_bypass_regNext_30_0_is_stationary_16;
  reg        [15:0]   io_in_c_bypass_regNext_30_1_data_16;
  reg                 io_in_c_bypass_regNext_30_1_is_stationary_16;
  reg        [15:0]   io_in_c_bypass_regNext_30_2_data_16;
  reg                 io_in_c_bypass_regNext_30_2_is_stationary_16;
  reg        [15:0]   io_in_c_bypass_regNext_30_3_data_16;
  reg                 io_in_c_bypass_regNext_30_3_is_stationary_16;
  reg        [15:0]   io_in_c_bypass_regNext_31_0_data_16;
  reg                 io_in_c_bypass_regNext_31_0_is_stationary_16;
  reg        [15:0]   io_in_c_bypass_regNext_31_1_data_16;
  reg                 io_in_c_bypass_regNext_31_1_is_stationary_16;
  reg        [15:0]   io_in_c_bypass_regNext_31_2_data_16;
  reg                 io_in_c_bypass_regNext_31_2_is_stationary_16;
  reg        [15:0]   io_in_c_bypass_regNext_31_3_data_16;
  reg                 io_in_c_bypass_regNext_31_3_is_stationary_16;
  reg        [15:0]   io_in_c_bypass_regNext_0_0_data_17;
  reg                 io_in_c_bypass_regNext_0_0_is_stationary_17;
  reg        [15:0]   io_in_c_bypass_regNext_0_1_data_17;
  reg                 io_in_c_bypass_regNext_0_1_is_stationary_17;
  reg        [15:0]   io_in_c_bypass_regNext_0_2_data_17;
  reg                 io_in_c_bypass_regNext_0_2_is_stationary_17;
  reg        [15:0]   io_in_c_bypass_regNext_0_3_data_17;
  reg                 io_in_c_bypass_regNext_0_3_is_stationary_17;
  reg        [15:0]   io_in_c_bypass_regNext_1_0_data_17;
  reg                 io_in_c_bypass_regNext_1_0_is_stationary_17;
  reg        [15:0]   io_in_c_bypass_regNext_1_1_data_17;
  reg                 io_in_c_bypass_regNext_1_1_is_stationary_17;
  reg        [15:0]   io_in_c_bypass_regNext_1_2_data_17;
  reg                 io_in_c_bypass_regNext_1_2_is_stationary_17;
  reg        [15:0]   io_in_c_bypass_regNext_1_3_data_17;
  reg                 io_in_c_bypass_regNext_1_3_is_stationary_17;
  reg        [15:0]   io_in_c_bypass_regNext_2_0_data_17;
  reg                 io_in_c_bypass_regNext_2_0_is_stationary_17;
  reg        [15:0]   io_in_c_bypass_regNext_2_1_data_17;
  reg                 io_in_c_bypass_regNext_2_1_is_stationary_17;
  reg        [15:0]   io_in_c_bypass_regNext_2_2_data_17;
  reg                 io_in_c_bypass_regNext_2_2_is_stationary_17;
  reg        [15:0]   io_in_c_bypass_regNext_2_3_data_17;
  reg                 io_in_c_bypass_regNext_2_3_is_stationary_17;
  reg        [15:0]   io_in_c_bypass_regNext_3_0_data_17;
  reg                 io_in_c_bypass_regNext_3_0_is_stationary_17;
  reg        [15:0]   io_in_c_bypass_regNext_3_1_data_17;
  reg                 io_in_c_bypass_regNext_3_1_is_stationary_17;
  reg        [15:0]   io_in_c_bypass_regNext_3_2_data_17;
  reg                 io_in_c_bypass_regNext_3_2_is_stationary_17;
  reg        [15:0]   io_in_c_bypass_regNext_3_3_data_17;
  reg                 io_in_c_bypass_regNext_3_3_is_stationary_17;
  reg        [15:0]   io_in_c_bypass_regNext_4_0_data_17;
  reg                 io_in_c_bypass_regNext_4_0_is_stationary_17;
  reg        [15:0]   io_in_c_bypass_regNext_4_1_data_17;
  reg                 io_in_c_bypass_regNext_4_1_is_stationary_17;
  reg        [15:0]   io_in_c_bypass_regNext_4_2_data_17;
  reg                 io_in_c_bypass_regNext_4_2_is_stationary_17;
  reg        [15:0]   io_in_c_bypass_regNext_4_3_data_17;
  reg                 io_in_c_bypass_regNext_4_3_is_stationary_17;
  reg        [15:0]   io_in_c_bypass_regNext_5_0_data_17;
  reg                 io_in_c_bypass_regNext_5_0_is_stationary_17;
  reg        [15:0]   io_in_c_bypass_regNext_5_1_data_17;
  reg                 io_in_c_bypass_regNext_5_1_is_stationary_17;
  reg        [15:0]   io_in_c_bypass_regNext_5_2_data_17;
  reg                 io_in_c_bypass_regNext_5_2_is_stationary_17;
  reg        [15:0]   io_in_c_bypass_regNext_5_3_data_17;
  reg                 io_in_c_bypass_regNext_5_3_is_stationary_17;
  reg        [15:0]   io_in_c_bypass_regNext_6_0_data_17;
  reg                 io_in_c_bypass_regNext_6_0_is_stationary_17;
  reg        [15:0]   io_in_c_bypass_regNext_6_1_data_17;
  reg                 io_in_c_bypass_regNext_6_1_is_stationary_17;
  reg        [15:0]   io_in_c_bypass_regNext_6_2_data_17;
  reg                 io_in_c_bypass_regNext_6_2_is_stationary_17;
  reg        [15:0]   io_in_c_bypass_regNext_6_3_data_17;
  reg                 io_in_c_bypass_regNext_6_3_is_stationary_17;
  reg        [15:0]   io_in_c_bypass_regNext_7_0_data_17;
  reg                 io_in_c_bypass_regNext_7_0_is_stationary_17;
  reg        [15:0]   io_in_c_bypass_regNext_7_1_data_17;
  reg                 io_in_c_bypass_regNext_7_1_is_stationary_17;
  reg        [15:0]   io_in_c_bypass_regNext_7_2_data_17;
  reg                 io_in_c_bypass_regNext_7_2_is_stationary_17;
  reg        [15:0]   io_in_c_bypass_regNext_7_3_data_17;
  reg                 io_in_c_bypass_regNext_7_3_is_stationary_17;
  reg        [15:0]   io_in_c_bypass_regNext_8_0_data_17;
  reg                 io_in_c_bypass_regNext_8_0_is_stationary_17;
  reg        [15:0]   io_in_c_bypass_regNext_8_1_data_17;
  reg                 io_in_c_bypass_regNext_8_1_is_stationary_17;
  reg        [15:0]   io_in_c_bypass_regNext_8_2_data_17;
  reg                 io_in_c_bypass_regNext_8_2_is_stationary_17;
  reg        [15:0]   io_in_c_bypass_regNext_8_3_data_17;
  reg                 io_in_c_bypass_regNext_8_3_is_stationary_17;
  reg        [15:0]   io_in_c_bypass_regNext_9_0_data_17;
  reg                 io_in_c_bypass_regNext_9_0_is_stationary_17;
  reg        [15:0]   io_in_c_bypass_regNext_9_1_data_17;
  reg                 io_in_c_bypass_regNext_9_1_is_stationary_17;
  reg        [15:0]   io_in_c_bypass_regNext_9_2_data_17;
  reg                 io_in_c_bypass_regNext_9_2_is_stationary_17;
  reg        [15:0]   io_in_c_bypass_regNext_9_3_data_17;
  reg                 io_in_c_bypass_regNext_9_3_is_stationary_17;
  reg        [15:0]   io_in_c_bypass_regNext_10_0_data_17;
  reg                 io_in_c_bypass_regNext_10_0_is_stationary_17;
  reg        [15:0]   io_in_c_bypass_regNext_10_1_data_17;
  reg                 io_in_c_bypass_regNext_10_1_is_stationary_17;
  reg        [15:0]   io_in_c_bypass_regNext_10_2_data_17;
  reg                 io_in_c_bypass_regNext_10_2_is_stationary_17;
  reg        [15:0]   io_in_c_bypass_regNext_10_3_data_17;
  reg                 io_in_c_bypass_regNext_10_3_is_stationary_17;
  reg        [15:0]   io_in_c_bypass_regNext_11_0_data_17;
  reg                 io_in_c_bypass_regNext_11_0_is_stationary_17;
  reg        [15:0]   io_in_c_bypass_regNext_11_1_data_17;
  reg                 io_in_c_bypass_regNext_11_1_is_stationary_17;
  reg        [15:0]   io_in_c_bypass_regNext_11_2_data_17;
  reg                 io_in_c_bypass_regNext_11_2_is_stationary_17;
  reg        [15:0]   io_in_c_bypass_regNext_11_3_data_17;
  reg                 io_in_c_bypass_regNext_11_3_is_stationary_17;
  reg        [15:0]   io_in_c_bypass_regNext_12_0_data_17;
  reg                 io_in_c_bypass_regNext_12_0_is_stationary_17;
  reg        [15:0]   io_in_c_bypass_regNext_12_1_data_17;
  reg                 io_in_c_bypass_regNext_12_1_is_stationary_17;
  reg        [15:0]   io_in_c_bypass_regNext_12_2_data_17;
  reg                 io_in_c_bypass_regNext_12_2_is_stationary_17;
  reg        [15:0]   io_in_c_bypass_regNext_12_3_data_17;
  reg                 io_in_c_bypass_regNext_12_3_is_stationary_17;
  reg        [15:0]   io_in_c_bypass_regNext_13_0_data_17;
  reg                 io_in_c_bypass_regNext_13_0_is_stationary_17;
  reg        [15:0]   io_in_c_bypass_regNext_13_1_data_17;
  reg                 io_in_c_bypass_regNext_13_1_is_stationary_17;
  reg        [15:0]   io_in_c_bypass_regNext_13_2_data_17;
  reg                 io_in_c_bypass_regNext_13_2_is_stationary_17;
  reg        [15:0]   io_in_c_bypass_regNext_13_3_data_17;
  reg                 io_in_c_bypass_regNext_13_3_is_stationary_17;
  reg        [15:0]   io_in_c_bypass_regNext_14_0_data_17;
  reg                 io_in_c_bypass_regNext_14_0_is_stationary_17;
  reg        [15:0]   io_in_c_bypass_regNext_14_1_data_17;
  reg                 io_in_c_bypass_regNext_14_1_is_stationary_17;
  reg        [15:0]   io_in_c_bypass_regNext_14_2_data_17;
  reg                 io_in_c_bypass_regNext_14_2_is_stationary_17;
  reg        [15:0]   io_in_c_bypass_regNext_14_3_data_17;
  reg                 io_in_c_bypass_regNext_14_3_is_stationary_17;
  reg        [15:0]   io_in_c_bypass_regNext_15_0_data_17;
  reg                 io_in_c_bypass_regNext_15_0_is_stationary_17;
  reg        [15:0]   io_in_c_bypass_regNext_15_1_data_17;
  reg                 io_in_c_bypass_regNext_15_1_is_stationary_17;
  reg        [15:0]   io_in_c_bypass_regNext_15_2_data_17;
  reg                 io_in_c_bypass_regNext_15_2_is_stationary_17;
  reg        [15:0]   io_in_c_bypass_regNext_15_3_data_17;
  reg                 io_in_c_bypass_regNext_15_3_is_stationary_17;
  reg        [15:0]   io_in_c_bypass_regNext_16_0_data_17;
  reg                 io_in_c_bypass_regNext_16_0_is_stationary_17;
  reg        [15:0]   io_in_c_bypass_regNext_16_1_data_17;
  reg                 io_in_c_bypass_regNext_16_1_is_stationary_17;
  reg        [15:0]   io_in_c_bypass_regNext_16_2_data_17;
  reg                 io_in_c_bypass_regNext_16_2_is_stationary_17;
  reg        [15:0]   io_in_c_bypass_regNext_16_3_data_17;
  reg                 io_in_c_bypass_regNext_16_3_is_stationary_17;
  reg        [15:0]   io_in_c_bypass_regNext_17_0_data_17;
  reg                 io_in_c_bypass_regNext_17_0_is_stationary_17;
  reg        [15:0]   io_in_c_bypass_regNext_17_1_data_17;
  reg                 io_in_c_bypass_regNext_17_1_is_stationary_17;
  reg        [15:0]   io_in_c_bypass_regNext_17_2_data_17;
  reg                 io_in_c_bypass_regNext_17_2_is_stationary_17;
  reg        [15:0]   io_in_c_bypass_regNext_17_3_data_17;
  reg                 io_in_c_bypass_regNext_17_3_is_stationary_17;
  reg        [15:0]   io_in_c_bypass_regNext_18_0_data_17;
  reg                 io_in_c_bypass_regNext_18_0_is_stationary_17;
  reg        [15:0]   io_in_c_bypass_regNext_18_1_data_17;
  reg                 io_in_c_bypass_regNext_18_1_is_stationary_17;
  reg        [15:0]   io_in_c_bypass_regNext_18_2_data_17;
  reg                 io_in_c_bypass_regNext_18_2_is_stationary_17;
  reg        [15:0]   io_in_c_bypass_regNext_18_3_data_17;
  reg                 io_in_c_bypass_regNext_18_3_is_stationary_17;
  reg        [15:0]   io_in_c_bypass_regNext_19_0_data_17;
  reg                 io_in_c_bypass_regNext_19_0_is_stationary_17;
  reg        [15:0]   io_in_c_bypass_regNext_19_1_data_17;
  reg                 io_in_c_bypass_regNext_19_1_is_stationary_17;
  reg        [15:0]   io_in_c_bypass_regNext_19_2_data_17;
  reg                 io_in_c_bypass_regNext_19_2_is_stationary_17;
  reg        [15:0]   io_in_c_bypass_regNext_19_3_data_17;
  reg                 io_in_c_bypass_regNext_19_3_is_stationary_17;
  reg        [15:0]   io_in_c_bypass_regNext_20_0_data_17;
  reg                 io_in_c_bypass_regNext_20_0_is_stationary_17;
  reg        [15:0]   io_in_c_bypass_regNext_20_1_data_17;
  reg                 io_in_c_bypass_regNext_20_1_is_stationary_17;
  reg        [15:0]   io_in_c_bypass_regNext_20_2_data_17;
  reg                 io_in_c_bypass_regNext_20_2_is_stationary_17;
  reg        [15:0]   io_in_c_bypass_regNext_20_3_data_17;
  reg                 io_in_c_bypass_regNext_20_3_is_stationary_17;
  reg        [15:0]   io_in_c_bypass_regNext_21_0_data_17;
  reg                 io_in_c_bypass_regNext_21_0_is_stationary_17;
  reg        [15:0]   io_in_c_bypass_regNext_21_1_data_17;
  reg                 io_in_c_bypass_regNext_21_1_is_stationary_17;
  reg        [15:0]   io_in_c_bypass_regNext_21_2_data_17;
  reg                 io_in_c_bypass_regNext_21_2_is_stationary_17;
  reg        [15:0]   io_in_c_bypass_regNext_21_3_data_17;
  reg                 io_in_c_bypass_regNext_21_3_is_stationary_17;
  reg        [15:0]   io_in_c_bypass_regNext_22_0_data_17;
  reg                 io_in_c_bypass_regNext_22_0_is_stationary_17;
  reg        [15:0]   io_in_c_bypass_regNext_22_1_data_17;
  reg                 io_in_c_bypass_regNext_22_1_is_stationary_17;
  reg        [15:0]   io_in_c_bypass_regNext_22_2_data_17;
  reg                 io_in_c_bypass_regNext_22_2_is_stationary_17;
  reg        [15:0]   io_in_c_bypass_regNext_22_3_data_17;
  reg                 io_in_c_bypass_regNext_22_3_is_stationary_17;
  reg        [15:0]   io_in_c_bypass_regNext_23_0_data_17;
  reg                 io_in_c_bypass_regNext_23_0_is_stationary_17;
  reg        [15:0]   io_in_c_bypass_regNext_23_1_data_17;
  reg                 io_in_c_bypass_regNext_23_1_is_stationary_17;
  reg        [15:0]   io_in_c_bypass_regNext_23_2_data_17;
  reg                 io_in_c_bypass_regNext_23_2_is_stationary_17;
  reg        [15:0]   io_in_c_bypass_regNext_23_3_data_17;
  reg                 io_in_c_bypass_regNext_23_3_is_stationary_17;
  reg        [15:0]   io_in_c_bypass_regNext_24_0_data_17;
  reg                 io_in_c_bypass_regNext_24_0_is_stationary_17;
  reg        [15:0]   io_in_c_bypass_regNext_24_1_data_17;
  reg                 io_in_c_bypass_regNext_24_1_is_stationary_17;
  reg        [15:0]   io_in_c_bypass_regNext_24_2_data_17;
  reg                 io_in_c_bypass_regNext_24_2_is_stationary_17;
  reg        [15:0]   io_in_c_bypass_regNext_24_3_data_17;
  reg                 io_in_c_bypass_regNext_24_3_is_stationary_17;
  reg        [15:0]   io_in_c_bypass_regNext_25_0_data_17;
  reg                 io_in_c_bypass_regNext_25_0_is_stationary_17;
  reg        [15:0]   io_in_c_bypass_regNext_25_1_data_17;
  reg                 io_in_c_bypass_regNext_25_1_is_stationary_17;
  reg        [15:0]   io_in_c_bypass_regNext_25_2_data_17;
  reg                 io_in_c_bypass_regNext_25_2_is_stationary_17;
  reg        [15:0]   io_in_c_bypass_regNext_25_3_data_17;
  reg                 io_in_c_bypass_regNext_25_3_is_stationary_17;
  reg        [15:0]   io_in_c_bypass_regNext_26_0_data_17;
  reg                 io_in_c_bypass_regNext_26_0_is_stationary_17;
  reg        [15:0]   io_in_c_bypass_regNext_26_1_data_17;
  reg                 io_in_c_bypass_regNext_26_1_is_stationary_17;
  reg        [15:0]   io_in_c_bypass_regNext_26_2_data_17;
  reg                 io_in_c_bypass_regNext_26_2_is_stationary_17;
  reg        [15:0]   io_in_c_bypass_regNext_26_3_data_17;
  reg                 io_in_c_bypass_regNext_26_3_is_stationary_17;
  reg        [15:0]   io_in_c_bypass_regNext_27_0_data_17;
  reg                 io_in_c_bypass_regNext_27_0_is_stationary_17;
  reg        [15:0]   io_in_c_bypass_regNext_27_1_data_17;
  reg                 io_in_c_bypass_regNext_27_1_is_stationary_17;
  reg        [15:0]   io_in_c_bypass_regNext_27_2_data_17;
  reg                 io_in_c_bypass_regNext_27_2_is_stationary_17;
  reg        [15:0]   io_in_c_bypass_regNext_27_3_data_17;
  reg                 io_in_c_bypass_regNext_27_3_is_stationary_17;
  reg        [15:0]   io_in_c_bypass_regNext_28_0_data_17;
  reg                 io_in_c_bypass_regNext_28_0_is_stationary_17;
  reg        [15:0]   io_in_c_bypass_regNext_28_1_data_17;
  reg                 io_in_c_bypass_regNext_28_1_is_stationary_17;
  reg        [15:0]   io_in_c_bypass_regNext_28_2_data_17;
  reg                 io_in_c_bypass_regNext_28_2_is_stationary_17;
  reg        [15:0]   io_in_c_bypass_regNext_28_3_data_17;
  reg                 io_in_c_bypass_regNext_28_3_is_stationary_17;
  reg        [15:0]   io_in_c_bypass_regNext_29_0_data_17;
  reg                 io_in_c_bypass_regNext_29_0_is_stationary_17;
  reg        [15:0]   io_in_c_bypass_regNext_29_1_data_17;
  reg                 io_in_c_bypass_regNext_29_1_is_stationary_17;
  reg        [15:0]   io_in_c_bypass_regNext_29_2_data_17;
  reg                 io_in_c_bypass_regNext_29_2_is_stationary_17;
  reg        [15:0]   io_in_c_bypass_regNext_29_3_data_17;
  reg                 io_in_c_bypass_regNext_29_3_is_stationary_17;
  reg        [15:0]   io_in_c_bypass_regNext_30_0_data_17;
  reg                 io_in_c_bypass_regNext_30_0_is_stationary_17;
  reg        [15:0]   io_in_c_bypass_regNext_30_1_data_17;
  reg                 io_in_c_bypass_regNext_30_1_is_stationary_17;
  reg        [15:0]   io_in_c_bypass_regNext_30_2_data_17;
  reg                 io_in_c_bypass_regNext_30_2_is_stationary_17;
  reg        [15:0]   io_in_c_bypass_regNext_30_3_data_17;
  reg                 io_in_c_bypass_regNext_30_3_is_stationary_17;
  reg        [15:0]   io_in_c_bypass_regNext_31_0_data_17;
  reg                 io_in_c_bypass_regNext_31_0_is_stationary_17;
  reg        [15:0]   io_in_c_bypass_regNext_31_1_data_17;
  reg                 io_in_c_bypass_regNext_31_1_is_stationary_17;
  reg        [15:0]   io_in_c_bypass_regNext_31_2_data_17;
  reg                 io_in_c_bypass_regNext_31_2_is_stationary_17;
  reg        [15:0]   io_in_c_bypass_regNext_31_3_data_17;
  reg                 io_in_c_bypass_regNext_31_3_is_stationary_17;
  reg        [15:0]   io_in_c_bypass_regNext_0_0_data_18;
  reg                 io_in_c_bypass_regNext_0_0_is_stationary_18;
  reg        [15:0]   io_in_c_bypass_regNext_0_1_data_18;
  reg                 io_in_c_bypass_regNext_0_1_is_stationary_18;
  reg        [15:0]   io_in_c_bypass_regNext_0_2_data_18;
  reg                 io_in_c_bypass_regNext_0_2_is_stationary_18;
  reg        [15:0]   io_in_c_bypass_regNext_0_3_data_18;
  reg                 io_in_c_bypass_regNext_0_3_is_stationary_18;
  reg        [15:0]   io_in_c_bypass_regNext_1_0_data_18;
  reg                 io_in_c_bypass_regNext_1_0_is_stationary_18;
  reg        [15:0]   io_in_c_bypass_regNext_1_1_data_18;
  reg                 io_in_c_bypass_regNext_1_1_is_stationary_18;
  reg        [15:0]   io_in_c_bypass_regNext_1_2_data_18;
  reg                 io_in_c_bypass_regNext_1_2_is_stationary_18;
  reg        [15:0]   io_in_c_bypass_regNext_1_3_data_18;
  reg                 io_in_c_bypass_regNext_1_3_is_stationary_18;
  reg        [15:0]   io_in_c_bypass_regNext_2_0_data_18;
  reg                 io_in_c_bypass_regNext_2_0_is_stationary_18;
  reg        [15:0]   io_in_c_bypass_regNext_2_1_data_18;
  reg                 io_in_c_bypass_regNext_2_1_is_stationary_18;
  reg        [15:0]   io_in_c_bypass_regNext_2_2_data_18;
  reg                 io_in_c_bypass_regNext_2_2_is_stationary_18;
  reg        [15:0]   io_in_c_bypass_regNext_2_3_data_18;
  reg                 io_in_c_bypass_regNext_2_3_is_stationary_18;
  reg        [15:0]   io_in_c_bypass_regNext_3_0_data_18;
  reg                 io_in_c_bypass_regNext_3_0_is_stationary_18;
  reg        [15:0]   io_in_c_bypass_regNext_3_1_data_18;
  reg                 io_in_c_bypass_regNext_3_1_is_stationary_18;
  reg        [15:0]   io_in_c_bypass_regNext_3_2_data_18;
  reg                 io_in_c_bypass_regNext_3_2_is_stationary_18;
  reg        [15:0]   io_in_c_bypass_regNext_3_3_data_18;
  reg                 io_in_c_bypass_regNext_3_3_is_stationary_18;
  reg        [15:0]   io_in_c_bypass_regNext_4_0_data_18;
  reg                 io_in_c_bypass_regNext_4_0_is_stationary_18;
  reg        [15:0]   io_in_c_bypass_regNext_4_1_data_18;
  reg                 io_in_c_bypass_regNext_4_1_is_stationary_18;
  reg        [15:0]   io_in_c_bypass_regNext_4_2_data_18;
  reg                 io_in_c_bypass_regNext_4_2_is_stationary_18;
  reg        [15:0]   io_in_c_bypass_regNext_4_3_data_18;
  reg                 io_in_c_bypass_regNext_4_3_is_stationary_18;
  reg        [15:0]   io_in_c_bypass_regNext_5_0_data_18;
  reg                 io_in_c_bypass_regNext_5_0_is_stationary_18;
  reg        [15:0]   io_in_c_bypass_regNext_5_1_data_18;
  reg                 io_in_c_bypass_regNext_5_1_is_stationary_18;
  reg        [15:0]   io_in_c_bypass_regNext_5_2_data_18;
  reg                 io_in_c_bypass_regNext_5_2_is_stationary_18;
  reg        [15:0]   io_in_c_bypass_regNext_5_3_data_18;
  reg                 io_in_c_bypass_regNext_5_3_is_stationary_18;
  reg        [15:0]   io_in_c_bypass_regNext_6_0_data_18;
  reg                 io_in_c_bypass_regNext_6_0_is_stationary_18;
  reg        [15:0]   io_in_c_bypass_regNext_6_1_data_18;
  reg                 io_in_c_bypass_regNext_6_1_is_stationary_18;
  reg        [15:0]   io_in_c_bypass_regNext_6_2_data_18;
  reg                 io_in_c_bypass_regNext_6_2_is_stationary_18;
  reg        [15:0]   io_in_c_bypass_regNext_6_3_data_18;
  reg                 io_in_c_bypass_regNext_6_3_is_stationary_18;
  reg        [15:0]   io_in_c_bypass_regNext_7_0_data_18;
  reg                 io_in_c_bypass_regNext_7_0_is_stationary_18;
  reg        [15:0]   io_in_c_bypass_regNext_7_1_data_18;
  reg                 io_in_c_bypass_regNext_7_1_is_stationary_18;
  reg        [15:0]   io_in_c_bypass_regNext_7_2_data_18;
  reg                 io_in_c_bypass_regNext_7_2_is_stationary_18;
  reg        [15:0]   io_in_c_bypass_regNext_7_3_data_18;
  reg                 io_in_c_bypass_regNext_7_3_is_stationary_18;
  reg        [15:0]   io_in_c_bypass_regNext_8_0_data_18;
  reg                 io_in_c_bypass_regNext_8_0_is_stationary_18;
  reg        [15:0]   io_in_c_bypass_regNext_8_1_data_18;
  reg                 io_in_c_bypass_regNext_8_1_is_stationary_18;
  reg        [15:0]   io_in_c_bypass_regNext_8_2_data_18;
  reg                 io_in_c_bypass_regNext_8_2_is_stationary_18;
  reg        [15:0]   io_in_c_bypass_regNext_8_3_data_18;
  reg                 io_in_c_bypass_regNext_8_3_is_stationary_18;
  reg        [15:0]   io_in_c_bypass_regNext_9_0_data_18;
  reg                 io_in_c_bypass_regNext_9_0_is_stationary_18;
  reg        [15:0]   io_in_c_bypass_regNext_9_1_data_18;
  reg                 io_in_c_bypass_regNext_9_1_is_stationary_18;
  reg        [15:0]   io_in_c_bypass_regNext_9_2_data_18;
  reg                 io_in_c_bypass_regNext_9_2_is_stationary_18;
  reg        [15:0]   io_in_c_bypass_regNext_9_3_data_18;
  reg                 io_in_c_bypass_regNext_9_3_is_stationary_18;
  reg        [15:0]   io_in_c_bypass_regNext_10_0_data_18;
  reg                 io_in_c_bypass_regNext_10_0_is_stationary_18;
  reg        [15:0]   io_in_c_bypass_regNext_10_1_data_18;
  reg                 io_in_c_bypass_regNext_10_1_is_stationary_18;
  reg        [15:0]   io_in_c_bypass_regNext_10_2_data_18;
  reg                 io_in_c_bypass_regNext_10_2_is_stationary_18;
  reg        [15:0]   io_in_c_bypass_regNext_10_3_data_18;
  reg                 io_in_c_bypass_regNext_10_3_is_stationary_18;
  reg        [15:0]   io_in_c_bypass_regNext_11_0_data_18;
  reg                 io_in_c_bypass_regNext_11_0_is_stationary_18;
  reg        [15:0]   io_in_c_bypass_regNext_11_1_data_18;
  reg                 io_in_c_bypass_regNext_11_1_is_stationary_18;
  reg        [15:0]   io_in_c_bypass_regNext_11_2_data_18;
  reg                 io_in_c_bypass_regNext_11_2_is_stationary_18;
  reg        [15:0]   io_in_c_bypass_regNext_11_3_data_18;
  reg                 io_in_c_bypass_regNext_11_3_is_stationary_18;
  reg        [15:0]   io_in_c_bypass_regNext_12_0_data_18;
  reg                 io_in_c_bypass_regNext_12_0_is_stationary_18;
  reg        [15:0]   io_in_c_bypass_regNext_12_1_data_18;
  reg                 io_in_c_bypass_regNext_12_1_is_stationary_18;
  reg        [15:0]   io_in_c_bypass_regNext_12_2_data_18;
  reg                 io_in_c_bypass_regNext_12_2_is_stationary_18;
  reg        [15:0]   io_in_c_bypass_regNext_12_3_data_18;
  reg                 io_in_c_bypass_regNext_12_3_is_stationary_18;
  reg        [15:0]   io_in_c_bypass_regNext_13_0_data_18;
  reg                 io_in_c_bypass_regNext_13_0_is_stationary_18;
  reg        [15:0]   io_in_c_bypass_regNext_13_1_data_18;
  reg                 io_in_c_bypass_regNext_13_1_is_stationary_18;
  reg        [15:0]   io_in_c_bypass_regNext_13_2_data_18;
  reg                 io_in_c_bypass_regNext_13_2_is_stationary_18;
  reg        [15:0]   io_in_c_bypass_regNext_13_3_data_18;
  reg                 io_in_c_bypass_regNext_13_3_is_stationary_18;
  reg        [15:0]   io_in_c_bypass_regNext_14_0_data_18;
  reg                 io_in_c_bypass_regNext_14_0_is_stationary_18;
  reg        [15:0]   io_in_c_bypass_regNext_14_1_data_18;
  reg                 io_in_c_bypass_regNext_14_1_is_stationary_18;
  reg        [15:0]   io_in_c_bypass_regNext_14_2_data_18;
  reg                 io_in_c_bypass_regNext_14_2_is_stationary_18;
  reg        [15:0]   io_in_c_bypass_regNext_14_3_data_18;
  reg                 io_in_c_bypass_regNext_14_3_is_stationary_18;
  reg        [15:0]   io_in_c_bypass_regNext_15_0_data_18;
  reg                 io_in_c_bypass_regNext_15_0_is_stationary_18;
  reg        [15:0]   io_in_c_bypass_regNext_15_1_data_18;
  reg                 io_in_c_bypass_regNext_15_1_is_stationary_18;
  reg        [15:0]   io_in_c_bypass_regNext_15_2_data_18;
  reg                 io_in_c_bypass_regNext_15_2_is_stationary_18;
  reg        [15:0]   io_in_c_bypass_regNext_15_3_data_18;
  reg                 io_in_c_bypass_regNext_15_3_is_stationary_18;
  reg        [15:0]   io_in_c_bypass_regNext_16_0_data_18;
  reg                 io_in_c_bypass_regNext_16_0_is_stationary_18;
  reg        [15:0]   io_in_c_bypass_regNext_16_1_data_18;
  reg                 io_in_c_bypass_regNext_16_1_is_stationary_18;
  reg        [15:0]   io_in_c_bypass_regNext_16_2_data_18;
  reg                 io_in_c_bypass_regNext_16_2_is_stationary_18;
  reg        [15:0]   io_in_c_bypass_regNext_16_3_data_18;
  reg                 io_in_c_bypass_regNext_16_3_is_stationary_18;
  reg        [15:0]   io_in_c_bypass_regNext_17_0_data_18;
  reg                 io_in_c_bypass_regNext_17_0_is_stationary_18;
  reg        [15:0]   io_in_c_bypass_regNext_17_1_data_18;
  reg                 io_in_c_bypass_regNext_17_1_is_stationary_18;
  reg        [15:0]   io_in_c_bypass_regNext_17_2_data_18;
  reg                 io_in_c_bypass_regNext_17_2_is_stationary_18;
  reg        [15:0]   io_in_c_bypass_regNext_17_3_data_18;
  reg                 io_in_c_bypass_regNext_17_3_is_stationary_18;
  reg        [15:0]   io_in_c_bypass_regNext_18_0_data_18;
  reg                 io_in_c_bypass_regNext_18_0_is_stationary_18;
  reg        [15:0]   io_in_c_bypass_regNext_18_1_data_18;
  reg                 io_in_c_bypass_regNext_18_1_is_stationary_18;
  reg        [15:0]   io_in_c_bypass_regNext_18_2_data_18;
  reg                 io_in_c_bypass_regNext_18_2_is_stationary_18;
  reg        [15:0]   io_in_c_bypass_regNext_18_3_data_18;
  reg                 io_in_c_bypass_regNext_18_3_is_stationary_18;
  reg        [15:0]   io_in_c_bypass_regNext_19_0_data_18;
  reg                 io_in_c_bypass_regNext_19_0_is_stationary_18;
  reg        [15:0]   io_in_c_bypass_regNext_19_1_data_18;
  reg                 io_in_c_bypass_regNext_19_1_is_stationary_18;
  reg        [15:0]   io_in_c_bypass_regNext_19_2_data_18;
  reg                 io_in_c_bypass_regNext_19_2_is_stationary_18;
  reg        [15:0]   io_in_c_bypass_regNext_19_3_data_18;
  reg                 io_in_c_bypass_regNext_19_3_is_stationary_18;
  reg        [15:0]   io_in_c_bypass_regNext_20_0_data_18;
  reg                 io_in_c_bypass_regNext_20_0_is_stationary_18;
  reg        [15:0]   io_in_c_bypass_regNext_20_1_data_18;
  reg                 io_in_c_bypass_regNext_20_1_is_stationary_18;
  reg        [15:0]   io_in_c_bypass_regNext_20_2_data_18;
  reg                 io_in_c_bypass_regNext_20_2_is_stationary_18;
  reg        [15:0]   io_in_c_bypass_regNext_20_3_data_18;
  reg                 io_in_c_bypass_regNext_20_3_is_stationary_18;
  reg        [15:0]   io_in_c_bypass_regNext_21_0_data_18;
  reg                 io_in_c_bypass_regNext_21_0_is_stationary_18;
  reg        [15:0]   io_in_c_bypass_regNext_21_1_data_18;
  reg                 io_in_c_bypass_regNext_21_1_is_stationary_18;
  reg        [15:0]   io_in_c_bypass_regNext_21_2_data_18;
  reg                 io_in_c_bypass_regNext_21_2_is_stationary_18;
  reg        [15:0]   io_in_c_bypass_regNext_21_3_data_18;
  reg                 io_in_c_bypass_regNext_21_3_is_stationary_18;
  reg        [15:0]   io_in_c_bypass_regNext_22_0_data_18;
  reg                 io_in_c_bypass_regNext_22_0_is_stationary_18;
  reg        [15:0]   io_in_c_bypass_regNext_22_1_data_18;
  reg                 io_in_c_bypass_regNext_22_1_is_stationary_18;
  reg        [15:0]   io_in_c_bypass_regNext_22_2_data_18;
  reg                 io_in_c_bypass_regNext_22_2_is_stationary_18;
  reg        [15:0]   io_in_c_bypass_regNext_22_3_data_18;
  reg                 io_in_c_bypass_regNext_22_3_is_stationary_18;
  reg        [15:0]   io_in_c_bypass_regNext_23_0_data_18;
  reg                 io_in_c_bypass_regNext_23_0_is_stationary_18;
  reg        [15:0]   io_in_c_bypass_regNext_23_1_data_18;
  reg                 io_in_c_bypass_regNext_23_1_is_stationary_18;
  reg        [15:0]   io_in_c_bypass_regNext_23_2_data_18;
  reg                 io_in_c_bypass_regNext_23_2_is_stationary_18;
  reg        [15:0]   io_in_c_bypass_regNext_23_3_data_18;
  reg                 io_in_c_bypass_regNext_23_3_is_stationary_18;
  reg        [15:0]   io_in_c_bypass_regNext_24_0_data_18;
  reg                 io_in_c_bypass_regNext_24_0_is_stationary_18;
  reg        [15:0]   io_in_c_bypass_regNext_24_1_data_18;
  reg                 io_in_c_bypass_regNext_24_1_is_stationary_18;
  reg        [15:0]   io_in_c_bypass_regNext_24_2_data_18;
  reg                 io_in_c_bypass_regNext_24_2_is_stationary_18;
  reg        [15:0]   io_in_c_bypass_regNext_24_3_data_18;
  reg                 io_in_c_bypass_regNext_24_3_is_stationary_18;
  reg        [15:0]   io_in_c_bypass_regNext_25_0_data_18;
  reg                 io_in_c_bypass_regNext_25_0_is_stationary_18;
  reg        [15:0]   io_in_c_bypass_regNext_25_1_data_18;
  reg                 io_in_c_bypass_regNext_25_1_is_stationary_18;
  reg        [15:0]   io_in_c_bypass_regNext_25_2_data_18;
  reg                 io_in_c_bypass_regNext_25_2_is_stationary_18;
  reg        [15:0]   io_in_c_bypass_regNext_25_3_data_18;
  reg                 io_in_c_bypass_regNext_25_3_is_stationary_18;
  reg        [15:0]   io_in_c_bypass_regNext_26_0_data_18;
  reg                 io_in_c_bypass_regNext_26_0_is_stationary_18;
  reg        [15:0]   io_in_c_bypass_regNext_26_1_data_18;
  reg                 io_in_c_bypass_regNext_26_1_is_stationary_18;
  reg        [15:0]   io_in_c_bypass_regNext_26_2_data_18;
  reg                 io_in_c_bypass_regNext_26_2_is_stationary_18;
  reg        [15:0]   io_in_c_bypass_regNext_26_3_data_18;
  reg                 io_in_c_bypass_regNext_26_3_is_stationary_18;
  reg        [15:0]   io_in_c_bypass_regNext_27_0_data_18;
  reg                 io_in_c_bypass_regNext_27_0_is_stationary_18;
  reg        [15:0]   io_in_c_bypass_regNext_27_1_data_18;
  reg                 io_in_c_bypass_regNext_27_1_is_stationary_18;
  reg        [15:0]   io_in_c_bypass_regNext_27_2_data_18;
  reg                 io_in_c_bypass_regNext_27_2_is_stationary_18;
  reg        [15:0]   io_in_c_bypass_regNext_27_3_data_18;
  reg                 io_in_c_bypass_regNext_27_3_is_stationary_18;
  reg        [15:0]   io_in_c_bypass_regNext_28_0_data_18;
  reg                 io_in_c_bypass_regNext_28_0_is_stationary_18;
  reg        [15:0]   io_in_c_bypass_regNext_28_1_data_18;
  reg                 io_in_c_bypass_regNext_28_1_is_stationary_18;
  reg        [15:0]   io_in_c_bypass_regNext_28_2_data_18;
  reg                 io_in_c_bypass_regNext_28_2_is_stationary_18;
  reg        [15:0]   io_in_c_bypass_regNext_28_3_data_18;
  reg                 io_in_c_bypass_regNext_28_3_is_stationary_18;
  reg        [15:0]   io_in_c_bypass_regNext_29_0_data_18;
  reg                 io_in_c_bypass_regNext_29_0_is_stationary_18;
  reg        [15:0]   io_in_c_bypass_regNext_29_1_data_18;
  reg                 io_in_c_bypass_regNext_29_1_is_stationary_18;
  reg        [15:0]   io_in_c_bypass_regNext_29_2_data_18;
  reg                 io_in_c_bypass_regNext_29_2_is_stationary_18;
  reg        [15:0]   io_in_c_bypass_regNext_29_3_data_18;
  reg                 io_in_c_bypass_regNext_29_3_is_stationary_18;
  reg        [15:0]   io_in_c_bypass_regNext_30_0_data_18;
  reg                 io_in_c_bypass_regNext_30_0_is_stationary_18;
  reg        [15:0]   io_in_c_bypass_regNext_30_1_data_18;
  reg                 io_in_c_bypass_regNext_30_1_is_stationary_18;
  reg        [15:0]   io_in_c_bypass_regNext_30_2_data_18;
  reg                 io_in_c_bypass_regNext_30_2_is_stationary_18;
  reg        [15:0]   io_in_c_bypass_regNext_30_3_data_18;
  reg                 io_in_c_bypass_regNext_30_3_is_stationary_18;
  reg        [15:0]   io_in_c_bypass_regNext_31_0_data_18;
  reg                 io_in_c_bypass_regNext_31_0_is_stationary_18;
  reg        [15:0]   io_in_c_bypass_regNext_31_1_data_18;
  reg                 io_in_c_bypass_regNext_31_1_is_stationary_18;
  reg        [15:0]   io_in_c_bypass_regNext_31_2_data_18;
  reg                 io_in_c_bypass_regNext_31_2_is_stationary_18;
  reg        [15:0]   io_in_c_bypass_regNext_31_3_data_18;
  reg                 io_in_c_bypass_regNext_31_3_is_stationary_18;
  reg        [15:0]   io_in_c_bypass_regNext_0_0_data_19;
  reg                 io_in_c_bypass_regNext_0_0_is_stationary_19;
  reg        [15:0]   io_in_c_bypass_regNext_0_1_data_19;
  reg                 io_in_c_bypass_regNext_0_1_is_stationary_19;
  reg        [15:0]   io_in_c_bypass_regNext_0_2_data_19;
  reg                 io_in_c_bypass_regNext_0_2_is_stationary_19;
  reg        [15:0]   io_in_c_bypass_regNext_0_3_data_19;
  reg                 io_in_c_bypass_regNext_0_3_is_stationary_19;
  reg        [15:0]   io_in_c_bypass_regNext_1_0_data_19;
  reg                 io_in_c_bypass_regNext_1_0_is_stationary_19;
  reg        [15:0]   io_in_c_bypass_regNext_1_1_data_19;
  reg                 io_in_c_bypass_regNext_1_1_is_stationary_19;
  reg        [15:0]   io_in_c_bypass_regNext_1_2_data_19;
  reg                 io_in_c_bypass_regNext_1_2_is_stationary_19;
  reg        [15:0]   io_in_c_bypass_regNext_1_3_data_19;
  reg                 io_in_c_bypass_regNext_1_3_is_stationary_19;
  reg        [15:0]   io_in_c_bypass_regNext_2_0_data_19;
  reg                 io_in_c_bypass_regNext_2_0_is_stationary_19;
  reg        [15:0]   io_in_c_bypass_regNext_2_1_data_19;
  reg                 io_in_c_bypass_regNext_2_1_is_stationary_19;
  reg        [15:0]   io_in_c_bypass_regNext_2_2_data_19;
  reg                 io_in_c_bypass_regNext_2_2_is_stationary_19;
  reg        [15:0]   io_in_c_bypass_regNext_2_3_data_19;
  reg                 io_in_c_bypass_regNext_2_3_is_stationary_19;
  reg        [15:0]   io_in_c_bypass_regNext_3_0_data_19;
  reg                 io_in_c_bypass_regNext_3_0_is_stationary_19;
  reg        [15:0]   io_in_c_bypass_regNext_3_1_data_19;
  reg                 io_in_c_bypass_regNext_3_1_is_stationary_19;
  reg        [15:0]   io_in_c_bypass_regNext_3_2_data_19;
  reg                 io_in_c_bypass_regNext_3_2_is_stationary_19;
  reg        [15:0]   io_in_c_bypass_regNext_3_3_data_19;
  reg                 io_in_c_bypass_regNext_3_3_is_stationary_19;
  reg        [15:0]   io_in_c_bypass_regNext_4_0_data_19;
  reg                 io_in_c_bypass_regNext_4_0_is_stationary_19;
  reg        [15:0]   io_in_c_bypass_regNext_4_1_data_19;
  reg                 io_in_c_bypass_regNext_4_1_is_stationary_19;
  reg        [15:0]   io_in_c_bypass_regNext_4_2_data_19;
  reg                 io_in_c_bypass_regNext_4_2_is_stationary_19;
  reg        [15:0]   io_in_c_bypass_regNext_4_3_data_19;
  reg                 io_in_c_bypass_regNext_4_3_is_stationary_19;
  reg        [15:0]   io_in_c_bypass_regNext_5_0_data_19;
  reg                 io_in_c_bypass_regNext_5_0_is_stationary_19;
  reg        [15:0]   io_in_c_bypass_regNext_5_1_data_19;
  reg                 io_in_c_bypass_regNext_5_1_is_stationary_19;
  reg        [15:0]   io_in_c_bypass_regNext_5_2_data_19;
  reg                 io_in_c_bypass_regNext_5_2_is_stationary_19;
  reg        [15:0]   io_in_c_bypass_regNext_5_3_data_19;
  reg                 io_in_c_bypass_regNext_5_3_is_stationary_19;
  reg        [15:0]   io_in_c_bypass_regNext_6_0_data_19;
  reg                 io_in_c_bypass_regNext_6_0_is_stationary_19;
  reg        [15:0]   io_in_c_bypass_regNext_6_1_data_19;
  reg                 io_in_c_bypass_regNext_6_1_is_stationary_19;
  reg        [15:0]   io_in_c_bypass_regNext_6_2_data_19;
  reg                 io_in_c_bypass_regNext_6_2_is_stationary_19;
  reg        [15:0]   io_in_c_bypass_regNext_6_3_data_19;
  reg                 io_in_c_bypass_regNext_6_3_is_stationary_19;
  reg        [15:0]   io_in_c_bypass_regNext_7_0_data_19;
  reg                 io_in_c_bypass_regNext_7_0_is_stationary_19;
  reg        [15:0]   io_in_c_bypass_regNext_7_1_data_19;
  reg                 io_in_c_bypass_regNext_7_1_is_stationary_19;
  reg        [15:0]   io_in_c_bypass_regNext_7_2_data_19;
  reg                 io_in_c_bypass_regNext_7_2_is_stationary_19;
  reg        [15:0]   io_in_c_bypass_regNext_7_3_data_19;
  reg                 io_in_c_bypass_regNext_7_3_is_stationary_19;
  reg        [15:0]   io_in_c_bypass_regNext_8_0_data_19;
  reg                 io_in_c_bypass_regNext_8_0_is_stationary_19;
  reg        [15:0]   io_in_c_bypass_regNext_8_1_data_19;
  reg                 io_in_c_bypass_regNext_8_1_is_stationary_19;
  reg        [15:0]   io_in_c_bypass_regNext_8_2_data_19;
  reg                 io_in_c_bypass_regNext_8_2_is_stationary_19;
  reg        [15:0]   io_in_c_bypass_regNext_8_3_data_19;
  reg                 io_in_c_bypass_regNext_8_3_is_stationary_19;
  reg        [15:0]   io_in_c_bypass_regNext_9_0_data_19;
  reg                 io_in_c_bypass_regNext_9_0_is_stationary_19;
  reg        [15:0]   io_in_c_bypass_regNext_9_1_data_19;
  reg                 io_in_c_bypass_regNext_9_1_is_stationary_19;
  reg        [15:0]   io_in_c_bypass_regNext_9_2_data_19;
  reg                 io_in_c_bypass_regNext_9_2_is_stationary_19;
  reg        [15:0]   io_in_c_bypass_regNext_9_3_data_19;
  reg                 io_in_c_bypass_regNext_9_3_is_stationary_19;
  reg        [15:0]   io_in_c_bypass_regNext_10_0_data_19;
  reg                 io_in_c_bypass_regNext_10_0_is_stationary_19;
  reg        [15:0]   io_in_c_bypass_regNext_10_1_data_19;
  reg                 io_in_c_bypass_regNext_10_1_is_stationary_19;
  reg        [15:0]   io_in_c_bypass_regNext_10_2_data_19;
  reg                 io_in_c_bypass_regNext_10_2_is_stationary_19;
  reg        [15:0]   io_in_c_bypass_regNext_10_3_data_19;
  reg                 io_in_c_bypass_regNext_10_3_is_stationary_19;
  reg        [15:0]   io_in_c_bypass_regNext_11_0_data_19;
  reg                 io_in_c_bypass_regNext_11_0_is_stationary_19;
  reg        [15:0]   io_in_c_bypass_regNext_11_1_data_19;
  reg                 io_in_c_bypass_regNext_11_1_is_stationary_19;
  reg        [15:0]   io_in_c_bypass_regNext_11_2_data_19;
  reg                 io_in_c_bypass_regNext_11_2_is_stationary_19;
  reg        [15:0]   io_in_c_bypass_regNext_11_3_data_19;
  reg                 io_in_c_bypass_regNext_11_3_is_stationary_19;
  reg        [15:0]   io_in_c_bypass_regNext_12_0_data_19;
  reg                 io_in_c_bypass_regNext_12_0_is_stationary_19;
  reg        [15:0]   io_in_c_bypass_regNext_12_1_data_19;
  reg                 io_in_c_bypass_regNext_12_1_is_stationary_19;
  reg        [15:0]   io_in_c_bypass_regNext_12_2_data_19;
  reg                 io_in_c_bypass_regNext_12_2_is_stationary_19;
  reg        [15:0]   io_in_c_bypass_regNext_12_3_data_19;
  reg                 io_in_c_bypass_regNext_12_3_is_stationary_19;
  reg        [15:0]   io_in_c_bypass_regNext_13_0_data_19;
  reg                 io_in_c_bypass_regNext_13_0_is_stationary_19;
  reg        [15:0]   io_in_c_bypass_regNext_13_1_data_19;
  reg                 io_in_c_bypass_regNext_13_1_is_stationary_19;
  reg        [15:0]   io_in_c_bypass_regNext_13_2_data_19;
  reg                 io_in_c_bypass_regNext_13_2_is_stationary_19;
  reg        [15:0]   io_in_c_bypass_regNext_13_3_data_19;
  reg                 io_in_c_bypass_regNext_13_3_is_stationary_19;
  reg        [15:0]   io_in_c_bypass_regNext_14_0_data_19;
  reg                 io_in_c_bypass_regNext_14_0_is_stationary_19;
  reg        [15:0]   io_in_c_bypass_regNext_14_1_data_19;
  reg                 io_in_c_bypass_regNext_14_1_is_stationary_19;
  reg        [15:0]   io_in_c_bypass_regNext_14_2_data_19;
  reg                 io_in_c_bypass_regNext_14_2_is_stationary_19;
  reg        [15:0]   io_in_c_bypass_regNext_14_3_data_19;
  reg                 io_in_c_bypass_regNext_14_3_is_stationary_19;
  reg        [15:0]   io_in_c_bypass_regNext_15_0_data_19;
  reg                 io_in_c_bypass_regNext_15_0_is_stationary_19;
  reg        [15:0]   io_in_c_bypass_regNext_15_1_data_19;
  reg                 io_in_c_bypass_regNext_15_1_is_stationary_19;
  reg        [15:0]   io_in_c_bypass_regNext_15_2_data_19;
  reg                 io_in_c_bypass_regNext_15_2_is_stationary_19;
  reg        [15:0]   io_in_c_bypass_regNext_15_3_data_19;
  reg                 io_in_c_bypass_regNext_15_3_is_stationary_19;
  reg        [15:0]   io_in_c_bypass_regNext_16_0_data_19;
  reg                 io_in_c_bypass_regNext_16_0_is_stationary_19;
  reg        [15:0]   io_in_c_bypass_regNext_16_1_data_19;
  reg                 io_in_c_bypass_regNext_16_1_is_stationary_19;
  reg        [15:0]   io_in_c_bypass_regNext_16_2_data_19;
  reg                 io_in_c_bypass_regNext_16_2_is_stationary_19;
  reg        [15:0]   io_in_c_bypass_regNext_16_3_data_19;
  reg                 io_in_c_bypass_regNext_16_3_is_stationary_19;
  reg        [15:0]   io_in_c_bypass_regNext_17_0_data_19;
  reg                 io_in_c_bypass_regNext_17_0_is_stationary_19;
  reg        [15:0]   io_in_c_bypass_regNext_17_1_data_19;
  reg                 io_in_c_bypass_regNext_17_1_is_stationary_19;
  reg        [15:0]   io_in_c_bypass_regNext_17_2_data_19;
  reg                 io_in_c_bypass_regNext_17_2_is_stationary_19;
  reg        [15:0]   io_in_c_bypass_regNext_17_3_data_19;
  reg                 io_in_c_bypass_regNext_17_3_is_stationary_19;
  reg        [15:0]   io_in_c_bypass_regNext_18_0_data_19;
  reg                 io_in_c_bypass_regNext_18_0_is_stationary_19;
  reg        [15:0]   io_in_c_bypass_regNext_18_1_data_19;
  reg                 io_in_c_bypass_regNext_18_1_is_stationary_19;
  reg        [15:0]   io_in_c_bypass_regNext_18_2_data_19;
  reg                 io_in_c_bypass_regNext_18_2_is_stationary_19;
  reg        [15:0]   io_in_c_bypass_regNext_18_3_data_19;
  reg                 io_in_c_bypass_regNext_18_3_is_stationary_19;
  reg        [15:0]   io_in_c_bypass_regNext_19_0_data_19;
  reg                 io_in_c_bypass_regNext_19_0_is_stationary_19;
  reg        [15:0]   io_in_c_bypass_regNext_19_1_data_19;
  reg                 io_in_c_bypass_regNext_19_1_is_stationary_19;
  reg        [15:0]   io_in_c_bypass_regNext_19_2_data_19;
  reg                 io_in_c_bypass_regNext_19_2_is_stationary_19;
  reg        [15:0]   io_in_c_bypass_regNext_19_3_data_19;
  reg                 io_in_c_bypass_regNext_19_3_is_stationary_19;
  reg        [15:0]   io_in_c_bypass_regNext_20_0_data_19;
  reg                 io_in_c_bypass_regNext_20_0_is_stationary_19;
  reg        [15:0]   io_in_c_bypass_regNext_20_1_data_19;
  reg                 io_in_c_bypass_regNext_20_1_is_stationary_19;
  reg        [15:0]   io_in_c_bypass_regNext_20_2_data_19;
  reg                 io_in_c_bypass_regNext_20_2_is_stationary_19;
  reg        [15:0]   io_in_c_bypass_regNext_20_3_data_19;
  reg                 io_in_c_bypass_regNext_20_3_is_stationary_19;
  reg        [15:0]   io_in_c_bypass_regNext_21_0_data_19;
  reg                 io_in_c_bypass_regNext_21_0_is_stationary_19;
  reg        [15:0]   io_in_c_bypass_regNext_21_1_data_19;
  reg                 io_in_c_bypass_regNext_21_1_is_stationary_19;
  reg        [15:0]   io_in_c_bypass_regNext_21_2_data_19;
  reg                 io_in_c_bypass_regNext_21_2_is_stationary_19;
  reg        [15:0]   io_in_c_bypass_regNext_21_3_data_19;
  reg                 io_in_c_bypass_regNext_21_3_is_stationary_19;
  reg        [15:0]   io_in_c_bypass_regNext_22_0_data_19;
  reg                 io_in_c_bypass_regNext_22_0_is_stationary_19;
  reg        [15:0]   io_in_c_bypass_regNext_22_1_data_19;
  reg                 io_in_c_bypass_regNext_22_1_is_stationary_19;
  reg        [15:0]   io_in_c_bypass_regNext_22_2_data_19;
  reg                 io_in_c_bypass_regNext_22_2_is_stationary_19;
  reg        [15:0]   io_in_c_bypass_regNext_22_3_data_19;
  reg                 io_in_c_bypass_regNext_22_3_is_stationary_19;
  reg        [15:0]   io_in_c_bypass_regNext_23_0_data_19;
  reg                 io_in_c_bypass_regNext_23_0_is_stationary_19;
  reg        [15:0]   io_in_c_bypass_regNext_23_1_data_19;
  reg                 io_in_c_bypass_regNext_23_1_is_stationary_19;
  reg        [15:0]   io_in_c_bypass_regNext_23_2_data_19;
  reg                 io_in_c_bypass_regNext_23_2_is_stationary_19;
  reg        [15:0]   io_in_c_bypass_regNext_23_3_data_19;
  reg                 io_in_c_bypass_regNext_23_3_is_stationary_19;
  reg        [15:0]   io_in_c_bypass_regNext_24_0_data_19;
  reg                 io_in_c_bypass_regNext_24_0_is_stationary_19;
  reg        [15:0]   io_in_c_bypass_regNext_24_1_data_19;
  reg                 io_in_c_bypass_regNext_24_1_is_stationary_19;
  reg        [15:0]   io_in_c_bypass_regNext_24_2_data_19;
  reg                 io_in_c_bypass_regNext_24_2_is_stationary_19;
  reg        [15:0]   io_in_c_bypass_regNext_24_3_data_19;
  reg                 io_in_c_bypass_regNext_24_3_is_stationary_19;
  reg        [15:0]   io_in_c_bypass_regNext_25_0_data_19;
  reg                 io_in_c_bypass_regNext_25_0_is_stationary_19;
  reg        [15:0]   io_in_c_bypass_regNext_25_1_data_19;
  reg                 io_in_c_bypass_regNext_25_1_is_stationary_19;
  reg        [15:0]   io_in_c_bypass_regNext_25_2_data_19;
  reg                 io_in_c_bypass_regNext_25_2_is_stationary_19;
  reg        [15:0]   io_in_c_bypass_regNext_25_3_data_19;
  reg                 io_in_c_bypass_regNext_25_3_is_stationary_19;
  reg        [15:0]   io_in_c_bypass_regNext_26_0_data_19;
  reg                 io_in_c_bypass_regNext_26_0_is_stationary_19;
  reg        [15:0]   io_in_c_bypass_regNext_26_1_data_19;
  reg                 io_in_c_bypass_regNext_26_1_is_stationary_19;
  reg        [15:0]   io_in_c_bypass_regNext_26_2_data_19;
  reg                 io_in_c_bypass_regNext_26_2_is_stationary_19;
  reg        [15:0]   io_in_c_bypass_regNext_26_3_data_19;
  reg                 io_in_c_bypass_regNext_26_3_is_stationary_19;
  reg        [15:0]   io_in_c_bypass_regNext_27_0_data_19;
  reg                 io_in_c_bypass_regNext_27_0_is_stationary_19;
  reg        [15:0]   io_in_c_bypass_regNext_27_1_data_19;
  reg                 io_in_c_bypass_regNext_27_1_is_stationary_19;
  reg        [15:0]   io_in_c_bypass_regNext_27_2_data_19;
  reg                 io_in_c_bypass_regNext_27_2_is_stationary_19;
  reg        [15:0]   io_in_c_bypass_regNext_27_3_data_19;
  reg                 io_in_c_bypass_regNext_27_3_is_stationary_19;
  reg        [15:0]   io_in_c_bypass_regNext_28_0_data_19;
  reg                 io_in_c_bypass_regNext_28_0_is_stationary_19;
  reg        [15:0]   io_in_c_bypass_regNext_28_1_data_19;
  reg                 io_in_c_bypass_regNext_28_1_is_stationary_19;
  reg        [15:0]   io_in_c_bypass_regNext_28_2_data_19;
  reg                 io_in_c_bypass_regNext_28_2_is_stationary_19;
  reg        [15:0]   io_in_c_bypass_regNext_28_3_data_19;
  reg                 io_in_c_bypass_regNext_28_3_is_stationary_19;
  reg        [15:0]   io_in_c_bypass_regNext_29_0_data_19;
  reg                 io_in_c_bypass_regNext_29_0_is_stationary_19;
  reg        [15:0]   io_in_c_bypass_regNext_29_1_data_19;
  reg                 io_in_c_bypass_regNext_29_1_is_stationary_19;
  reg        [15:0]   io_in_c_bypass_regNext_29_2_data_19;
  reg                 io_in_c_bypass_regNext_29_2_is_stationary_19;
  reg        [15:0]   io_in_c_bypass_regNext_29_3_data_19;
  reg                 io_in_c_bypass_regNext_29_3_is_stationary_19;
  reg        [15:0]   io_in_c_bypass_regNext_30_0_data_19;
  reg                 io_in_c_bypass_regNext_30_0_is_stationary_19;
  reg        [15:0]   io_in_c_bypass_regNext_30_1_data_19;
  reg                 io_in_c_bypass_regNext_30_1_is_stationary_19;
  reg        [15:0]   io_in_c_bypass_regNext_30_2_data_19;
  reg                 io_in_c_bypass_regNext_30_2_is_stationary_19;
  reg        [15:0]   io_in_c_bypass_regNext_30_3_data_19;
  reg                 io_in_c_bypass_regNext_30_3_is_stationary_19;
  reg        [15:0]   io_in_c_bypass_regNext_31_0_data_19;
  reg                 io_in_c_bypass_regNext_31_0_is_stationary_19;
  reg        [15:0]   io_in_c_bypass_regNext_31_1_data_19;
  reg                 io_in_c_bypass_regNext_31_1_is_stationary_19;
  reg        [15:0]   io_in_c_bypass_regNext_31_2_data_19;
  reg                 io_in_c_bypass_regNext_31_2_is_stationary_19;
  reg        [15:0]   io_in_c_bypass_regNext_31_3_data_19;
  reg                 io_in_c_bypass_regNext_31_3_is_stationary_19;
  reg        [15:0]   io_in_c_bypass_regNext_0_0_data_20;
  reg                 io_in_c_bypass_regNext_0_0_is_stationary_20;
  reg        [15:0]   io_in_c_bypass_regNext_0_1_data_20;
  reg                 io_in_c_bypass_regNext_0_1_is_stationary_20;
  reg        [15:0]   io_in_c_bypass_regNext_0_2_data_20;
  reg                 io_in_c_bypass_regNext_0_2_is_stationary_20;
  reg        [15:0]   io_in_c_bypass_regNext_0_3_data_20;
  reg                 io_in_c_bypass_regNext_0_3_is_stationary_20;
  reg        [15:0]   io_in_c_bypass_regNext_1_0_data_20;
  reg                 io_in_c_bypass_regNext_1_0_is_stationary_20;
  reg        [15:0]   io_in_c_bypass_regNext_1_1_data_20;
  reg                 io_in_c_bypass_regNext_1_1_is_stationary_20;
  reg        [15:0]   io_in_c_bypass_regNext_1_2_data_20;
  reg                 io_in_c_bypass_regNext_1_2_is_stationary_20;
  reg        [15:0]   io_in_c_bypass_regNext_1_3_data_20;
  reg                 io_in_c_bypass_regNext_1_3_is_stationary_20;
  reg        [15:0]   io_in_c_bypass_regNext_2_0_data_20;
  reg                 io_in_c_bypass_regNext_2_0_is_stationary_20;
  reg        [15:0]   io_in_c_bypass_regNext_2_1_data_20;
  reg                 io_in_c_bypass_regNext_2_1_is_stationary_20;
  reg        [15:0]   io_in_c_bypass_regNext_2_2_data_20;
  reg                 io_in_c_bypass_regNext_2_2_is_stationary_20;
  reg        [15:0]   io_in_c_bypass_regNext_2_3_data_20;
  reg                 io_in_c_bypass_regNext_2_3_is_stationary_20;
  reg        [15:0]   io_in_c_bypass_regNext_3_0_data_20;
  reg                 io_in_c_bypass_regNext_3_0_is_stationary_20;
  reg        [15:0]   io_in_c_bypass_regNext_3_1_data_20;
  reg                 io_in_c_bypass_regNext_3_1_is_stationary_20;
  reg        [15:0]   io_in_c_bypass_regNext_3_2_data_20;
  reg                 io_in_c_bypass_regNext_3_2_is_stationary_20;
  reg        [15:0]   io_in_c_bypass_regNext_3_3_data_20;
  reg                 io_in_c_bypass_regNext_3_3_is_stationary_20;
  reg        [15:0]   io_in_c_bypass_regNext_4_0_data_20;
  reg                 io_in_c_bypass_regNext_4_0_is_stationary_20;
  reg        [15:0]   io_in_c_bypass_regNext_4_1_data_20;
  reg                 io_in_c_bypass_regNext_4_1_is_stationary_20;
  reg        [15:0]   io_in_c_bypass_regNext_4_2_data_20;
  reg                 io_in_c_bypass_regNext_4_2_is_stationary_20;
  reg        [15:0]   io_in_c_bypass_regNext_4_3_data_20;
  reg                 io_in_c_bypass_regNext_4_3_is_stationary_20;
  reg        [15:0]   io_in_c_bypass_regNext_5_0_data_20;
  reg                 io_in_c_bypass_regNext_5_0_is_stationary_20;
  reg        [15:0]   io_in_c_bypass_regNext_5_1_data_20;
  reg                 io_in_c_bypass_regNext_5_1_is_stationary_20;
  reg        [15:0]   io_in_c_bypass_regNext_5_2_data_20;
  reg                 io_in_c_bypass_regNext_5_2_is_stationary_20;
  reg        [15:0]   io_in_c_bypass_regNext_5_3_data_20;
  reg                 io_in_c_bypass_regNext_5_3_is_stationary_20;
  reg        [15:0]   io_in_c_bypass_regNext_6_0_data_20;
  reg                 io_in_c_bypass_regNext_6_0_is_stationary_20;
  reg        [15:0]   io_in_c_bypass_regNext_6_1_data_20;
  reg                 io_in_c_bypass_regNext_6_1_is_stationary_20;
  reg        [15:0]   io_in_c_bypass_regNext_6_2_data_20;
  reg                 io_in_c_bypass_regNext_6_2_is_stationary_20;
  reg        [15:0]   io_in_c_bypass_regNext_6_3_data_20;
  reg                 io_in_c_bypass_regNext_6_3_is_stationary_20;
  reg        [15:0]   io_in_c_bypass_regNext_7_0_data_20;
  reg                 io_in_c_bypass_regNext_7_0_is_stationary_20;
  reg        [15:0]   io_in_c_bypass_regNext_7_1_data_20;
  reg                 io_in_c_bypass_regNext_7_1_is_stationary_20;
  reg        [15:0]   io_in_c_bypass_regNext_7_2_data_20;
  reg                 io_in_c_bypass_regNext_7_2_is_stationary_20;
  reg        [15:0]   io_in_c_bypass_regNext_7_3_data_20;
  reg                 io_in_c_bypass_regNext_7_3_is_stationary_20;
  reg        [15:0]   io_in_c_bypass_regNext_8_0_data_20;
  reg                 io_in_c_bypass_regNext_8_0_is_stationary_20;
  reg        [15:0]   io_in_c_bypass_regNext_8_1_data_20;
  reg                 io_in_c_bypass_regNext_8_1_is_stationary_20;
  reg        [15:0]   io_in_c_bypass_regNext_8_2_data_20;
  reg                 io_in_c_bypass_regNext_8_2_is_stationary_20;
  reg        [15:0]   io_in_c_bypass_regNext_8_3_data_20;
  reg                 io_in_c_bypass_regNext_8_3_is_stationary_20;
  reg        [15:0]   io_in_c_bypass_regNext_9_0_data_20;
  reg                 io_in_c_bypass_regNext_9_0_is_stationary_20;
  reg        [15:0]   io_in_c_bypass_regNext_9_1_data_20;
  reg                 io_in_c_bypass_regNext_9_1_is_stationary_20;
  reg        [15:0]   io_in_c_bypass_regNext_9_2_data_20;
  reg                 io_in_c_bypass_regNext_9_2_is_stationary_20;
  reg        [15:0]   io_in_c_bypass_regNext_9_3_data_20;
  reg                 io_in_c_bypass_regNext_9_3_is_stationary_20;
  reg        [15:0]   io_in_c_bypass_regNext_10_0_data_20;
  reg                 io_in_c_bypass_regNext_10_0_is_stationary_20;
  reg        [15:0]   io_in_c_bypass_regNext_10_1_data_20;
  reg                 io_in_c_bypass_regNext_10_1_is_stationary_20;
  reg        [15:0]   io_in_c_bypass_regNext_10_2_data_20;
  reg                 io_in_c_bypass_regNext_10_2_is_stationary_20;
  reg        [15:0]   io_in_c_bypass_regNext_10_3_data_20;
  reg                 io_in_c_bypass_regNext_10_3_is_stationary_20;
  reg        [15:0]   io_in_c_bypass_regNext_11_0_data_20;
  reg                 io_in_c_bypass_regNext_11_0_is_stationary_20;
  reg        [15:0]   io_in_c_bypass_regNext_11_1_data_20;
  reg                 io_in_c_bypass_regNext_11_1_is_stationary_20;
  reg        [15:0]   io_in_c_bypass_regNext_11_2_data_20;
  reg                 io_in_c_bypass_regNext_11_2_is_stationary_20;
  reg        [15:0]   io_in_c_bypass_regNext_11_3_data_20;
  reg                 io_in_c_bypass_regNext_11_3_is_stationary_20;
  reg        [15:0]   io_in_c_bypass_regNext_12_0_data_20;
  reg                 io_in_c_bypass_regNext_12_0_is_stationary_20;
  reg        [15:0]   io_in_c_bypass_regNext_12_1_data_20;
  reg                 io_in_c_bypass_regNext_12_1_is_stationary_20;
  reg        [15:0]   io_in_c_bypass_regNext_12_2_data_20;
  reg                 io_in_c_bypass_regNext_12_2_is_stationary_20;
  reg        [15:0]   io_in_c_bypass_regNext_12_3_data_20;
  reg                 io_in_c_bypass_regNext_12_3_is_stationary_20;
  reg        [15:0]   io_in_c_bypass_regNext_13_0_data_20;
  reg                 io_in_c_bypass_regNext_13_0_is_stationary_20;
  reg        [15:0]   io_in_c_bypass_regNext_13_1_data_20;
  reg                 io_in_c_bypass_regNext_13_1_is_stationary_20;
  reg        [15:0]   io_in_c_bypass_regNext_13_2_data_20;
  reg                 io_in_c_bypass_regNext_13_2_is_stationary_20;
  reg        [15:0]   io_in_c_bypass_regNext_13_3_data_20;
  reg                 io_in_c_bypass_regNext_13_3_is_stationary_20;
  reg        [15:0]   io_in_c_bypass_regNext_14_0_data_20;
  reg                 io_in_c_bypass_regNext_14_0_is_stationary_20;
  reg        [15:0]   io_in_c_bypass_regNext_14_1_data_20;
  reg                 io_in_c_bypass_regNext_14_1_is_stationary_20;
  reg        [15:0]   io_in_c_bypass_regNext_14_2_data_20;
  reg                 io_in_c_bypass_regNext_14_2_is_stationary_20;
  reg        [15:0]   io_in_c_bypass_regNext_14_3_data_20;
  reg                 io_in_c_bypass_regNext_14_3_is_stationary_20;
  reg        [15:0]   io_in_c_bypass_regNext_15_0_data_20;
  reg                 io_in_c_bypass_regNext_15_0_is_stationary_20;
  reg        [15:0]   io_in_c_bypass_regNext_15_1_data_20;
  reg                 io_in_c_bypass_regNext_15_1_is_stationary_20;
  reg        [15:0]   io_in_c_bypass_regNext_15_2_data_20;
  reg                 io_in_c_bypass_regNext_15_2_is_stationary_20;
  reg        [15:0]   io_in_c_bypass_regNext_15_3_data_20;
  reg                 io_in_c_bypass_regNext_15_3_is_stationary_20;
  reg        [15:0]   io_in_c_bypass_regNext_16_0_data_20;
  reg                 io_in_c_bypass_regNext_16_0_is_stationary_20;
  reg        [15:0]   io_in_c_bypass_regNext_16_1_data_20;
  reg                 io_in_c_bypass_regNext_16_1_is_stationary_20;
  reg        [15:0]   io_in_c_bypass_regNext_16_2_data_20;
  reg                 io_in_c_bypass_regNext_16_2_is_stationary_20;
  reg        [15:0]   io_in_c_bypass_regNext_16_3_data_20;
  reg                 io_in_c_bypass_regNext_16_3_is_stationary_20;
  reg        [15:0]   io_in_c_bypass_regNext_17_0_data_20;
  reg                 io_in_c_bypass_regNext_17_0_is_stationary_20;
  reg        [15:0]   io_in_c_bypass_regNext_17_1_data_20;
  reg                 io_in_c_bypass_regNext_17_1_is_stationary_20;
  reg        [15:0]   io_in_c_bypass_regNext_17_2_data_20;
  reg                 io_in_c_bypass_regNext_17_2_is_stationary_20;
  reg        [15:0]   io_in_c_bypass_regNext_17_3_data_20;
  reg                 io_in_c_bypass_regNext_17_3_is_stationary_20;
  reg        [15:0]   io_in_c_bypass_regNext_18_0_data_20;
  reg                 io_in_c_bypass_regNext_18_0_is_stationary_20;
  reg        [15:0]   io_in_c_bypass_regNext_18_1_data_20;
  reg                 io_in_c_bypass_regNext_18_1_is_stationary_20;
  reg        [15:0]   io_in_c_bypass_regNext_18_2_data_20;
  reg                 io_in_c_bypass_regNext_18_2_is_stationary_20;
  reg        [15:0]   io_in_c_bypass_regNext_18_3_data_20;
  reg                 io_in_c_bypass_regNext_18_3_is_stationary_20;
  reg        [15:0]   io_in_c_bypass_regNext_19_0_data_20;
  reg                 io_in_c_bypass_regNext_19_0_is_stationary_20;
  reg        [15:0]   io_in_c_bypass_regNext_19_1_data_20;
  reg                 io_in_c_bypass_regNext_19_1_is_stationary_20;
  reg        [15:0]   io_in_c_bypass_regNext_19_2_data_20;
  reg                 io_in_c_bypass_regNext_19_2_is_stationary_20;
  reg        [15:0]   io_in_c_bypass_regNext_19_3_data_20;
  reg                 io_in_c_bypass_regNext_19_3_is_stationary_20;
  reg        [15:0]   io_in_c_bypass_regNext_20_0_data_20;
  reg                 io_in_c_bypass_regNext_20_0_is_stationary_20;
  reg        [15:0]   io_in_c_bypass_regNext_20_1_data_20;
  reg                 io_in_c_bypass_regNext_20_1_is_stationary_20;
  reg        [15:0]   io_in_c_bypass_regNext_20_2_data_20;
  reg                 io_in_c_bypass_regNext_20_2_is_stationary_20;
  reg        [15:0]   io_in_c_bypass_regNext_20_3_data_20;
  reg                 io_in_c_bypass_regNext_20_3_is_stationary_20;
  reg        [15:0]   io_in_c_bypass_regNext_21_0_data_20;
  reg                 io_in_c_bypass_regNext_21_0_is_stationary_20;
  reg        [15:0]   io_in_c_bypass_regNext_21_1_data_20;
  reg                 io_in_c_bypass_regNext_21_1_is_stationary_20;
  reg        [15:0]   io_in_c_bypass_regNext_21_2_data_20;
  reg                 io_in_c_bypass_regNext_21_2_is_stationary_20;
  reg        [15:0]   io_in_c_bypass_regNext_21_3_data_20;
  reg                 io_in_c_bypass_regNext_21_3_is_stationary_20;
  reg        [15:0]   io_in_c_bypass_regNext_22_0_data_20;
  reg                 io_in_c_bypass_regNext_22_0_is_stationary_20;
  reg        [15:0]   io_in_c_bypass_regNext_22_1_data_20;
  reg                 io_in_c_bypass_regNext_22_1_is_stationary_20;
  reg        [15:0]   io_in_c_bypass_regNext_22_2_data_20;
  reg                 io_in_c_bypass_regNext_22_2_is_stationary_20;
  reg        [15:0]   io_in_c_bypass_regNext_22_3_data_20;
  reg                 io_in_c_bypass_regNext_22_3_is_stationary_20;
  reg        [15:0]   io_in_c_bypass_regNext_23_0_data_20;
  reg                 io_in_c_bypass_regNext_23_0_is_stationary_20;
  reg        [15:0]   io_in_c_bypass_regNext_23_1_data_20;
  reg                 io_in_c_bypass_regNext_23_1_is_stationary_20;
  reg        [15:0]   io_in_c_bypass_regNext_23_2_data_20;
  reg                 io_in_c_bypass_regNext_23_2_is_stationary_20;
  reg        [15:0]   io_in_c_bypass_regNext_23_3_data_20;
  reg                 io_in_c_bypass_regNext_23_3_is_stationary_20;
  reg        [15:0]   io_in_c_bypass_regNext_24_0_data_20;
  reg                 io_in_c_bypass_regNext_24_0_is_stationary_20;
  reg        [15:0]   io_in_c_bypass_regNext_24_1_data_20;
  reg                 io_in_c_bypass_regNext_24_1_is_stationary_20;
  reg        [15:0]   io_in_c_bypass_regNext_24_2_data_20;
  reg                 io_in_c_bypass_regNext_24_2_is_stationary_20;
  reg        [15:0]   io_in_c_bypass_regNext_24_3_data_20;
  reg                 io_in_c_bypass_regNext_24_3_is_stationary_20;
  reg        [15:0]   io_in_c_bypass_regNext_25_0_data_20;
  reg                 io_in_c_bypass_regNext_25_0_is_stationary_20;
  reg        [15:0]   io_in_c_bypass_regNext_25_1_data_20;
  reg                 io_in_c_bypass_regNext_25_1_is_stationary_20;
  reg        [15:0]   io_in_c_bypass_regNext_25_2_data_20;
  reg                 io_in_c_bypass_regNext_25_2_is_stationary_20;
  reg        [15:0]   io_in_c_bypass_regNext_25_3_data_20;
  reg                 io_in_c_bypass_regNext_25_3_is_stationary_20;
  reg        [15:0]   io_in_c_bypass_regNext_26_0_data_20;
  reg                 io_in_c_bypass_regNext_26_0_is_stationary_20;
  reg        [15:0]   io_in_c_bypass_regNext_26_1_data_20;
  reg                 io_in_c_bypass_regNext_26_1_is_stationary_20;
  reg        [15:0]   io_in_c_bypass_regNext_26_2_data_20;
  reg                 io_in_c_bypass_regNext_26_2_is_stationary_20;
  reg        [15:0]   io_in_c_bypass_regNext_26_3_data_20;
  reg                 io_in_c_bypass_regNext_26_3_is_stationary_20;
  reg        [15:0]   io_in_c_bypass_regNext_27_0_data_20;
  reg                 io_in_c_bypass_regNext_27_0_is_stationary_20;
  reg        [15:0]   io_in_c_bypass_regNext_27_1_data_20;
  reg                 io_in_c_bypass_regNext_27_1_is_stationary_20;
  reg        [15:0]   io_in_c_bypass_regNext_27_2_data_20;
  reg                 io_in_c_bypass_regNext_27_2_is_stationary_20;
  reg        [15:0]   io_in_c_bypass_regNext_27_3_data_20;
  reg                 io_in_c_bypass_regNext_27_3_is_stationary_20;
  reg        [15:0]   io_in_c_bypass_regNext_28_0_data_20;
  reg                 io_in_c_bypass_regNext_28_0_is_stationary_20;
  reg        [15:0]   io_in_c_bypass_regNext_28_1_data_20;
  reg                 io_in_c_bypass_regNext_28_1_is_stationary_20;
  reg        [15:0]   io_in_c_bypass_regNext_28_2_data_20;
  reg                 io_in_c_bypass_regNext_28_2_is_stationary_20;
  reg        [15:0]   io_in_c_bypass_regNext_28_3_data_20;
  reg                 io_in_c_bypass_regNext_28_3_is_stationary_20;
  reg        [15:0]   io_in_c_bypass_regNext_29_0_data_20;
  reg                 io_in_c_bypass_regNext_29_0_is_stationary_20;
  reg        [15:0]   io_in_c_bypass_regNext_29_1_data_20;
  reg                 io_in_c_bypass_regNext_29_1_is_stationary_20;
  reg        [15:0]   io_in_c_bypass_regNext_29_2_data_20;
  reg                 io_in_c_bypass_regNext_29_2_is_stationary_20;
  reg        [15:0]   io_in_c_bypass_regNext_29_3_data_20;
  reg                 io_in_c_bypass_regNext_29_3_is_stationary_20;
  reg        [15:0]   io_in_c_bypass_regNext_30_0_data_20;
  reg                 io_in_c_bypass_regNext_30_0_is_stationary_20;
  reg        [15:0]   io_in_c_bypass_regNext_30_1_data_20;
  reg                 io_in_c_bypass_regNext_30_1_is_stationary_20;
  reg        [15:0]   io_in_c_bypass_regNext_30_2_data_20;
  reg                 io_in_c_bypass_regNext_30_2_is_stationary_20;
  reg        [15:0]   io_in_c_bypass_regNext_30_3_data_20;
  reg                 io_in_c_bypass_regNext_30_3_is_stationary_20;
  reg        [15:0]   io_in_c_bypass_regNext_31_0_data_20;
  reg                 io_in_c_bypass_regNext_31_0_is_stationary_20;
  reg        [15:0]   io_in_c_bypass_regNext_31_1_data_20;
  reg                 io_in_c_bypass_regNext_31_1_is_stationary_20;
  reg        [15:0]   io_in_c_bypass_regNext_31_2_data_20;
  reg                 io_in_c_bypass_regNext_31_2_is_stationary_20;
  reg        [15:0]   io_in_c_bypass_regNext_31_3_data_20;
  reg                 io_in_c_bypass_regNext_31_3_is_stationary_20;
  reg        [15:0]   io_in_c_bypass_regNext_0_0_data_21;
  reg                 io_in_c_bypass_regNext_0_0_is_stationary_21;
  reg        [15:0]   io_in_c_bypass_regNext_0_1_data_21;
  reg                 io_in_c_bypass_regNext_0_1_is_stationary_21;
  reg        [15:0]   io_in_c_bypass_regNext_0_2_data_21;
  reg                 io_in_c_bypass_regNext_0_2_is_stationary_21;
  reg        [15:0]   io_in_c_bypass_regNext_0_3_data_21;
  reg                 io_in_c_bypass_regNext_0_3_is_stationary_21;
  reg        [15:0]   io_in_c_bypass_regNext_1_0_data_21;
  reg                 io_in_c_bypass_regNext_1_0_is_stationary_21;
  reg        [15:0]   io_in_c_bypass_regNext_1_1_data_21;
  reg                 io_in_c_bypass_regNext_1_1_is_stationary_21;
  reg        [15:0]   io_in_c_bypass_regNext_1_2_data_21;
  reg                 io_in_c_bypass_regNext_1_2_is_stationary_21;
  reg        [15:0]   io_in_c_bypass_regNext_1_3_data_21;
  reg                 io_in_c_bypass_regNext_1_3_is_stationary_21;
  reg        [15:0]   io_in_c_bypass_regNext_2_0_data_21;
  reg                 io_in_c_bypass_regNext_2_0_is_stationary_21;
  reg        [15:0]   io_in_c_bypass_regNext_2_1_data_21;
  reg                 io_in_c_bypass_regNext_2_1_is_stationary_21;
  reg        [15:0]   io_in_c_bypass_regNext_2_2_data_21;
  reg                 io_in_c_bypass_regNext_2_2_is_stationary_21;
  reg        [15:0]   io_in_c_bypass_regNext_2_3_data_21;
  reg                 io_in_c_bypass_regNext_2_3_is_stationary_21;
  reg        [15:0]   io_in_c_bypass_regNext_3_0_data_21;
  reg                 io_in_c_bypass_regNext_3_0_is_stationary_21;
  reg        [15:0]   io_in_c_bypass_regNext_3_1_data_21;
  reg                 io_in_c_bypass_regNext_3_1_is_stationary_21;
  reg        [15:0]   io_in_c_bypass_regNext_3_2_data_21;
  reg                 io_in_c_bypass_regNext_3_2_is_stationary_21;
  reg        [15:0]   io_in_c_bypass_regNext_3_3_data_21;
  reg                 io_in_c_bypass_regNext_3_3_is_stationary_21;
  reg        [15:0]   io_in_c_bypass_regNext_4_0_data_21;
  reg                 io_in_c_bypass_regNext_4_0_is_stationary_21;
  reg        [15:0]   io_in_c_bypass_regNext_4_1_data_21;
  reg                 io_in_c_bypass_regNext_4_1_is_stationary_21;
  reg        [15:0]   io_in_c_bypass_regNext_4_2_data_21;
  reg                 io_in_c_bypass_regNext_4_2_is_stationary_21;
  reg        [15:0]   io_in_c_bypass_regNext_4_3_data_21;
  reg                 io_in_c_bypass_regNext_4_3_is_stationary_21;
  reg        [15:0]   io_in_c_bypass_regNext_5_0_data_21;
  reg                 io_in_c_bypass_regNext_5_0_is_stationary_21;
  reg        [15:0]   io_in_c_bypass_regNext_5_1_data_21;
  reg                 io_in_c_bypass_regNext_5_1_is_stationary_21;
  reg        [15:0]   io_in_c_bypass_regNext_5_2_data_21;
  reg                 io_in_c_bypass_regNext_5_2_is_stationary_21;
  reg        [15:0]   io_in_c_bypass_regNext_5_3_data_21;
  reg                 io_in_c_bypass_regNext_5_3_is_stationary_21;
  reg        [15:0]   io_in_c_bypass_regNext_6_0_data_21;
  reg                 io_in_c_bypass_regNext_6_0_is_stationary_21;
  reg        [15:0]   io_in_c_bypass_regNext_6_1_data_21;
  reg                 io_in_c_bypass_regNext_6_1_is_stationary_21;
  reg        [15:0]   io_in_c_bypass_regNext_6_2_data_21;
  reg                 io_in_c_bypass_regNext_6_2_is_stationary_21;
  reg        [15:0]   io_in_c_bypass_regNext_6_3_data_21;
  reg                 io_in_c_bypass_regNext_6_3_is_stationary_21;
  reg        [15:0]   io_in_c_bypass_regNext_7_0_data_21;
  reg                 io_in_c_bypass_regNext_7_0_is_stationary_21;
  reg        [15:0]   io_in_c_bypass_regNext_7_1_data_21;
  reg                 io_in_c_bypass_regNext_7_1_is_stationary_21;
  reg        [15:0]   io_in_c_bypass_regNext_7_2_data_21;
  reg                 io_in_c_bypass_regNext_7_2_is_stationary_21;
  reg        [15:0]   io_in_c_bypass_regNext_7_3_data_21;
  reg                 io_in_c_bypass_regNext_7_3_is_stationary_21;
  reg        [15:0]   io_in_c_bypass_regNext_8_0_data_21;
  reg                 io_in_c_bypass_regNext_8_0_is_stationary_21;
  reg        [15:0]   io_in_c_bypass_regNext_8_1_data_21;
  reg                 io_in_c_bypass_regNext_8_1_is_stationary_21;
  reg        [15:0]   io_in_c_bypass_regNext_8_2_data_21;
  reg                 io_in_c_bypass_regNext_8_2_is_stationary_21;
  reg        [15:0]   io_in_c_bypass_regNext_8_3_data_21;
  reg                 io_in_c_bypass_regNext_8_3_is_stationary_21;
  reg        [15:0]   io_in_c_bypass_regNext_9_0_data_21;
  reg                 io_in_c_bypass_regNext_9_0_is_stationary_21;
  reg        [15:0]   io_in_c_bypass_regNext_9_1_data_21;
  reg                 io_in_c_bypass_regNext_9_1_is_stationary_21;
  reg        [15:0]   io_in_c_bypass_regNext_9_2_data_21;
  reg                 io_in_c_bypass_regNext_9_2_is_stationary_21;
  reg        [15:0]   io_in_c_bypass_regNext_9_3_data_21;
  reg                 io_in_c_bypass_regNext_9_3_is_stationary_21;
  reg        [15:0]   io_in_c_bypass_regNext_10_0_data_21;
  reg                 io_in_c_bypass_regNext_10_0_is_stationary_21;
  reg        [15:0]   io_in_c_bypass_regNext_10_1_data_21;
  reg                 io_in_c_bypass_regNext_10_1_is_stationary_21;
  reg        [15:0]   io_in_c_bypass_regNext_10_2_data_21;
  reg                 io_in_c_bypass_regNext_10_2_is_stationary_21;
  reg        [15:0]   io_in_c_bypass_regNext_10_3_data_21;
  reg                 io_in_c_bypass_regNext_10_3_is_stationary_21;
  reg        [15:0]   io_in_c_bypass_regNext_11_0_data_21;
  reg                 io_in_c_bypass_regNext_11_0_is_stationary_21;
  reg        [15:0]   io_in_c_bypass_regNext_11_1_data_21;
  reg                 io_in_c_bypass_regNext_11_1_is_stationary_21;
  reg        [15:0]   io_in_c_bypass_regNext_11_2_data_21;
  reg                 io_in_c_bypass_regNext_11_2_is_stationary_21;
  reg        [15:0]   io_in_c_bypass_regNext_11_3_data_21;
  reg                 io_in_c_bypass_regNext_11_3_is_stationary_21;
  reg        [15:0]   io_in_c_bypass_regNext_12_0_data_21;
  reg                 io_in_c_bypass_regNext_12_0_is_stationary_21;
  reg        [15:0]   io_in_c_bypass_regNext_12_1_data_21;
  reg                 io_in_c_bypass_regNext_12_1_is_stationary_21;
  reg        [15:0]   io_in_c_bypass_regNext_12_2_data_21;
  reg                 io_in_c_bypass_regNext_12_2_is_stationary_21;
  reg        [15:0]   io_in_c_bypass_regNext_12_3_data_21;
  reg                 io_in_c_bypass_regNext_12_3_is_stationary_21;
  reg        [15:0]   io_in_c_bypass_regNext_13_0_data_21;
  reg                 io_in_c_bypass_regNext_13_0_is_stationary_21;
  reg        [15:0]   io_in_c_bypass_regNext_13_1_data_21;
  reg                 io_in_c_bypass_regNext_13_1_is_stationary_21;
  reg        [15:0]   io_in_c_bypass_regNext_13_2_data_21;
  reg                 io_in_c_bypass_regNext_13_2_is_stationary_21;
  reg        [15:0]   io_in_c_bypass_regNext_13_3_data_21;
  reg                 io_in_c_bypass_regNext_13_3_is_stationary_21;
  reg        [15:0]   io_in_c_bypass_regNext_14_0_data_21;
  reg                 io_in_c_bypass_regNext_14_0_is_stationary_21;
  reg        [15:0]   io_in_c_bypass_regNext_14_1_data_21;
  reg                 io_in_c_bypass_regNext_14_1_is_stationary_21;
  reg        [15:0]   io_in_c_bypass_regNext_14_2_data_21;
  reg                 io_in_c_bypass_regNext_14_2_is_stationary_21;
  reg        [15:0]   io_in_c_bypass_regNext_14_3_data_21;
  reg                 io_in_c_bypass_regNext_14_3_is_stationary_21;
  reg        [15:0]   io_in_c_bypass_regNext_15_0_data_21;
  reg                 io_in_c_bypass_regNext_15_0_is_stationary_21;
  reg        [15:0]   io_in_c_bypass_regNext_15_1_data_21;
  reg                 io_in_c_bypass_regNext_15_1_is_stationary_21;
  reg        [15:0]   io_in_c_bypass_regNext_15_2_data_21;
  reg                 io_in_c_bypass_regNext_15_2_is_stationary_21;
  reg        [15:0]   io_in_c_bypass_regNext_15_3_data_21;
  reg                 io_in_c_bypass_regNext_15_3_is_stationary_21;
  reg        [15:0]   io_in_c_bypass_regNext_16_0_data_21;
  reg                 io_in_c_bypass_regNext_16_0_is_stationary_21;
  reg        [15:0]   io_in_c_bypass_regNext_16_1_data_21;
  reg                 io_in_c_bypass_regNext_16_1_is_stationary_21;
  reg        [15:0]   io_in_c_bypass_regNext_16_2_data_21;
  reg                 io_in_c_bypass_regNext_16_2_is_stationary_21;
  reg        [15:0]   io_in_c_bypass_regNext_16_3_data_21;
  reg                 io_in_c_bypass_regNext_16_3_is_stationary_21;
  reg        [15:0]   io_in_c_bypass_regNext_17_0_data_21;
  reg                 io_in_c_bypass_regNext_17_0_is_stationary_21;
  reg        [15:0]   io_in_c_bypass_regNext_17_1_data_21;
  reg                 io_in_c_bypass_regNext_17_1_is_stationary_21;
  reg        [15:0]   io_in_c_bypass_regNext_17_2_data_21;
  reg                 io_in_c_bypass_regNext_17_2_is_stationary_21;
  reg        [15:0]   io_in_c_bypass_regNext_17_3_data_21;
  reg                 io_in_c_bypass_regNext_17_3_is_stationary_21;
  reg        [15:0]   io_in_c_bypass_regNext_18_0_data_21;
  reg                 io_in_c_bypass_regNext_18_0_is_stationary_21;
  reg        [15:0]   io_in_c_bypass_regNext_18_1_data_21;
  reg                 io_in_c_bypass_regNext_18_1_is_stationary_21;
  reg        [15:0]   io_in_c_bypass_regNext_18_2_data_21;
  reg                 io_in_c_bypass_regNext_18_2_is_stationary_21;
  reg        [15:0]   io_in_c_bypass_regNext_18_3_data_21;
  reg                 io_in_c_bypass_regNext_18_3_is_stationary_21;
  reg        [15:0]   io_in_c_bypass_regNext_19_0_data_21;
  reg                 io_in_c_bypass_regNext_19_0_is_stationary_21;
  reg        [15:0]   io_in_c_bypass_regNext_19_1_data_21;
  reg                 io_in_c_bypass_regNext_19_1_is_stationary_21;
  reg        [15:0]   io_in_c_bypass_regNext_19_2_data_21;
  reg                 io_in_c_bypass_regNext_19_2_is_stationary_21;
  reg        [15:0]   io_in_c_bypass_regNext_19_3_data_21;
  reg                 io_in_c_bypass_regNext_19_3_is_stationary_21;
  reg        [15:0]   io_in_c_bypass_regNext_20_0_data_21;
  reg                 io_in_c_bypass_regNext_20_0_is_stationary_21;
  reg        [15:0]   io_in_c_bypass_regNext_20_1_data_21;
  reg                 io_in_c_bypass_regNext_20_1_is_stationary_21;
  reg        [15:0]   io_in_c_bypass_regNext_20_2_data_21;
  reg                 io_in_c_bypass_regNext_20_2_is_stationary_21;
  reg        [15:0]   io_in_c_bypass_regNext_20_3_data_21;
  reg                 io_in_c_bypass_regNext_20_3_is_stationary_21;
  reg        [15:0]   io_in_c_bypass_regNext_21_0_data_21;
  reg                 io_in_c_bypass_regNext_21_0_is_stationary_21;
  reg        [15:0]   io_in_c_bypass_regNext_21_1_data_21;
  reg                 io_in_c_bypass_regNext_21_1_is_stationary_21;
  reg        [15:0]   io_in_c_bypass_regNext_21_2_data_21;
  reg                 io_in_c_bypass_regNext_21_2_is_stationary_21;
  reg        [15:0]   io_in_c_bypass_regNext_21_3_data_21;
  reg                 io_in_c_bypass_regNext_21_3_is_stationary_21;
  reg        [15:0]   io_in_c_bypass_regNext_22_0_data_21;
  reg                 io_in_c_bypass_regNext_22_0_is_stationary_21;
  reg        [15:0]   io_in_c_bypass_regNext_22_1_data_21;
  reg                 io_in_c_bypass_regNext_22_1_is_stationary_21;
  reg        [15:0]   io_in_c_bypass_regNext_22_2_data_21;
  reg                 io_in_c_bypass_regNext_22_2_is_stationary_21;
  reg        [15:0]   io_in_c_bypass_regNext_22_3_data_21;
  reg                 io_in_c_bypass_regNext_22_3_is_stationary_21;
  reg        [15:0]   io_in_c_bypass_regNext_23_0_data_21;
  reg                 io_in_c_bypass_regNext_23_0_is_stationary_21;
  reg        [15:0]   io_in_c_bypass_regNext_23_1_data_21;
  reg                 io_in_c_bypass_regNext_23_1_is_stationary_21;
  reg        [15:0]   io_in_c_bypass_regNext_23_2_data_21;
  reg                 io_in_c_bypass_regNext_23_2_is_stationary_21;
  reg        [15:0]   io_in_c_bypass_regNext_23_3_data_21;
  reg                 io_in_c_bypass_regNext_23_3_is_stationary_21;
  reg        [15:0]   io_in_c_bypass_regNext_24_0_data_21;
  reg                 io_in_c_bypass_regNext_24_0_is_stationary_21;
  reg        [15:0]   io_in_c_bypass_regNext_24_1_data_21;
  reg                 io_in_c_bypass_regNext_24_1_is_stationary_21;
  reg        [15:0]   io_in_c_bypass_regNext_24_2_data_21;
  reg                 io_in_c_bypass_regNext_24_2_is_stationary_21;
  reg        [15:0]   io_in_c_bypass_regNext_24_3_data_21;
  reg                 io_in_c_bypass_regNext_24_3_is_stationary_21;
  reg        [15:0]   io_in_c_bypass_regNext_25_0_data_21;
  reg                 io_in_c_bypass_regNext_25_0_is_stationary_21;
  reg        [15:0]   io_in_c_bypass_regNext_25_1_data_21;
  reg                 io_in_c_bypass_regNext_25_1_is_stationary_21;
  reg        [15:0]   io_in_c_bypass_regNext_25_2_data_21;
  reg                 io_in_c_bypass_regNext_25_2_is_stationary_21;
  reg        [15:0]   io_in_c_bypass_regNext_25_3_data_21;
  reg                 io_in_c_bypass_regNext_25_3_is_stationary_21;
  reg        [15:0]   io_in_c_bypass_regNext_26_0_data_21;
  reg                 io_in_c_bypass_regNext_26_0_is_stationary_21;
  reg        [15:0]   io_in_c_bypass_regNext_26_1_data_21;
  reg                 io_in_c_bypass_regNext_26_1_is_stationary_21;
  reg        [15:0]   io_in_c_bypass_regNext_26_2_data_21;
  reg                 io_in_c_bypass_regNext_26_2_is_stationary_21;
  reg        [15:0]   io_in_c_bypass_regNext_26_3_data_21;
  reg                 io_in_c_bypass_regNext_26_3_is_stationary_21;
  reg        [15:0]   io_in_c_bypass_regNext_27_0_data_21;
  reg                 io_in_c_bypass_regNext_27_0_is_stationary_21;
  reg        [15:0]   io_in_c_bypass_regNext_27_1_data_21;
  reg                 io_in_c_bypass_regNext_27_1_is_stationary_21;
  reg        [15:0]   io_in_c_bypass_regNext_27_2_data_21;
  reg                 io_in_c_bypass_regNext_27_2_is_stationary_21;
  reg        [15:0]   io_in_c_bypass_regNext_27_3_data_21;
  reg                 io_in_c_bypass_regNext_27_3_is_stationary_21;
  reg        [15:0]   io_in_c_bypass_regNext_28_0_data_21;
  reg                 io_in_c_bypass_regNext_28_0_is_stationary_21;
  reg        [15:0]   io_in_c_bypass_regNext_28_1_data_21;
  reg                 io_in_c_bypass_regNext_28_1_is_stationary_21;
  reg        [15:0]   io_in_c_bypass_regNext_28_2_data_21;
  reg                 io_in_c_bypass_regNext_28_2_is_stationary_21;
  reg        [15:0]   io_in_c_bypass_regNext_28_3_data_21;
  reg                 io_in_c_bypass_regNext_28_3_is_stationary_21;
  reg        [15:0]   io_in_c_bypass_regNext_29_0_data_21;
  reg                 io_in_c_bypass_regNext_29_0_is_stationary_21;
  reg        [15:0]   io_in_c_bypass_regNext_29_1_data_21;
  reg                 io_in_c_bypass_regNext_29_1_is_stationary_21;
  reg        [15:0]   io_in_c_bypass_regNext_29_2_data_21;
  reg                 io_in_c_bypass_regNext_29_2_is_stationary_21;
  reg        [15:0]   io_in_c_bypass_regNext_29_3_data_21;
  reg                 io_in_c_bypass_regNext_29_3_is_stationary_21;
  reg        [15:0]   io_in_c_bypass_regNext_30_0_data_21;
  reg                 io_in_c_bypass_regNext_30_0_is_stationary_21;
  reg        [15:0]   io_in_c_bypass_regNext_30_1_data_21;
  reg                 io_in_c_bypass_regNext_30_1_is_stationary_21;
  reg        [15:0]   io_in_c_bypass_regNext_30_2_data_21;
  reg                 io_in_c_bypass_regNext_30_2_is_stationary_21;
  reg        [15:0]   io_in_c_bypass_regNext_30_3_data_21;
  reg                 io_in_c_bypass_regNext_30_3_is_stationary_21;
  reg        [15:0]   io_in_c_bypass_regNext_31_0_data_21;
  reg                 io_in_c_bypass_regNext_31_0_is_stationary_21;
  reg        [15:0]   io_in_c_bypass_regNext_31_1_data_21;
  reg                 io_in_c_bypass_regNext_31_1_is_stationary_21;
  reg        [15:0]   io_in_c_bypass_regNext_31_2_data_21;
  reg                 io_in_c_bypass_regNext_31_2_is_stationary_21;
  reg        [15:0]   io_in_c_bypass_regNext_31_3_data_21;
  reg                 io_in_c_bypass_regNext_31_3_is_stationary_21;
  reg        [15:0]   io_in_c_bypass_regNext_0_0_data_22;
  reg                 io_in_c_bypass_regNext_0_0_is_stationary_22;
  reg        [15:0]   io_in_c_bypass_regNext_0_1_data_22;
  reg                 io_in_c_bypass_regNext_0_1_is_stationary_22;
  reg        [15:0]   io_in_c_bypass_regNext_0_2_data_22;
  reg                 io_in_c_bypass_regNext_0_2_is_stationary_22;
  reg        [15:0]   io_in_c_bypass_regNext_0_3_data_22;
  reg                 io_in_c_bypass_regNext_0_3_is_stationary_22;
  reg        [15:0]   io_in_c_bypass_regNext_1_0_data_22;
  reg                 io_in_c_bypass_regNext_1_0_is_stationary_22;
  reg        [15:0]   io_in_c_bypass_regNext_1_1_data_22;
  reg                 io_in_c_bypass_regNext_1_1_is_stationary_22;
  reg        [15:0]   io_in_c_bypass_regNext_1_2_data_22;
  reg                 io_in_c_bypass_regNext_1_2_is_stationary_22;
  reg        [15:0]   io_in_c_bypass_regNext_1_3_data_22;
  reg                 io_in_c_bypass_regNext_1_3_is_stationary_22;
  reg        [15:0]   io_in_c_bypass_regNext_2_0_data_22;
  reg                 io_in_c_bypass_regNext_2_0_is_stationary_22;
  reg        [15:0]   io_in_c_bypass_regNext_2_1_data_22;
  reg                 io_in_c_bypass_regNext_2_1_is_stationary_22;
  reg        [15:0]   io_in_c_bypass_regNext_2_2_data_22;
  reg                 io_in_c_bypass_regNext_2_2_is_stationary_22;
  reg        [15:0]   io_in_c_bypass_regNext_2_3_data_22;
  reg                 io_in_c_bypass_regNext_2_3_is_stationary_22;
  reg        [15:0]   io_in_c_bypass_regNext_3_0_data_22;
  reg                 io_in_c_bypass_regNext_3_0_is_stationary_22;
  reg        [15:0]   io_in_c_bypass_regNext_3_1_data_22;
  reg                 io_in_c_bypass_regNext_3_1_is_stationary_22;
  reg        [15:0]   io_in_c_bypass_regNext_3_2_data_22;
  reg                 io_in_c_bypass_regNext_3_2_is_stationary_22;
  reg        [15:0]   io_in_c_bypass_regNext_3_3_data_22;
  reg                 io_in_c_bypass_regNext_3_3_is_stationary_22;
  reg        [15:0]   io_in_c_bypass_regNext_4_0_data_22;
  reg                 io_in_c_bypass_regNext_4_0_is_stationary_22;
  reg        [15:0]   io_in_c_bypass_regNext_4_1_data_22;
  reg                 io_in_c_bypass_regNext_4_1_is_stationary_22;
  reg        [15:0]   io_in_c_bypass_regNext_4_2_data_22;
  reg                 io_in_c_bypass_regNext_4_2_is_stationary_22;
  reg        [15:0]   io_in_c_bypass_regNext_4_3_data_22;
  reg                 io_in_c_bypass_regNext_4_3_is_stationary_22;
  reg        [15:0]   io_in_c_bypass_regNext_5_0_data_22;
  reg                 io_in_c_bypass_regNext_5_0_is_stationary_22;
  reg        [15:0]   io_in_c_bypass_regNext_5_1_data_22;
  reg                 io_in_c_bypass_regNext_5_1_is_stationary_22;
  reg        [15:0]   io_in_c_bypass_regNext_5_2_data_22;
  reg                 io_in_c_bypass_regNext_5_2_is_stationary_22;
  reg        [15:0]   io_in_c_bypass_regNext_5_3_data_22;
  reg                 io_in_c_bypass_regNext_5_3_is_stationary_22;
  reg        [15:0]   io_in_c_bypass_regNext_6_0_data_22;
  reg                 io_in_c_bypass_regNext_6_0_is_stationary_22;
  reg        [15:0]   io_in_c_bypass_regNext_6_1_data_22;
  reg                 io_in_c_bypass_regNext_6_1_is_stationary_22;
  reg        [15:0]   io_in_c_bypass_regNext_6_2_data_22;
  reg                 io_in_c_bypass_regNext_6_2_is_stationary_22;
  reg        [15:0]   io_in_c_bypass_regNext_6_3_data_22;
  reg                 io_in_c_bypass_regNext_6_3_is_stationary_22;
  reg        [15:0]   io_in_c_bypass_regNext_7_0_data_22;
  reg                 io_in_c_bypass_regNext_7_0_is_stationary_22;
  reg        [15:0]   io_in_c_bypass_regNext_7_1_data_22;
  reg                 io_in_c_bypass_regNext_7_1_is_stationary_22;
  reg        [15:0]   io_in_c_bypass_regNext_7_2_data_22;
  reg                 io_in_c_bypass_regNext_7_2_is_stationary_22;
  reg        [15:0]   io_in_c_bypass_regNext_7_3_data_22;
  reg                 io_in_c_bypass_regNext_7_3_is_stationary_22;
  reg        [15:0]   io_in_c_bypass_regNext_8_0_data_22;
  reg                 io_in_c_bypass_regNext_8_0_is_stationary_22;
  reg        [15:0]   io_in_c_bypass_regNext_8_1_data_22;
  reg                 io_in_c_bypass_regNext_8_1_is_stationary_22;
  reg        [15:0]   io_in_c_bypass_regNext_8_2_data_22;
  reg                 io_in_c_bypass_regNext_8_2_is_stationary_22;
  reg        [15:0]   io_in_c_bypass_regNext_8_3_data_22;
  reg                 io_in_c_bypass_regNext_8_3_is_stationary_22;
  reg        [15:0]   io_in_c_bypass_regNext_9_0_data_22;
  reg                 io_in_c_bypass_regNext_9_0_is_stationary_22;
  reg        [15:0]   io_in_c_bypass_regNext_9_1_data_22;
  reg                 io_in_c_bypass_regNext_9_1_is_stationary_22;
  reg        [15:0]   io_in_c_bypass_regNext_9_2_data_22;
  reg                 io_in_c_bypass_regNext_9_2_is_stationary_22;
  reg        [15:0]   io_in_c_bypass_regNext_9_3_data_22;
  reg                 io_in_c_bypass_regNext_9_3_is_stationary_22;
  reg        [15:0]   io_in_c_bypass_regNext_10_0_data_22;
  reg                 io_in_c_bypass_regNext_10_0_is_stationary_22;
  reg        [15:0]   io_in_c_bypass_regNext_10_1_data_22;
  reg                 io_in_c_bypass_regNext_10_1_is_stationary_22;
  reg        [15:0]   io_in_c_bypass_regNext_10_2_data_22;
  reg                 io_in_c_bypass_regNext_10_2_is_stationary_22;
  reg        [15:0]   io_in_c_bypass_regNext_10_3_data_22;
  reg                 io_in_c_bypass_regNext_10_3_is_stationary_22;
  reg        [15:0]   io_in_c_bypass_regNext_11_0_data_22;
  reg                 io_in_c_bypass_regNext_11_0_is_stationary_22;
  reg        [15:0]   io_in_c_bypass_regNext_11_1_data_22;
  reg                 io_in_c_bypass_regNext_11_1_is_stationary_22;
  reg        [15:0]   io_in_c_bypass_regNext_11_2_data_22;
  reg                 io_in_c_bypass_regNext_11_2_is_stationary_22;
  reg        [15:0]   io_in_c_bypass_regNext_11_3_data_22;
  reg                 io_in_c_bypass_regNext_11_3_is_stationary_22;
  reg        [15:0]   io_in_c_bypass_regNext_12_0_data_22;
  reg                 io_in_c_bypass_regNext_12_0_is_stationary_22;
  reg        [15:0]   io_in_c_bypass_regNext_12_1_data_22;
  reg                 io_in_c_bypass_regNext_12_1_is_stationary_22;
  reg        [15:0]   io_in_c_bypass_regNext_12_2_data_22;
  reg                 io_in_c_bypass_regNext_12_2_is_stationary_22;
  reg        [15:0]   io_in_c_bypass_regNext_12_3_data_22;
  reg                 io_in_c_bypass_regNext_12_3_is_stationary_22;
  reg        [15:0]   io_in_c_bypass_regNext_13_0_data_22;
  reg                 io_in_c_bypass_regNext_13_0_is_stationary_22;
  reg        [15:0]   io_in_c_bypass_regNext_13_1_data_22;
  reg                 io_in_c_bypass_regNext_13_1_is_stationary_22;
  reg        [15:0]   io_in_c_bypass_regNext_13_2_data_22;
  reg                 io_in_c_bypass_regNext_13_2_is_stationary_22;
  reg        [15:0]   io_in_c_bypass_regNext_13_3_data_22;
  reg                 io_in_c_bypass_regNext_13_3_is_stationary_22;
  reg        [15:0]   io_in_c_bypass_regNext_14_0_data_22;
  reg                 io_in_c_bypass_regNext_14_0_is_stationary_22;
  reg        [15:0]   io_in_c_bypass_regNext_14_1_data_22;
  reg                 io_in_c_bypass_regNext_14_1_is_stationary_22;
  reg        [15:0]   io_in_c_bypass_regNext_14_2_data_22;
  reg                 io_in_c_bypass_regNext_14_2_is_stationary_22;
  reg        [15:0]   io_in_c_bypass_regNext_14_3_data_22;
  reg                 io_in_c_bypass_regNext_14_3_is_stationary_22;
  reg        [15:0]   io_in_c_bypass_regNext_15_0_data_22;
  reg                 io_in_c_bypass_regNext_15_0_is_stationary_22;
  reg        [15:0]   io_in_c_bypass_regNext_15_1_data_22;
  reg                 io_in_c_bypass_regNext_15_1_is_stationary_22;
  reg        [15:0]   io_in_c_bypass_regNext_15_2_data_22;
  reg                 io_in_c_bypass_regNext_15_2_is_stationary_22;
  reg        [15:0]   io_in_c_bypass_regNext_15_3_data_22;
  reg                 io_in_c_bypass_regNext_15_3_is_stationary_22;
  reg        [15:0]   io_in_c_bypass_regNext_16_0_data_22;
  reg                 io_in_c_bypass_regNext_16_0_is_stationary_22;
  reg        [15:0]   io_in_c_bypass_regNext_16_1_data_22;
  reg                 io_in_c_bypass_regNext_16_1_is_stationary_22;
  reg        [15:0]   io_in_c_bypass_regNext_16_2_data_22;
  reg                 io_in_c_bypass_regNext_16_2_is_stationary_22;
  reg        [15:0]   io_in_c_bypass_regNext_16_3_data_22;
  reg                 io_in_c_bypass_regNext_16_3_is_stationary_22;
  reg        [15:0]   io_in_c_bypass_regNext_17_0_data_22;
  reg                 io_in_c_bypass_regNext_17_0_is_stationary_22;
  reg        [15:0]   io_in_c_bypass_regNext_17_1_data_22;
  reg                 io_in_c_bypass_regNext_17_1_is_stationary_22;
  reg        [15:0]   io_in_c_bypass_regNext_17_2_data_22;
  reg                 io_in_c_bypass_regNext_17_2_is_stationary_22;
  reg        [15:0]   io_in_c_bypass_regNext_17_3_data_22;
  reg                 io_in_c_bypass_regNext_17_3_is_stationary_22;
  reg        [15:0]   io_in_c_bypass_regNext_18_0_data_22;
  reg                 io_in_c_bypass_regNext_18_0_is_stationary_22;
  reg        [15:0]   io_in_c_bypass_regNext_18_1_data_22;
  reg                 io_in_c_bypass_regNext_18_1_is_stationary_22;
  reg        [15:0]   io_in_c_bypass_regNext_18_2_data_22;
  reg                 io_in_c_bypass_regNext_18_2_is_stationary_22;
  reg        [15:0]   io_in_c_bypass_regNext_18_3_data_22;
  reg                 io_in_c_bypass_regNext_18_3_is_stationary_22;
  reg        [15:0]   io_in_c_bypass_regNext_19_0_data_22;
  reg                 io_in_c_bypass_regNext_19_0_is_stationary_22;
  reg        [15:0]   io_in_c_bypass_regNext_19_1_data_22;
  reg                 io_in_c_bypass_regNext_19_1_is_stationary_22;
  reg        [15:0]   io_in_c_bypass_regNext_19_2_data_22;
  reg                 io_in_c_bypass_regNext_19_2_is_stationary_22;
  reg        [15:0]   io_in_c_bypass_regNext_19_3_data_22;
  reg                 io_in_c_bypass_regNext_19_3_is_stationary_22;
  reg        [15:0]   io_in_c_bypass_regNext_20_0_data_22;
  reg                 io_in_c_bypass_regNext_20_0_is_stationary_22;
  reg        [15:0]   io_in_c_bypass_regNext_20_1_data_22;
  reg                 io_in_c_bypass_regNext_20_1_is_stationary_22;
  reg        [15:0]   io_in_c_bypass_regNext_20_2_data_22;
  reg                 io_in_c_bypass_regNext_20_2_is_stationary_22;
  reg        [15:0]   io_in_c_bypass_regNext_20_3_data_22;
  reg                 io_in_c_bypass_regNext_20_3_is_stationary_22;
  reg        [15:0]   io_in_c_bypass_regNext_21_0_data_22;
  reg                 io_in_c_bypass_regNext_21_0_is_stationary_22;
  reg        [15:0]   io_in_c_bypass_regNext_21_1_data_22;
  reg                 io_in_c_bypass_regNext_21_1_is_stationary_22;
  reg        [15:0]   io_in_c_bypass_regNext_21_2_data_22;
  reg                 io_in_c_bypass_regNext_21_2_is_stationary_22;
  reg        [15:0]   io_in_c_bypass_regNext_21_3_data_22;
  reg                 io_in_c_bypass_regNext_21_3_is_stationary_22;
  reg        [15:0]   io_in_c_bypass_regNext_22_0_data_22;
  reg                 io_in_c_bypass_regNext_22_0_is_stationary_22;
  reg        [15:0]   io_in_c_bypass_regNext_22_1_data_22;
  reg                 io_in_c_bypass_regNext_22_1_is_stationary_22;
  reg        [15:0]   io_in_c_bypass_regNext_22_2_data_22;
  reg                 io_in_c_bypass_regNext_22_2_is_stationary_22;
  reg        [15:0]   io_in_c_bypass_regNext_22_3_data_22;
  reg                 io_in_c_bypass_regNext_22_3_is_stationary_22;
  reg        [15:0]   io_in_c_bypass_regNext_23_0_data_22;
  reg                 io_in_c_bypass_regNext_23_0_is_stationary_22;
  reg        [15:0]   io_in_c_bypass_regNext_23_1_data_22;
  reg                 io_in_c_bypass_regNext_23_1_is_stationary_22;
  reg        [15:0]   io_in_c_bypass_regNext_23_2_data_22;
  reg                 io_in_c_bypass_regNext_23_2_is_stationary_22;
  reg        [15:0]   io_in_c_bypass_regNext_23_3_data_22;
  reg                 io_in_c_bypass_regNext_23_3_is_stationary_22;
  reg        [15:0]   io_in_c_bypass_regNext_24_0_data_22;
  reg                 io_in_c_bypass_regNext_24_0_is_stationary_22;
  reg        [15:0]   io_in_c_bypass_regNext_24_1_data_22;
  reg                 io_in_c_bypass_regNext_24_1_is_stationary_22;
  reg        [15:0]   io_in_c_bypass_regNext_24_2_data_22;
  reg                 io_in_c_bypass_regNext_24_2_is_stationary_22;
  reg        [15:0]   io_in_c_bypass_regNext_24_3_data_22;
  reg                 io_in_c_bypass_regNext_24_3_is_stationary_22;
  reg        [15:0]   io_in_c_bypass_regNext_25_0_data_22;
  reg                 io_in_c_bypass_regNext_25_0_is_stationary_22;
  reg        [15:0]   io_in_c_bypass_regNext_25_1_data_22;
  reg                 io_in_c_bypass_regNext_25_1_is_stationary_22;
  reg        [15:0]   io_in_c_bypass_regNext_25_2_data_22;
  reg                 io_in_c_bypass_regNext_25_2_is_stationary_22;
  reg        [15:0]   io_in_c_bypass_regNext_25_3_data_22;
  reg                 io_in_c_bypass_regNext_25_3_is_stationary_22;
  reg        [15:0]   io_in_c_bypass_regNext_26_0_data_22;
  reg                 io_in_c_bypass_regNext_26_0_is_stationary_22;
  reg        [15:0]   io_in_c_bypass_regNext_26_1_data_22;
  reg                 io_in_c_bypass_regNext_26_1_is_stationary_22;
  reg        [15:0]   io_in_c_bypass_regNext_26_2_data_22;
  reg                 io_in_c_bypass_regNext_26_2_is_stationary_22;
  reg        [15:0]   io_in_c_bypass_regNext_26_3_data_22;
  reg                 io_in_c_bypass_regNext_26_3_is_stationary_22;
  reg        [15:0]   io_in_c_bypass_regNext_27_0_data_22;
  reg                 io_in_c_bypass_regNext_27_0_is_stationary_22;
  reg        [15:0]   io_in_c_bypass_regNext_27_1_data_22;
  reg                 io_in_c_bypass_regNext_27_1_is_stationary_22;
  reg        [15:0]   io_in_c_bypass_regNext_27_2_data_22;
  reg                 io_in_c_bypass_regNext_27_2_is_stationary_22;
  reg        [15:0]   io_in_c_bypass_regNext_27_3_data_22;
  reg                 io_in_c_bypass_regNext_27_3_is_stationary_22;
  reg        [15:0]   io_in_c_bypass_regNext_28_0_data_22;
  reg                 io_in_c_bypass_regNext_28_0_is_stationary_22;
  reg        [15:0]   io_in_c_bypass_regNext_28_1_data_22;
  reg                 io_in_c_bypass_regNext_28_1_is_stationary_22;
  reg        [15:0]   io_in_c_bypass_regNext_28_2_data_22;
  reg                 io_in_c_bypass_regNext_28_2_is_stationary_22;
  reg        [15:0]   io_in_c_bypass_regNext_28_3_data_22;
  reg                 io_in_c_bypass_regNext_28_3_is_stationary_22;
  reg        [15:0]   io_in_c_bypass_regNext_29_0_data_22;
  reg                 io_in_c_bypass_regNext_29_0_is_stationary_22;
  reg        [15:0]   io_in_c_bypass_regNext_29_1_data_22;
  reg                 io_in_c_bypass_regNext_29_1_is_stationary_22;
  reg        [15:0]   io_in_c_bypass_regNext_29_2_data_22;
  reg                 io_in_c_bypass_regNext_29_2_is_stationary_22;
  reg        [15:0]   io_in_c_bypass_regNext_29_3_data_22;
  reg                 io_in_c_bypass_regNext_29_3_is_stationary_22;
  reg        [15:0]   io_in_c_bypass_regNext_30_0_data_22;
  reg                 io_in_c_bypass_regNext_30_0_is_stationary_22;
  reg        [15:0]   io_in_c_bypass_regNext_30_1_data_22;
  reg                 io_in_c_bypass_regNext_30_1_is_stationary_22;
  reg        [15:0]   io_in_c_bypass_regNext_30_2_data_22;
  reg                 io_in_c_bypass_regNext_30_2_is_stationary_22;
  reg        [15:0]   io_in_c_bypass_regNext_30_3_data_22;
  reg                 io_in_c_bypass_regNext_30_3_is_stationary_22;
  reg        [15:0]   io_in_c_bypass_regNext_31_0_data_22;
  reg                 io_in_c_bypass_regNext_31_0_is_stationary_22;
  reg        [15:0]   io_in_c_bypass_regNext_31_1_data_22;
  reg                 io_in_c_bypass_regNext_31_1_is_stationary_22;
  reg        [15:0]   io_in_c_bypass_regNext_31_2_data_22;
  reg                 io_in_c_bypass_regNext_31_2_is_stationary_22;
  reg        [15:0]   io_in_c_bypass_regNext_31_3_data_22;
  reg                 io_in_c_bypass_regNext_31_3_is_stationary_22;
  reg        [15:0]   io_in_c_bypass_regNext_0_0_data_23;
  reg                 io_in_c_bypass_regNext_0_0_is_stationary_23;
  reg        [15:0]   io_in_c_bypass_regNext_0_1_data_23;
  reg                 io_in_c_bypass_regNext_0_1_is_stationary_23;
  reg        [15:0]   io_in_c_bypass_regNext_0_2_data_23;
  reg                 io_in_c_bypass_regNext_0_2_is_stationary_23;
  reg        [15:0]   io_in_c_bypass_regNext_0_3_data_23;
  reg                 io_in_c_bypass_regNext_0_3_is_stationary_23;
  reg        [15:0]   io_in_c_bypass_regNext_1_0_data_23;
  reg                 io_in_c_bypass_regNext_1_0_is_stationary_23;
  reg        [15:0]   io_in_c_bypass_regNext_1_1_data_23;
  reg                 io_in_c_bypass_regNext_1_1_is_stationary_23;
  reg        [15:0]   io_in_c_bypass_regNext_1_2_data_23;
  reg                 io_in_c_bypass_regNext_1_2_is_stationary_23;
  reg        [15:0]   io_in_c_bypass_regNext_1_3_data_23;
  reg                 io_in_c_bypass_regNext_1_3_is_stationary_23;
  reg        [15:0]   io_in_c_bypass_regNext_2_0_data_23;
  reg                 io_in_c_bypass_regNext_2_0_is_stationary_23;
  reg        [15:0]   io_in_c_bypass_regNext_2_1_data_23;
  reg                 io_in_c_bypass_regNext_2_1_is_stationary_23;
  reg        [15:0]   io_in_c_bypass_regNext_2_2_data_23;
  reg                 io_in_c_bypass_regNext_2_2_is_stationary_23;
  reg        [15:0]   io_in_c_bypass_regNext_2_3_data_23;
  reg                 io_in_c_bypass_regNext_2_3_is_stationary_23;
  reg        [15:0]   io_in_c_bypass_regNext_3_0_data_23;
  reg                 io_in_c_bypass_regNext_3_0_is_stationary_23;
  reg        [15:0]   io_in_c_bypass_regNext_3_1_data_23;
  reg                 io_in_c_bypass_regNext_3_1_is_stationary_23;
  reg        [15:0]   io_in_c_bypass_regNext_3_2_data_23;
  reg                 io_in_c_bypass_regNext_3_2_is_stationary_23;
  reg        [15:0]   io_in_c_bypass_regNext_3_3_data_23;
  reg                 io_in_c_bypass_regNext_3_3_is_stationary_23;
  reg        [15:0]   io_in_c_bypass_regNext_4_0_data_23;
  reg                 io_in_c_bypass_regNext_4_0_is_stationary_23;
  reg        [15:0]   io_in_c_bypass_regNext_4_1_data_23;
  reg                 io_in_c_bypass_regNext_4_1_is_stationary_23;
  reg        [15:0]   io_in_c_bypass_regNext_4_2_data_23;
  reg                 io_in_c_bypass_regNext_4_2_is_stationary_23;
  reg        [15:0]   io_in_c_bypass_regNext_4_3_data_23;
  reg                 io_in_c_bypass_regNext_4_3_is_stationary_23;
  reg        [15:0]   io_in_c_bypass_regNext_5_0_data_23;
  reg                 io_in_c_bypass_regNext_5_0_is_stationary_23;
  reg        [15:0]   io_in_c_bypass_regNext_5_1_data_23;
  reg                 io_in_c_bypass_regNext_5_1_is_stationary_23;
  reg        [15:0]   io_in_c_bypass_regNext_5_2_data_23;
  reg                 io_in_c_bypass_regNext_5_2_is_stationary_23;
  reg        [15:0]   io_in_c_bypass_regNext_5_3_data_23;
  reg                 io_in_c_bypass_regNext_5_3_is_stationary_23;
  reg        [15:0]   io_in_c_bypass_regNext_6_0_data_23;
  reg                 io_in_c_bypass_regNext_6_0_is_stationary_23;
  reg        [15:0]   io_in_c_bypass_regNext_6_1_data_23;
  reg                 io_in_c_bypass_regNext_6_1_is_stationary_23;
  reg        [15:0]   io_in_c_bypass_regNext_6_2_data_23;
  reg                 io_in_c_bypass_regNext_6_2_is_stationary_23;
  reg        [15:0]   io_in_c_bypass_regNext_6_3_data_23;
  reg                 io_in_c_bypass_regNext_6_3_is_stationary_23;
  reg        [15:0]   io_in_c_bypass_regNext_7_0_data_23;
  reg                 io_in_c_bypass_regNext_7_0_is_stationary_23;
  reg        [15:0]   io_in_c_bypass_regNext_7_1_data_23;
  reg                 io_in_c_bypass_regNext_7_1_is_stationary_23;
  reg        [15:0]   io_in_c_bypass_regNext_7_2_data_23;
  reg                 io_in_c_bypass_regNext_7_2_is_stationary_23;
  reg        [15:0]   io_in_c_bypass_regNext_7_3_data_23;
  reg                 io_in_c_bypass_regNext_7_3_is_stationary_23;
  reg        [15:0]   io_in_c_bypass_regNext_8_0_data_23;
  reg                 io_in_c_bypass_regNext_8_0_is_stationary_23;
  reg        [15:0]   io_in_c_bypass_regNext_8_1_data_23;
  reg                 io_in_c_bypass_regNext_8_1_is_stationary_23;
  reg        [15:0]   io_in_c_bypass_regNext_8_2_data_23;
  reg                 io_in_c_bypass_regNext_8_2_is_stationary_23;
  reg        [15:0]   io_in_c_bypass_regNext_8_3_data_23;
  reg                 io_in_c_bypass_regNext_8_3_is_stationary_23;
  reg        [15:0]   io_in_c_bypass_regNext_9_0_data_23;
  reg                 io_in_c_bypass_regNext_9_0_is_stationary_23;
  reg        [15:0]   io_in_c_bypass_regNext_9_1_data_23;
  reg                 io_in_c_bypass_regNext_9_1_is_stationary_23;
  reg        [15:0]   io_in_c_bypass_regNext_9_2_data_23;
  reg                 io_in_c_bypass_regNext_9_2_is_stationary_23;
  reg        [15:0]   io_in_c_bypass_regNext_9_3_data_23;
  reg                 io_in_c_bypass_regNext_9_3_is_stationary_23;
  reg        [15:0]   io_in_c_bypass_regNext_10_0_data_23;
  reg                 io_in_c_bypass_regNext_10_0_is_stationary_23;
  reg        [15:0]   io_in_c_bypass_regNext_10_1_data_23;
  reg                 io_in_c_bypass_regNext_10_1_is_stationary_23;
  reg        [15:0]   io_in_c_bypass_regNext_10_2_data_23;
  reg                 io_in_c_bypass_regNext_10_2_is_stationary_23;
  reg        [15:0]   io_in_c_bypass_regNext_10_3_data_23;
  reg                 io_in_c_bypass_regNext_10_3_is_stationary_23;
  reg        [15:0]   io_in_c_bypass_regNext_11_0_data_23;
  reg                 io_in_c_bypass_regNext_11_0_is_stationary_23;
  reg        [15:0]   io_in_c_bypass_regNext_11_1_data_23;
  reg                 io_in_c_bypass_regNext_11_1_is_stationary_23;
  reg        [15:0]   io_in_c_bypass_regNext_11_2_data_23;
  reg                 io_in_c_bypass_regNext_11_2_is_stationary_23;
  reg        [15:0]   io_in_c_bypass_regNext_11_3_data_23;
  reg                 io_in_c_bypass_regNext_11_3_is_stationary_23;
  reg        [15:0]   io_in_c_bypass_regNext_12_0_data_23;
  reg                 io_in_c_bypass_regNext_12_0_is_stationary_23;
  reg        [15:0]   io_in_c_bypass_regNext_12_1_data_23;
  reg                 io_in_c_bypass_regNext_12_1_is_stationary_23;
  reg        [15:0]   io_in_c_bypass_regNext_12_2_data_23;
  reg                 io_in_c_bypass_regNext_12_2_is_stationary_23;
  reg        [15:0]   io_in_c_bypass_regNext_12_3_data_23;
  reg                 io_in_c_bypass_regNext_12_3_is_stationary_23;
  reg        [15:0]   io_in_c_bypass_regNext_13_0_data_23;
  reg                 io_in_c_bypass_regNext_13_0_is_stationary_23;
  reg        [15:0]   io_in_c_bypass_regNext_13_1_data_23;
  reg                 io_in_c_bypass_regNext_13_1_is_stationary_23;
  reg        [15:0]   io_in_c_bypass_regNext_13_2_data_23;
  reg                 io_in_c_bypass_regNext_13_2_is_stationary_23;
  reg        [15:0]   io_in_c_bypass_regNext_13_3_data_23;
  reg                 io_in_c_bypass_regNext_13_3_is_stationary_23;
  reg        [15:0]   io_in_c_bypass_regNext_14_0_data_23;
  reg                 io_in_c_bypass_regNext_14_0_is_stationary_23;
  reg        [15:0]   io_in_c_bypass_regNext_14_1_data_23;
  reg                 io_in_c_bypass_regNext_14_1_is_stationary_23;
  reg        [15:0]   io_in_c_bypass_regNext_14_2_data_23;
  reg                 io_in_c_bypass_regNext_14_2_is_stationary_23;
  reg        [15:0]   io_in_c_bypass_regNext_14_3_data_23;
  reg                 io_in_c_bypass_regNext_14_3_is_stationary_23;
  reg        [15:0]   io_in_c_bypass_regNext_15_0_data_23;
  reg                 io_in_c_bypass_regNext_15_0_is_stationary_23;
  reg        [15:0]   io_in_c_bypass_regNext_15_1_data_23;
  reg                 io_in_c_bypass_regNext_15_1_is_stationary_23;
  reg        [15:0]   io_in_c_bypass_regNext_15_2_data_23;
  reg                 io_in_c_bypass_regNext_15_2_is_stationary_23;
  reg        [15:0]   io_in_c_bypass_regNext_15_3_data_23;
  reg                 io_in_c_bypass_regNext_15_3_is_stationary_23;
  reg        [15:0]   io_in_c_bypass_regNext_16_0_data_23;
  reg                 io_in_c_bypass_regNext_16_0_is_stationary_23;
  reg        [15:0]   io_in_c_bypass_regNext_16_1_data_23;
  reg                 io_in_c_bypass_regNext_16_1_is_stationary_23;
  reg        [15:0]   io_in_c_bypass_regNext_16_2_data_23;
  reg                 io_in_c_bypass_regNext_16_2_is_stationary_23;
  reg        [15:0]   io_in_c_bypass_regNext_16_3_data_23;
  reg                 io_in_c_bypass_regNext_16_3_is_stationary_23;
  reg        [15:0]   io_in_c_bypass_regNext_17_0_data_23;
  reg                 io_in_c_bypass_regNext_17_0_is_stationary_23;
  reg        [15:0]   io_in_c_bypass_regNext_17_1_data_23;
  reg                 io_in_c_bypass_regNext_17_1_is_stationary_23;
  reg        [15:0]   io_in_c_bypass_regNext_17_2_data_23;
  reg                 io_in_c_bypass_regNext_17_2_is_stationary_23;
  reg        [15:0]   io_in_c_bypass_regNext_17_3_data_23;
  reg                 io_in_c_bypass_regNext_17_3_is_stationary_23;
  reg        [15:0]   io_in_c_bypass_regNext_18_0_data_23;
  reg                 io_in_c_bypass_regNext_18_0_is_stationary_23;
  reg        [15:0]   io_in_c_bypass_regNext_18_1_data_23;
  reg                 io_in_c_bypass_regNext_18_1_is_stationary_23;
  reg        [15:0]   io_in_c_bypass_regNext_18_2_data_23;
  reg                 io_in_c_bypass_regNext_18_2_is_stationary_23;
  reg        [15:0]   io_in_c_bypass_regNext_18_3_data_23;
  reg                 io_in_c_bypass_regNext_18_3_is_stationary_23;
  reg        [15:0]   io_in_c_bypass_regNext_19_0_data_23;
  reg                 io_in_c_bypass_regNext_19_0_is_stationary_23;
  reg        [15:0]   io_in_c_bypass_regNext_19_1_data_23;
  reg                 io_in_c_bypass_regNext_19_1_is_stationary_23;
  reg        [15:0]   io_in_c_bypass_regNext_19_2_data_23;
  reg                 io_in_c_bypass_regNext_19_2_is_stationary_23;
  reg        [15:0]   io_in_c_bypass_regNext_19_3_data_23;
  reg                 io_in_c_bypass_regNext_19_3_is_stationary_23;
  reg        [15:0]   io_in_c_bypass_regNext_20_0_data_23;
  reg                 io_in_c_bypass_regNext_20_0_is_stationary_23;
  reg        [15:0]   io_in_c_bypass_regNext_20_1_data_23;
  reg                 io_in_c_bypass_regNext_20_1_is_stationary_23;
  reg        [15:0]   io_in_c_bypass_regNext_20_2_data_23;
  reg                 io_in_c_bypass_regNext_20_2_is_stationary_23;
  reg        [15:0]   io_in_c_bypass_regNext_20_3_data_23;
  reg                 io_in_c_bypass_regNext_20_3_is_stationary_23;
  reg        [15:0]   io_in_c_bypass_regNext_21_0_data_23;
  reg                 io_in_c_bypass_regNext_21_0_is_stationary_23;
  reg        [15:0]   io_in_c_bypass_regNext_21_1_data_23;
  reg                 io_in_c_bypass_regNext_21_1_is_stationary_23;
  reg        [15:0]   io_in_c_bypass_regNext_21_2_data_23;
  reg                 io_in_c_bypass_regNext_21_2_is_stationary_23;
  reg        [15:0]   io_in_c_bypass_regNext_21_3_data_23;
  reg                 io_in_c_bypass_regNext_21_3_is_stationary_23;
  reg        [15:0]   io_in_c_bypass_regNext_22_0_data_23;
  reg                 io_in_c_bypass_regNext_22_0_is_stationary_23;
  reg        [15:0]   io_in_c_bypass_regNext_22_1_data_23;
  reg                 io_in_c_bypass_regNext_22_1_is_stationary_23;
  reg        [15:0]   io_in_c_bypass_regNext_22_2_data_23;
  reg                 io_in_c_bypass_regNext_22_2_is_stationary_23;
  reg        [15:0]   io_in_c_bypass_regNext_22_3_data_23;
  reg                 io_in_c_bypass_regNext_22_3_is_stationary_23;
  reg        [15:0]   io_in_c_bypass_regNext_23_0_data_23;
  reg                 io_in_c_bypass_regNext_23_0_is_stationary_23;
  reg        [15:0]   io_in_c_bypass_regNext_23_1_data_23;
  reg                 io_in_c_bypass_regNext_23_1_is_stationary_23;
  reg        [15:0]   io_in_c_bypass_regNext_23_2_data_23;
  reg                 io_in_c_bypass_regNext_23_2_is_stationary_23;
  reg        [15:0]   io_in_c_bypass_regNext_23_3_data_23;
  reg                 io_in_c_bypass_regNext_23_3_is_stationary_23;
  reg        [15:0]   io_in_c_bypass_regNext_24_0_data_23;
  reg                 io_in_c_bypass_regNext_24_0_is_stationary_23;
  reg        [15:0]   io_in_c_bypass_regNext_24_1_data_23;
  reg                 io_in_c_bypass_regNext_24_1_is_stationary_23;
  reg        [15:0]   io_in_c_bypass_regNext_24_2_data_23;
  reg                 io_in_c_bypass_regNext_24_2_is_stationary_23;
  reg        [15:0]   io_in_c_bypass_regNext_24_3_data_23;
  reg                 io_in_c_bypass_regNext_24_3_is_stationary_23;
  reg        [15:0]   io_in_c_bypass_regNext_25_0_data_23;
  reg                 io_in_c_bypass_regNext_25_0_is_stationary_23;
  reg        [15:0]   io_in_c_bypass_regNext_25_1_data_23;
  reg                 io_in_c_bypass_regNext_25_1_is_stationary_23;
  reg        [15:0]   io_in_c_bypass_regNext_25_2_data_23;
  reg                 io_in_c_bypass_regNext_25_2_is_stationary_23;
  reg        [15:0]   io_in_c_bypass_regNext_25_3_data_23;
  reg                 io_in_c_bypass_regNext_25_3_is_stationary_23;
  reg        [15:0]   io_in_c_bypass_regNext_26_0_data_23;
  reg                 io_in_c_bypass_regNext_26_0_is_stationary_23;
  reg        [15:0]   io_in_c_bypass_regNext_26_1_data_23;
  reg                 io_in_c_bypass_regNext_26_1_is_stationary_23;
  reg        [15:0]   io_in_c_bypass_regNext_26_2_data_23;
  reg                 io_in_c_bypass_regNext_26_2_is_stationary_23;
  reg        [15:0]   io_in_c_bypass_regNext_26_3_data_23;
  reg                 io_in_c_bypass_regNext_26_3_is_stationary_23;
  reg        [15:0]   io_in_c_bypass_regNext_27_0_data_23;
  reg                 io_in_c_bypass_regNext_27_0_is_stationary_23;
  reg        [15:0]   io_in_c_bypass_regNext_27_1_data_23;
  reg                 io_in_c_bypass_regNext_27_1_is_stationary_23;
  reg        [15:0]   io_in_c_bypass_regNext_27_2_data_23;
  reg                 io_in_c_bypass_regNext_27_2_is_stationary_23;
  reg        [15:0]   io_in_c_bypass_regNext_27_3_data_23;
  reg                 io_in_c_bypass_regNext_27_3_is_stationary_23;
  reg        [15:0]   io_in_c_bypass_regNext_28_0_data_23;
  reg                 io_in_c_bypass_regNext_28_0_is_stationary_23;
  reg        [15:0]   io_in_c_bypass_regNext_28_1_data_23;
  reg                 io_in_c_bypass_regNext_28_1_is_stationary_23;
  reg        [15:0]   io_in_c_bypass_regNext_28_2_data_23;
  reg                 io_in_c_bypass_regNext_28_2_is_stationary_23;
  reg        [15:0]   io_in_c_bypass_regNext_28_3_data_23;
  reg                 io_in_c_bypass_regNext_28_3_is_stationary_23;
  reg        [15:0]   io_in_c_bypass_regNext_29_0_data_23;
  reg                 io_in_c_bypass_regNext_29_0_is_stationary_23;
  reg        [15:0]   io_in_c_bypass_regNext_29_1_data_23;
  reg                 io_in_c_bypass_regNext_29_1_is_stationary_23;
  reg        [15:0]   io_in_c_bypass_regNext_29_2_data_23;
  reg                 io_in_c_bypass_regNext_29_2_is_stationary_23;
  reg        [15:0]   io_in_c_bypass_regNext_29_3_data_23;
  reg                 io_in_c_bypass_regNext_29_3_is_stationary_23;
  reg        [15:0]   io_in_c_bypass_regNext_30_0_data_23;
  reg                 io_in_c_bypass_regNext_30_0_is_stationary_23;
  reg        [15:0]   io_in_c_bypass_regNext_30_1_data_23;
  reg                 io_in_c_bypass_regNext_30_1_is_stationary_23;
  reg        [15:0]   io_in_c_bypass_regNext_30_2_data_23;
  reg                 io_in_c_bypass_regNext_30_2_is_stationary_23;
  reg        [15:0]   io_in_c_bypass_regNext_30_3_data_23;
  reg                 io_in_c_bypass_regNext_30_3_is_stationary_23;
  reg        [15:0]   io_in_c_bypass_regNext_31_0_data_23;
  reg                 io_in_c_bypass_regNext_31_0_is_stationary_23;
  reg        [15:0]   io_in_c_bypass_regNext_31_1_data_23;
  reg                 io_in_c_bypass_regNext_31_1_is_stationary_23;
  reg        [15:0]   io_in_c_bypass_regNext_31_2_data_23;
  reg                 io_in_c_bypass_regNext_31_2_is_stationary_23;
  reg        [15:0]   io_in_c_bypass_regNext_31_3_data_23;
  reg                 io_in_c_bypass_regNext_31_3_is_stationary_23;
  reg        [15:0]   io_in_c_bypass_regNext_0_0_data_24;
  reg                 io_in_c_bypass_regNext_0_0_is_stationary_24;
  reg        [15:0]   io_in_c_bypass_regNext_0_1_data_24;
  reg                 io_in_c_bypass_regNext_0_1_is_stationary_24;
  reg        [15:0]   io_in_c_bypass_regNext_0_2_data_24;
  reg                 io_in_c_bypass_regNext_0_2_is_stationary_24;
  reg        [15:0]   io_in_c_bypass_regNext_0_3_data_24;
  reg                 io_in_c_bypass_regNext_0_3_is_stationary_24;
  reg        [15:0]   io_in_c_bypass_regNext_1_0_data_24;
  reg                 io_in_c_bypass_regNext_1_0_is_stationary_24;
  reg        [15:0]   io_in_c_bypass_regNext_1_1_data_24;
  reg                 io_in_c_bypass_regNext_1_1_is_stationary_24;
  reg        [15:0]   io_in_c_bypass_regNext_1_2_data_24;
  reg                 io_in_c_bypass_regNext_1_2_is_stationary_24;
  reg        [15:0]   io_in_c_bypass_regNext_1_3_data_24;
  reg                 io_in_c_bypass_regNext_1_3_is_stationary_24;
  reg        [15:0]   io_in_c_bypass_regNext_2_0_data_24;
  reg                 io_in_c_bypass_regNext_2_0_is_stationary_24;
  reg        [15:0]   io_in_c_bypass_regNext_2_1_data_24;
  reg                 io_in_c_bypass_regNext_2_1_is_stationary_24;
  reg        [15:0]   io_in_c_bypass_regNext_2_2_data_24;
  reg                 io_in_c_bypass_regNext_2_2_is_stationary_24;
  reg        [15:0]   io_in_c_bypass_regNext_2_3_data_24;
  reg                 io_in_c_bypass_regNext_2_3_is_stationary_24;
  reg        [15:0]   io_in_c_bypass_regNext_3_0_data_24;
  reg                 io_in_c_bypass_regNext_3_0_is_stationary_24;
  reg        [15:0]   io_in_c_bypass_regNext_3_1_data_24;
  reg                 io_in_c_bypass_regNext_3_1_is_stationary_24;
  reg        [15:0]   io_in_c_bypass_regNext_3_2_data_24;
  reg                 io_in_c_bypass_regNext_3_2_is_stationary_24;
  reg        [15:0]   io_in_c_bypass_regNext_3_3_data_24;
  reg                 io_in_c_bypass_regNext_3_3_is_stationary_24;
  reg        [15:0]   io_in_c_bypass_regNext_4_0_data_24;
  reg                 io_in_c_bypass_regNext_4_0_is_stationary_24;
  reg        [15:0]   io_in_c_bypass_regNext_4_1_data_24;
  reg                 io_in_c_bypass_regNext_4_1_is_stationary_24;
  reg        [15:0]   io_in_c_bypass_regNext_4_2_data_24;
  reg                 io_in_c_bypass_regNext_4_2_is_stationary_24;
  reg        [15:0]   io_in_c_bypass_regNext_4_3_data_24;
  reg                 io_in_c_bypass_regNext_4_3_is_stationary_24;
  reg        [15:0]   io_in_c_bypass_regNext_5_0_data_24;
  reg                 io_in_c_bypass_regNext_5_0_is_stationary_24;
  reg        [15:0]   io_in_c_bypass_regNext_5_1_data_24;
  reg                 io_in_c_bypass_regNext_5_1_is_stationary_24;
  reg        [15:0]   io_in_c_bypass_regNext_5_2_data_24;
  reg                 io_in_c_bypass_regNext_5_2_is_stationary_24;
  reg        [15:0]   io_in_c_bypass_regNext_5_3_data_24;
  reg                 io_in_c_bypass_regNext_5_3_is_stationary_24;
  reg        [15:0]   io_in_c_bypass_regNext_6_0_data_24;
  reg                 io_in_c_bypass_regNext_6_0_is_stationary_24;
  reg        [15:0]   io_in_c_bypass_regNext_6_1_data_24;
  reg                 io_in_c_bypass_regNext_6_1_is_stationary_24;
  reg        [15:0]   io_in_c_bypass_regNext_6_2_data_24;
  reg                 io_in_c_bypass_regNext_6_2_is_stationary_24;
  reg        [15:0]   io_in_c_bypass_regNext_6_3_data_24;
  reg                 io_in_c_bypass_regNext_6_3_is_stationary_24;
  reg        [15:0]   io_in_c_bypass_regNext_7_0_data_24;
  reg                 io_in_c_bypass_regNext_7_0_is_stationary_24;
  reg        [15:0]   io_in_c_bypass_regNext_7_1_data_24;
  reg                 io_in_c_bypass_regNext_7_1_is_stationary_24;
  reg        [15:0]   io_in_c_bypass_regNext_7_2_data_24;
  reg                 io_in_c_bypass_regNext_7_2_is_stationary_24;
  reg        [15:0]   io_in_c_bypass_regNext_7_3_data_24;
  reg                 io_in_c_bypass_regNext_7_3_is_stationary_24;
  reg        [15:0]   io_in_c_bypass_regNext_8_0_data_24;
  reg                 io_in_c_bypass_regNext_8_0_is_stationary_24;
  reg        [15:0]   io_in_c_bypass_regNext_8_1_data_24;
  reg                 io_in_c_bypass_regNext_8_1_is_stationary_24;
  reg        [15:0]   io_in_c_bypass_regNext_8_2_data_24;
  reg                 io_in_c_bypass_regNext_8_2_is_stationary_24;
  reg        [15:0]   io_in_c_bypass_regNext_8_3_data_24;
  reg                 io_in_c_bypass_regNext_8_3_is_stationary_24;
  reg        [15:0]   io_in_c_bypass_regNext_9_0_data_24;
  reg                 io_in_c_bypass_regNext_9_0_is_stationary_24;
  reg        [15:0]   io_in_c_bypass_regNext_9_1_data_24;
  reg                 io_in_c_bypass_regNext_9_1_is_stationary_24;
  reg        [15:0]   io_in_c_bypass_regNext_9_2_data_24;
  reg                 io_in_c_bypass_regNext_9_2_is_stationary_24;
  reg        [15:0]   io_in_c_bypass_regNext_9_3_data_24;
  reg                 io_in_c_bypass_regNext_9_3_is_stationary_24;
  reg        [15:0]   io_in_c_bypass_regNext_10_0_data_24;
  reg                 io_in_c_bypass_regNext_10_0_is_stationary_24;
  reg        [15:0]   io_in_c_bypass_regNext_10_1_data_24;
  reg                 io_in_c_bypass_regNext_10_1_is_stationary_24;
  reg        [15:0]   io_in_c_bypass_regNext_10_2_data_24;
  reg                 io_in_c_bypass_regNext_10_2_is_stationary_24;
  reg        [15:0]   io_in_c_bypass_regNext_10_3_data_24;
  reg                 io_in_c_bypass_regNext_10_3_is_stationary_24;
  reg        [15:0]   io_in_c_bypass_regNext_11_0_data_24;
  reg                 io_in_c_bypass_regNext_11_0_is_stationary_24;
  reg        [15:0]   io_in_c_bypass_regNext_11_1_data_24;
  reg                 io_in_c_bypass_regNext_11_1_is_stationary_24;
  reg        [15:0]   io_in_c_bypass_regNext_11_2_data_24;
  reg                 io_in_c_bypass_regNext_11_2_is_stationary_24;
  reg        [15:0]   io_in_c_bypass_regNext_11_3_data_24;
  reg                 io_in_c_bypass_regNext_11_3_is_stationary_24;
  reg        [15:0]   io_in_c_bypass_regNext_12_0_data_24;
  reg                 io_in_c_bypass_regNext_12_0_is_stationary_24;
  reg        [15:0]   io_in_c_bypass_regNext_12_1_data_24;
  reg                 io_in_c_bypass_regNext_12_1_is_stationary_24;
  reg        [15:0]   io_in_c_bypass_regNext_12_2_data_24;
  reg                 io_in_c_bypass_regNext_12_2_is_stationary_24;
  reg        [15:0]   io_in_c_bypass_regNext_12_3_data_24;
  reg                 io_in_c_bypass_regNext_12_3_is_stationary_24;
  reg        [15:0]   io_in_c_bypass_regNext_13_0_data_24;
  reg                 io_in_c_bypass_regNext_13_0_is_stationary_24;
  reg        [15:0]   io_in_c_bypass_regNext_13_1_data_24;
  reg                 io_in_c_bypass_regNext_13_1_is_stationary_24;
  reg        [15:0]   io_in_c_bypass_regNext_13_2_data_24;
  reg                 io_in_c_bypass_regNext_13_2_is_stationary_24;
  reg        [15:0]   io_in_c_bypass_regNext_13_3_data_24;
  reg                 io_in_c_bypass_regNext_13_3_is_stationary_24;
  reg        [15:0]   io_in_c_bypass_regNext_14_0_data_24;
  reg                 io_in_c_bypass_regNext_14_0_is_stationary_24;
  reg        [15:0]   io_in_c_bypass_regNext_14_1_data_24;
  reg                 io_in_c_bypass_regNext_14_1_is_stationary_24;
  reg        [15:0]   io_in_c_bypass_regNext_14_2_data_24;
  reg                 io_in_c_bypass_regNext_14_2_is_stationary_24;
  reg        [15:0]   io_in_c_bypass_regNext_14_3_data_24;
  reg                 io_in_c_bypass_regNext_14_3_is_stationary_24;
  reg        [15:0]   io_in_c_bypass_regNext_15_0_data_24;
  reg                 io_in_c_bypass_regNext_15_0_is_stationary_24;
  reg        [15:0]   io_in_c_bypass_regNext_15_1_data_24;
  reg                 io_in_c_bypass_regNext_15_1_is_stationary_24;
  reg        [15:0]   io_in_c_bypass_regNext_15_2_data_24;
  reg                 io_in_c_bypass_regNext_15_2_is_stationary_24;
  reg        [15:0]   io_in_c_bypass_regNext_15_3_data_24;
  reg                 io_in_c_bypass_regNext_15_3_is_stationary_24;
  reg        [15:0]   io_in_c_bypass_regNext_16_0_data_24;
  reg                 io_in_c_bypass_regNext_16_0_is_stationary_24;
  reg        [15:0]   io_in_c_bypass_regNext_16_1_data_24;
  reg                 io_in_c_bypass_regNext_16_1_is_stationary_24;
  reg        [15:0]   io_in_c_bypass_regNext_16_2_data_24;
  reg                 io_in_c_bypass_regNext_16_2_is_stationary_24;
  reg        [15:0]   io_in_c_bypass_regNext_16_3_data_24;
  reg                 io_in_c_bypass_regNext_16_3_is_stationary_24;
  reg        [15:0]   io_in_c_bypass_regNext_17_0_data_24;
  reg                 io_in_c_bypass_regNext_17_0_is_stationary_24;
  reg        [15:0]   io_in_c_bypass_regNext_17_1_data_24;
  reg                 io_in_c_bypass_regNext_17_1_is_stationary_24;
  reg        [15:0]   io_in_c_bypass_regNext_17_2_data_24;
  reg                 io_in_c_bypass_regNext_17_2_is_stationary_24;
  reg        [15:0]   io_in_c_bypass_regNext_17_3_data_24;
  reg                 io_in_c_bypass_regNext_17_3_is_stationary_24;
  reg        [15:0]   io_in_c_bypass_regNext_18_0_data_24;
  reg                 io_in_c_bypass_regNext_18_0_is_stationary_24;
  reg        [15:0]   io_in_c_bypass_regNext_18_1_data_24;
  reg                 io_in_c_bypass_regNext_18_1_is_stationary_24;
  reg        [15:0]   io_in_c_bypass_regNext_18_2_data_24;
  reg                 io_in_c_bypass_regNext_18_2_is_stationary_24;
  reg        [15:0]   io_in_c_bypass_regNext_18_3_data_24;
  reg                 io_in_c_bypass_regNext_18_3_is_stationary_24;
  reg        [15:0]   io_in_c_bypass_regNext_19_0_data_24;
  reg                 io_in_c_bypass_regNext_19_0_is_stationary_24;
  reg        [15:0]   io_in_c_bypass_regNext_19_1_data_24;
  reg                 io_in_c_bypass_regNext_19_1_is_stationary_24;
  reg        [15:0]   io_in_c_bypass_regNext_19_2_data_24;
  reg                 io_in_c_bypass_regNext_19_2_is_stationary_24;
  reg        [15:0]   io_in_c_bypass_regNext_19_3_data_24;
  reg                 io_in_c_bypass_regNext_19_3_is_stationary_24;
  reg        [15:0]   io_in_c_bypass_regNext_20_0_data_24;
  reg                 io_in_c_bypass_regNext_20_0_is_stationary_24;
  reg        [15:0]   io_in_c_bypass_regNext_20_1_data_24;
  reg                 io_in_c_bypass_regNext_20_1_is_stationary_24;
  reg        [15:0]   io_in_c_bypass_regNext_20_2_data_24;
  reg                 io_in_c_bypass_regNext_20_2_is_stationary_24;
  reg        [15:0]   io_in_c_bypass_regNext_20_3_data_24;
  reg                 io_in_c_bypass_regNext_20_3_is_stationary_24;
  reg        [15:0]   io_in_c_bypass_regNext_21_0_data_24;
  reg                 io_in_c_bypass_regNext_21_0_is_stationary_24;
  reg        [15:0]   io_in_c_bypass_regNext_21_1_data_24;
  reg                 io_in_c_bypass_regNext_21_1_is_stationary_24;
  reg        [15:0]   io_in_c_bypass_regNext_21_2_data_24;
  reg                 io_in_c_bypass_regNext_21_2_is_stationary_24;
  reg        [15:0]   io_in_c_bypass_regNext_21_3_data_24;
  reg                 io_in_c_bypass_regNext_21_3_is_stationary_24;
  reg        [15:0]   io_in_c_bypass_regNext_22_0_data_24;
  reg                 io_in_c_bypass_regNext_22_0_is_stationary_24;
  reg        [15:0]   io_in_c_bypass_regNext_22_1_data_24;
  reg                 io_in_c_bypass_regNext_22_1_is_stationary_24;
  reg        [15:0]   io_in_c_bypass_regNext_22_2_data_24;
  reg                 io_in_c_bypass_regNext_22_2_is_stationary_24;
  reg        [15:0]   io_in_c_bypass_regNext_22_3_data_24;
  reg                 io_in_c_bypass_regNext_22_3_is_stationary_24;
  reg        [15:0]   io_in_c_bypass_regNext_23_0_data_24;
  reg                 io_in_c_bypass_regNext_23_0_is_stationary_24;
  reg        [15:0]   io_in_c_bypass_regNext_23_1_data_24;
  reg                 io_in_c_bypass_regNext_23_1_is_stationary_24;
  reg        [15:0]   io_in_c_bypass_regNext_23_2_data_24;
  reg                 io_in_c_bypass_regNext_23_2_is_stationary_24;
  reg        [15:0]   io_in_c_bypass_regNext_23_3_data_24;
  reg                 io_in_c_bypass_regNext_23_3_is_stationary_24;
  reg        [15:0]   io_in_c_bypass_regNext_24_0_data_24;
  reg                 io_in_c_bypass_regNext_24_0_is_stationary_24;
  reg        [15:0]   io_in_c_bypass_regNext_24_1_data_24;
  reg                 io_in_c_bypass_regNext_24_1_is_stationary_24;
  reg        [15:0]   io_in_c_bypass_regNext_24_2_data_24;
  reg                 io_in_c_bypass_regNext_24_2_is_stationary_24;
  reg        [15:0]   io_in_c_bypass_regNext_24_3_data_24;
  reg                 io_in_c_bypass_regNext_24_3_is_stationary_24;
  reg        [15:0]   io_in_c_bypass_regNext_25_0_data_24;
  reg                 io_in_c_bypass_regNext_25_0_is_stationary_24;
  reg        [15:0]   io_in_c_bypass_regNext_25_1_data_24;
  reg                 io_in_c_bypass_regNext_25_1_is_stationary_24;
  reg        [15:0]   io_in_c_bypass_regNext_25_2_data_24;
  reg                 io_in_c_bypass_regNext_25_2_is_stationary_24;
  reg        [15:0]   io_in_c_bypass_regNext_25_3_data_24;
  reg                 io_in_c_bypass_regNext_25_3_is_stationary_24;
  reg        [15:0]   io_in_c_bypass_regNext_26_0_data_24;
  reg                 io_in_c_bypass_regNext_26_0_is_stationary_24;
  reg        [15:0]   io_in_c_bypass_regNext_26_1_data_24;
  reg                 io_in_c_bypass_regNext_26_1_is_stationary_24;
  reg        [15:0]   io_in_c_bypass_regNext_26_2_data_24;
  reg                 io_in_c_bypass_regNext_26_2_is_stationary_24;
  reg        [15:0]   io_in_c_bypass_regNext_26_3_data_24;
  reg                 io_in_c_bypass_regNext_26_3_is_stationary_24;
  reg        [15:0]   io_in_c_bypass_regNext_27_0_data_24;
  reg                 io_in_c_bypass_regNext_27_0_is_stationary_24;
  reg        [15:0]   io_in_c_bypass_regNext_27_1_data_24;
  reg                 io_in_c_bypass_regNext_27_1_is_stationary_24;
  reg        [15:0]   io_in_c_bypass_regNext_27_2_data_24;
  reg                 io_in_c_bypass_regNext_27_2_is_stationary_24;
  reg        [15:0]   io_in_c_bypass_regNext_27_3_data_24;
  reg                 io_in_c_bypass_regNext_27_3_is_stationary_24;
  reg        [15:0]   io_in_c_bypass_regNext_28_0_data_24;
  reg                 io_in_c_bypass_regNext_28_0_is_stationary_24;
  reg        [15:0]   io_in_c_bypass_regNext_28_1_data_24;
  reg                 io_in_c_bypass_regNext_28_1_is_stationary_24;
  reg        [15:0]   io_in_c_bypass_regNext_28_2_data_24;
  reg                 io_in_c_bypass_regNext_28_2_is_stationary_24;
  reg        [15:0]   io_in_c_bypass_regNext_28_3_data_24;
  reg                 io_in_c_bypass_regNext_28_3_is_stationary_24;
  reg        [15:0]   io_in_c_bypass_regNext_29_0_data_24;
  reg                 io_in_c_bypass_regNext_29_0_is_stationary_24;
  reg        [15:0]   io_in_c_bypass_regNext_29_1_data_24;
  reg                 io_in_c_bypass_regNext_29_1_is_stationary_24;
  reg        [15:0]   io_in_c_bypass_regNext_29_2_data_24;
  reg                 io_in_c_bypass_regNext_29_2_is_stationary_24;
  reg        [15:0]   io_in_c_bypass_regNext_29_3_data_24;
  reg                 io_in_c_bypass_regNext_29_3_is_stationary_24;
  reg        [15:0]   io_in_c_bypass_regNext_30_0_data_24;
  reg                 io_in_c_bypass_regNext_30_0_is_stationary_24;
  reg        [15:0]   io_in_c_bypass_regNext_30_1_data_24;
  reg                 io_in_c_bypass_regNext_30_1_is_stationary_24;
  reg        [15:0]   io_in_c_bypass_regNext_30_2_data_24;
  reg                 io_in_c_bypass_regNext_30_2_is_stationary_24;
  reg        [15:0]   io_in_c_bypass_regNext_30_3_data_24;
  reg                 io_in_c_bypass_regNext_30_3_is_stationary_24;
  reg        [15:0]   io_in_c_bypass_regNext_31_0_data_24;
  reg                 io_in_c_bypass_regNext_31_0_is_stationary_24;
  reg        [15:0]   io_in_c_bypass_regNext_31_1_data_24;
  reg                 io_in_c_bypass_regNext_31_1_is_stationary_24;
  reg        [15:0]   io_in_c_bypass_regNext_31_2_data_24;
  reg                 io_in_c_bypass_regNext_31_2_is_stationary_24;
  reg        [15:0]   io_in_c_bypass_regNext_31_3_data_24;
  reg                 io_in_c_bypass_regNext_31_3_is_stationary_24;
  reg        [15:0]   io_in_c_bypass_regNext_0_0_data_25;
  reg                 io_in_c_bypass_regNext_0_0_is_stationary_25;
  reg        [15:0]   io_in_c_bypass_regNext_0_1_data_25;
  reg                 io_in_c_bypass_regNext_0_1_is_stationary_25;
  reg        [15:0]   io_in_c_bypass_regNext_0_2_data_25;
  reg                 io_in_c_bypass_regNext_0_2_is_stationary_25;
  reg        [15:0]   io_in_c_bypass_regNext_0_3_data_25;
  reg                 io_in_c_bypass_regNext_0_3_is_stationary_25;
  reg        [15:0]   io_in_c_bypass_regNext_1_0_data_25;
  reg                 io_in_c_bypass_regNext_1_0_is_stationary_25;
  reg        [15:0]   io_in_c_bypass_regNext_1_1_data_25;
  reg                 io_in_c_bypass_regNext_1_1_is_stationary_25;
  reg        [15:0]   io_in_c_bypass_regNext_1_2_data_25;
  reg                 io_in_c_bypass_regNext_1_2_is_stationary_25;
  reg        [15:0]   io_in_c_bypass_regNext_1_3_data_25;
  reg                 io_in_c_bypass_regNext_1_3_is_stationary_25;
  reg        [15:0]   io_in_c_bypass_regNext_2_0_data_25;
  reg                 io_in_c_bypass_regNext_2_0_is_stationary_25;
  reg        [15:0]   io_in_c_bypass_regNext_2_1_data_25;
  reg                 io_in_c_bypass_regNext_2_1_is_stationary_25;
  reg        [15:0]   io_in_c_bypass_regNext_2_2_data_25;
  reg                 io_in_c_bypass_regNext_2_2_is_stationary_25;
  reg        [15:0]   io_in_c_bypass_regNext_2_3_data_25;
  reg                 io_in_c_bypass_regNext_2_3_is_stationary_25;
  reg        [15:0]   io_in_c_bypass_regNext_3_0_data_25;
  reg                 io_in_c_bypass_regNext_3_0_is_stationary_25;
  reg        [15:0]   io_in_c_bypass_regNext_3_1_data_25;
  reg                 io_in_c_bypass_regNext_3_1_is_stationary_25;
  reg        [15:0]   io_in_c_bypass_regNext_3_2_data_25;
  reg                 io_in_c_bypass_regNext_3_2_is_stationary_25;
  reg        [15:0]   io_in_c_bypass_regNext_3_3_data_25;
  reg                 io_in_c_bypass_regNext_3_3_is_stationary_25;
  reg        [15:0]   io_in_c_bypass_regNext_4_0_data_25;
  reg                 io_in_c_bypass_regNext_4_0_is_stationary_25;
  reg        [15:0]   io_in_c_bypass_regNext_4_1_data_25;
  reg                 io_in_c_bypass_regNext_4_1_is_stationary_25;
  reg        [15:0]   io_in_c_bypass_regNext_4_2_data_25;
  reg                 io_in_c_bypass_regNext_4_2_is_stationary_25;
  reg        [15:0]   io_in_c_bypass_regNext_4_3_data_25;
  reg                 io_in_c_bypass_regNext_4_3_is_stationary_25;
  reg        [15:0]   io_in_c_bypass_regNext_5_0_data_25;
  reg                 io_in_c_bypass_regNext_5_0_is_stationary_25;
  reg        [15:0]   io_in_c_bypass_regNext_5_1_data_25;
  reg                 io_in_c_bypass_regNext_5_1_is_stationary_25;
  reg        [15:0]   io_in_c_bypass_regNext_5_2_data_25;
  reg                 io_in_c_bypass_regNext_5_2_is_stationary_25;
  reg        [15:0]   io_in_c_bypass_regNext_5_3_data_25;
  reg                 io_in_c_bypass_regNext_5_3_is_stationary_25;
  reg        [15:0]   io_in_c_bypass_regNext_6_0_data_25;
  reg                 io_in_c_bypass_regNext_6_0_is_stationary_25;
  reg        [15:0]   io_in_c_bypass_regNext_6_1_data_25;
  reg                 io_in_c_bypass_regNext_6_1_is_stationary_25;
  reg        [15:0]   io_in_c_bypass_regNext_6_2_data_25;
  reg                 io_in_c_bypass_regNext_6_2_is_stationary_25;
  reg        [15:0]   io_in_c_bypass_regNext_6_3_data_25;
  reg                 io_in_c_bypass_regNext_6_3_is_stationary_25;
  reg        [15:0]   io_in_c_bypass_regNext_7_0_data_25;
  reg                 io_in_c_bypass_regNext_7_0_is_stationary_25;
  reg        [15:0]   io_in_c_bypass_regNext_7_1_data_25;
  reg                 io_in_c_bypass_regNext_7_1_is_stationary_25;
  reg        [15:0]   io_in_c_bypass_regNext_7_2_data_25;
  reg                 io_in_c_bypass_regNext_7_2_is_stationary_25;
  reg        [15:0]   io_in_c_bypass_regNext_7_3_data_25;
  reg                 io_in_c_bypass_regNext_7_3_is_stationary_25;
  reg        [15:0]   io_in_c_bypass_regNext_8_0_data_25;
  reg                 io_in_c_bypass_regNext_8_0_is_stationary_25;
  reg        [15:0]   io_in_c_bypass_regNext_8_1_data_25;
  reg                 io_in_c_bypass_regNext_8_1_is_stationary_25;
  reg        [15:0]   io_in_c_bypass_regNext_8_2_data_25;
  reg                 io_in_c_bypass_regNext_8_2_is_stationary_25;
  reg        [15:0]   io_in_c_bypass_regNext_8_3_data_25;
  reg                 io_in_c_bypass_regNext_8_3_is_stationary_25;
  reg        [15:0]   io_in_c_bypass_regNext_9_0_data_25;
  reg                 io_in_c_bypass_regNext_9_0_is_stationary_25;
  reg        [15:0]   io_in_c_bypass_regNext_9_1_data_25;
  reg                 io_in_c_bypass_regNext_9_1_is_stationary_25;
  reg        [15:0]   io_in_c_bypass_regNext_9_2_data_25;
  reg                 io_in_c_bypass_regNext_9_2_is_stationary_25;
  reg        [15:0]   io_in_c_bypass_regNext_9_3_data_25;
  reg                 io_in_c_bypass_regNext_9_3_is_stationary_25;
  reg        [15:0]   io_in_c_bypass_regNext_10_0_data_25;
  reg                 io_in_c_bypass_regNext_10_0_is_stationary_25;
  reg        [15:0]   io_in_c_bypass_regNext_10_1_data_25;
  reg                 io_in_c_bypass_regNext_10_1_is_stationary_25;
  reg        [15:0]   io_in_c_bypass_regNext_10_2_data_25;
  reg                 io_in_c_bypass_regNext_10_2_is_stationary_25;
  reg        [15:0]   io_in_c_bypass_regNext_10_3_data_25;
  reg                 io_in_c_bypass_regNext_10_3_is_stationary_25;
  reg        [15:0]   io_in_c_bypass_regNext_11_0_data_25;
  reg                 io_in_c_bypass_regNext_11_0_is_stationary_25;
  reg        [15:0]   io_in_c_bypass_regNext_11_1_data_25;
  reg                 io_in_c_bypass_regNext_11_1_is_stationary_25;
  reg        [15:0]   io_in_c_bypass_regNext_11_2_data_25;
  reg                 io_in_c_bypass_regNext_11_2_is_stationary_25;
  reg        [15:0]   io_in_c_bypass_regNext_11_3_data_25;
  reg                 io_in_c_bypass_regNext_11_3_is_stationary_25;
  reg        [15:0]   io_in_c_bypass_regNext_12_0_data_25;
  reg                 io_in_c_bypass_regNext_12_0_is_stationary_25;
  reg        [15:0]   io_in_c_bypass_regNext_12_1_data_25;
  reg                 io_in_c_bypass_regNext_12_1_is_stationary_25;
  reg        [15:0]   io_in_c_bypass_regNext_12_2_data_25;
  reg                 io_in_c_bypass_regNext_12_2_is_stationary_25;
  reg        [15:0]   io_in_c_bypass_regNext_12_3_data_25;
  reg                 io_in_c_bypass_regNext_12_3_is_stationary_25;
  reg        [15:0]   io_in_c_bypass_regNext_13_0_data_25;
  reg                 io_in_c_bypass_regNext_13_0_is_stationary_25;
  reg        [15:0]   io_in_c_bypass_regNext_13_1_data_25;
  reg                 io_in_c_bypass_regNext_13_1_is_stationary_25;
  reg        [15:0]   io_in_c_bypass_regNext_13_2_data_25;
  reg                 io_in_c_bypass_regNext_13_2_is_stationary_25;
  reg        [15:0]   io_in_c_bypass_regNext_13_3_data_25;
  reg                 io_in_c_bypass_regNext_13_3_is_stationary_25;
  reg        [15:0]   io_in_c_bypass_regNext_14_0_data_25;
  reg                 io_in_c_bypass_regNext_14_0_is_stationary_25;
  reg        [15:0]   io_in_c_bypass_regNext_14_1_data_25;
  reg                 io_in_c_bypass_regNext_14_1_is_stationary_25;
  reg        [15:0]   io_in_c_bypass_regNext_14_2_data_25;
  reg                 io_in_c_bypass_regNext_14_2_is_stationary_25;
  reg        [15:0]   io_in_c_bypass_regNext_14_3_data_25;
  reg                 io_in_c_bypass_regNext_14_3_is_stationary_25;
  reg        [15:0]   io_in_c_bypass_regNext_15_0_data_25;
  reg                 io_in_c_bypass_regNext_15_0_is_stationary_25;
  reg        [15:0]   io_in_c_bypass_regNext_15_1_data_25;
  reg                 io_in_c_bypass_regNext_15_1_is_stationary_25;
  reg        [15:0]   io_in_c_bypass_regNext_15_2_data_25;
  reg                 io_in_c_bypass_regNext_15_2_is_stationary_25;
  reg        [15:0]   io_in_c_bypass_regNext_15_3_data_25;
  reg                 io_in_c_bypass_regNext_15_3_is_stationary_25;
  reg        [15:0]   io_in_c_bypass_regNext_16_0_data_25;
  reg                 io_in_c_bypass_regNext_16_0_is_stationary_25;
  reg        [15:0]   io_in_c_bypass_regNext_16_1_data_25;
  reg                 io_in_c_bypass_regNext_16_1_is_stationary_25;
  reg        [15:0]   io_in_c_bypass_regNext_16_2_data_25;
  reg                 io_in_c_bypass_regNext_16_2_is_stationary_25;
  reg        [15:0]   io_in_c_bypass_regNext_16_3_data_25;
  reg                 io_in_c_bypass_regNext_16_3_is_stationary_25;
  reg        [15:0]   io_in_c_bypass_regNext_17_0_data_25;
  reg                 io_in_c_bypass_regNext_17_0_is_stationary_25;
  reg        [15:0]   io_in_c_bypass_regNext_17_1_data_25;
  reg                 io_in_c_bypass_regNext_17_1_is_stationary_25;
  reg        [15:0]   io_in_c_bypass_regNext_17_2_data_25;
  reg                 io_in_c_bypass_regNext_17_2_is_stationary_25;
  reg        [15:0]   io_in_c_bypass_regNext_17_3_data_25;
  reg                 io_in_c_bypass_regNext_17_3_is_stationary_25;
  reg        [15:0]   io_in_c_bypass_regNext_18_0_data_25;
  reg                 io_in_c_bypass_regNext_18_0_is_stationary_25;
  reg        [15:0]   io_in_c_bypass_regNext_18_1_data_25;
  reg                 io_in_c_bypass_regNext_18_1_is_stationary_25;
  reg        [15:0]   io_in_c_bypass_regNext_18_2_data_25;
  reg                 io_in_c_bypass_regNext_18_2_is_stationary_25;
  reg        [15:0]   io_in_c_bypass_regNext_18_3_data_25;
  reg                 io_in_c_bypass_regNext_18_3_is_stationary_25;
  reg        [15:0]   io_in_c_bypass_regNext_19_0_data_25;
  reg                 io_in_c_bypass_regNext_19_0_is_stationary_25;
  reg        [15:0]   io_in_c_bypass_regNext_19_1_data_25;
  reg                 io_in_c_bypass_regNext_19_1_is_stationary_25;
  reg        [15:0]   io_in_c_bypass_regNext_19_2_data_25;
  reg                 io_in_c_bypass_regNext_19_2_is_stationary_25;
  reg        [15:0]   io_in_c_bypass_regNext_19_3_data_25;
  reg                 io_in_c_bypass_regNext_19_3_is_stationary_25;
  reg        [15:0]   io_in_c_bypass_regNext_20_0_data_25;
  reg                 io_in_c_bypass_regNext_20_0_is_stationary_25;
  reg        [15:0]   io_in_c_bypass_regNext_20_1_data_25;
  reg                 io_in_c_bypass_regNext_20_1_is_stationary_25;
  reg        [15:0]   io_in_c_bypass_regNext_20_2_data_25;
  reg                 io_in_c_bypass_regNext_20_2_is_stationary_25;
  reg        [15:0]   io_in_c_bypass_regNext_20_3_data_25;
  reg                 io_in_c_bypass_regNext_20_3_is_stationary_25;
  reg        [15:0]   io_in_c_bypass_regNext_21_0_data_25;
  reg                 io_in_c_bypass_regNext_21_0_is_stationary_25;
  reg        [15:0]   io_in_c_bypass_regNext_21_1_data_25;
  reg                 io_in_c_bypass_regNext_21_1_is_stationary_25;
  reg        [15:0]   io_in_c_bypass_regNext_21_2_data_25;
  reg                 io_in_c_bypass_regNext_21_2_is_stationary_25;
  reg        [15:0]   io_in_c_bypass_regNext_21_3_data_25;
  reg                 io_in_c_bypass_regNext_21_3_is_stationary_25;
  reg        [15:0]   io_in_c_bypass_regNext_22_0_data_25;
  reg                 io_in_c_bypass_regNext_22_0_is_stationary_25;
  reg        [15:0]   io_in_c_bypass_regNext_22_1_data_25;
  reg                 io_in_c_bypass_regNext_22_1_is_stationary_25;
  reg        [15:0]   io_in_c_bypass_regNext_22_2_data_25;
  reg                 io_in_c_bypass_regNext_22_2_is_stationary_25;
  reg        [15:0]   io_in_c_bypass_regNext_22_3_data_25;
  reg                 io_in_c_bypass_regNext_22_3_is_stationary_25;
  reg        [15:0]   io_in_c_bypass_regNext_23_0_data_25;
  reg                 io_in_c_bypass_regNext_23_0_is_stationary_25;
  reg        [15:0]   io_in_c_bypass_regNext_23_1_data_25;
  reg                 io_in_c_bypass_regNext_23_1_is_stationary_25;
  reg        [15:0]   io_in_c_bypass_regNext_23_2_data_25;
  reg                 io_in_c_bypass_regNext_23_2_is_stationary_25;
  reg        [15:0]   io_in_c_bypass_regNext_23_3_data_25;
  reg                 io_in_c_bypass_regNext_23_3_is_stationary_25;
  reg        [15:0]   io_in_c_bypass_regNext_24_0_data_25;
  reg                 io_in_c_bypass_regNext_24_0_is_stationary_25;
  reg        [15:0]   io_in_c_bypass_regNext_24_1_data_25;
  reg                 io_in_c_bypass_regNext_24_1_is_stationary_25;
  reg        [15:0]   io_in_c_bypass_regNext_24_2_data_25;
  reg                 io_in_c_bypass_regNext_24_2_is_stationary_25;
  reg        [15:0]   io_in_c_bypass_regNext_24_3_data_25;
  reg                 io_in_c_bypass_regNext_24_3_is_stationary_25;
  reg        [15:0]   io_in_c_bypass_regNext_25_0_data_25;
  reg                 io_in_c_bypass_regNext_25_0_is_stationary_25;
  reg        [15:0]   io_in_c_bypass_regNext_25_1_data_25;
  reg                 io_in_c_bypass_regNext_25_1_is_stationary_25;
  reg        [15:0]   io_in_c_bypass_regNext_25_2_data_25;
  reg                 io_in_c_bypass_regNext_25_2_is_stationary_25;
  reg        [15:0]   io_in_c_bypass_regNext_25_3_data_25;
  reg                 io_in_c_bypass_regNext_25_3_is_stationary_25;
  reg        [15:0]   io_in_c_bypass_regNext_26_0_data_25;
  reg                 io_in_c_bypass_regNext_26_0_is_stationary_25;
  reg        [15:0]   io_in_c_bypass_regNext_26_1_data_25;
  reg                 io_in_c_bypass_regNext_26_1_is_stationary_25;
  reg        [15:0]   io_in_c_bypass_regNext_26_2_data_25;
  reg                 io_in_c_bypass_regNext_26_2_is_stationary_25;
  reg        [15:0]   io_in_c_bypass_regNext_26_3_data_25;
  reg                 io_in_c_bypass_regNext_26_3_is_stationary_25;
  reg        [15:0]   io_in_c_bypass_regNext_27_0_data_25;
  reg                 io_in_c_bypass_regNext_27_0_is_stationary_25;
  reg        [15:0]   io_in_c_bypass_regNext_27_1_data_25;
  reg                 io_in_c_bypass_regNext_27_1_is_stationary_25;
  reg        [15:0]   io_in_c_bypass_regNext_27_2_data_25;
  reg                 io_in_c_bypass_regNext_27_2_is_stationary_25;
  reg        [15:0]   io_in_c_bypass_regNext_27_3_data_25;
  reg                 io_in_c_bypass_regNext_27_3_is_stationary_25;
  reg        [15:0]   io_in_c_bypass_regNext_28_0_data_25;
  reg                 io_in_c_bypass_regNext_28_0_is_stationary_25;
  reg        [15:0]   io_in_c_bypass_regNext_28_1_data_25;
  reg                 io_in_c_bypass_regNext_28_1_is_stationary_25;
  reg        [15:0]   io_in_c_bypass_regNext_28_2_data_25;
  reg                 io_in_c_bypass_regNext_28_2_is_stationary_25;
  reg        [15:0]   io_in_c_bypass_regNext_28_3_data_25;
  reg                 io_in_c_bypass_regNext_28_3_is_stationary_25;
  reg        [15:0]   io_in_c_bypass_regNext_29_0_data_25;
  reg                 io_in_c_bypass_regNext_29_0_is_stationary_25;
  reg        [15:0]   io_in_c_bypass_regNext_29_1_data_25;
  reg                 io_in_c_bypass_regNext_29_1_is_stationary_25;
  reg        [15:0]   io_in_c_bypass_regNext_29_2_data_25;
  reg                 io_in_c_bypass_regNext_29_2_is_stationary_25;
  reg        [15:0]   io_in_c_bypass_regNext_29_3_data_25;
  reg                 io_in_c_bypass_regNext_29_3_is_stationary_25;
  reg        [15:0]   io_in_c_bypass_regNext_30_0_data_25;
  reg                 io_in_c_bypass_regNext_30_0_is_stationary_25;
  reg        [15:0]   io_in_c_bypass_regNext_30_1_data_25;
  reg                 io_in_c_bypass_regNext_30_1_is_stationary_25;
  reg        [15:0]   io_in_c_bypass_regNext_30_2_data_25;
  reg                 io_in_c_bypass_regNext_30_2_is_stationary_25;
  reg        [15:0]   io_in_c_bypass_regNext_30_3_data_25;
  reg                 io_in_c_bypass_regNext_30_3_is_stationary_25;
  reg        [15:0]   io_in_c_bypass_regNext_31_0_data_25;
  reg                 io_in_c_bypass_regNext_31_0_is_stationary_25;
  reg        [15:0]   io_in_c_bypass_regNext_31_1_data_25;
  reg                 io_in_c_bypass_regNext_31_1_is_stationary_25;
  reg        [15:0]   io_in_c_bypass_regNext_31_2_data_25;
  reg                 io_in_c_bypass_regNext_31_2_is_stationary_25;
  reg        [15:0]   io_in_c_bypass_regNext_31_3_data_25;
  reg                 io_in_c_bypass_regNext_31_3_is_stationary_25;
  reg        [15:0]   io_in_c_bypass_regNext_0_0_data_26;
  reg                 io_in_c_bypass_regNext_0_0_is_stationary_26;
  reg        [15:0]   io_in_c_bypass_regNext_0_1_data_26;
  reg                 io_in_c_bypass_regNext_0_1_is_stationary_26;
  reg        [15:0]   io_in_c_bypass_regNext_0_2_data_26;
  reg                 io_in_c_bypass_regNext_0_2_is_stationary_26;
  reg        [15:0]   io_in_c_bypass_regNext_0_3_data_26;
  reg                 io_in_c_bypass_regNext_0_3_is_stationary_26;
  reg        [15:0]   io_in_c_bypass_regNext_1_0_data_26;
  reg                 io_in_c_bypass_regNext_1_0_is_stationary_26;
  reg        [15:0]   io_in_c_bypass_regNext_1_1_data_26;
  reg                 io_in_c_bypass_regNext_1_1_is_stationary_26;
  reg        [15:0]   io_in_c_bypass_regNext_1_2_data_26;
  reg                 io_in_c_bypass_regNext_1_2_is_stationary_26;
  reg        [15:0]   io_in_c_bypass_regNext_1_3_data_26;
  reg                 io_in_c_bypass_regNext_1_3_is_stationary_26;
  reg        [15:0]   io_in_c_bypass_regNext_2_0_data_26;
  reg                 io_in_c_bypass_regNext_2_0_is_stationary_26;
  reg        [15:0]   io_in_c_bypass_regNext_2_1_data_26;
  reg                 io_in_c_bypass_regNext_2_1_is_stationary_26;
  reg        [15:0]   io_in_c_bypass_regNext_2_2_data_26;
  reg                 io_in_c_bypass_regNext_2_2_is_stationary_26;
  reg        [15:0]   io_in_c_bypass_regNext_2_3_data_26;
  reg                 io_in_c_bypass_regNext_2_3_is_stationary_26;
  reg        [15:0]   io_in_c_bypass_regNext_3_0_data_26;
  reg                 io_in_c_bypass_regNext_3_0_is_stationary_26;
  reg        [15:0]   io_in_c_bypass_regNext_3_1_data_26;
  reg                 io_in_c_bypass_regNext_3_1_is_stationary_26;
  reg        [15:0]   io_in_c_bypass_regNext_3_2_data_26;
  reg                 io_in_c_bypass_regNext_3_2_is_stationary_26;
  reg        [15:0]   io_in_c_bypass_regNext_3_3_data_26;
  reg                 io_in_c_bypass_regNext_3_3_is_stationary_26;
  reg        [15:0]   io_in_c_bypass_regNext_4_0_data_26;
  reg                 io_in_c_bypass_regNext_4_0_is_stationary_26;
  reg        [15:0]   io_in_c_bypass_regNext_4_1_data_26;
  reg                 io_in_c_bypass_regNext_4_1_is_stationary_26;
  reg        [15:0]   io_in_c_bypass_regNext_4_2_data_26;
  reg                 io_in_c_bypass_regNext_4_2_is_stationary_26;
  reg        [15:0]   io_in_c_bypass_regNext_4_3_data_26;
  reg                 io_in_c_bypass_regNext_4_3_is_stationary_26;
  reg        [15:0]   io_in_c_bypass_regNext_5_0_data_26;
  reg                 io_in_c_bypass_regNext_5_0_is_stationary_26;
  reg        [15:0]   io_in_c_bypass_regNext_5_1_data_26;
  reg                 io_in_c_bypass_regNext_5_1_is_stationary_26;
  reg        [15:0]   io_in_c_bypass_regNext_5_2_data_26;
  reg                 io_in_c_bypass_regNext_5_2_is_stationary_26;
  reg        [15:0]   io_in_c_bypass_regNext_5_3_data_26;
  reg                 io_in_c_bypass_regNext_5_3_is_stationary_26;
  reg        [15:0]   io_in_c_bypass_regNext_6_0_data_26;
  reg                 io_in_c_bypass_regNext_6_0_is_stationary_26;
  reg        [15:0]   io_in_c_bypass_regNext_6_1_data_26;
  reg                 io_in_c_bypass_regNext_6_1_is_stationary_26;
  reg        [15:0]   io_in_c_bypass_regNext_6_2_data_26;
  reg                 io_in_c_bypass_regNext_6_2_is_stationary_26;
  reg        [15:0]   io_in_c_bypass_regNext_6_3_data_26;
  reg                 io_in_c_bypass_regNext_6_3_is_stationary_26;
  reg        [15:0]   io_in_c_bypass_regNext_7_0_data_26;
  reg                 io_in_c_bypass_regNext_7_0_is_stationary_26;
  reg        [15:0]   io_in_c_bypass_regNext_7_1_data_26;
  reg                 io_in_c_bypass_regNext_7_1_is_stationary_26;
  reg        [15:0]   io_in_c_bypass_regNext_7_2_data_26;
  reg                 io_in_c_bypass_regNext_7_2_is_stationary_26;
  reg        [15:0]   io_in_c_bypass_regNext_7_3_data_26;
  reg                 io_in_c_bypass_regNext_7_3_is_stationary_26;
  reg        [15:0]   io_in_c_bypass_regNext_8_0_data_26;
  reg                 io_in_c_bypass_regNext_8_0_is_stationary_26;
  reg        [15:0]   io_in_c_bypass_regNext_8_1_data_26;
  reg                 io_in_c_bypass_regNext_8_1_is_stationary_26;
  reg        [15:0]   io_in_c_bypass_regNext_8_2_data_26;
  reg                 io_in_c_bypass_regNext_8_2_is_stationary_26;
  reg        [15:0]   io_in_c_bypass_regNext_8_3_data_26;
  reg                 io_in_c_bypass_regNext_8_3_is_stationary_26;
  reg        [15:0]   io_in_c_bypass_regNext_9_0_data_26;
  reg                 io_in_c_bypass_regNext_9_0_is_stationary_26;
  reg        [15:0]   io_in_c_bypass_regNext_9_1_data_26;
  reg                 io_in_c_bypass_regNext_9_1_is_stationary_26;
  reg        [15:0]   io_in_c_bypass_regNext_9_2_data_26;
  reg                 io_in_c_bypass_regNext_9_2_is_stationary_26;
  reg        [15:0]   io_in_c_bypass_regNext_9_3_data_26;
  reg                 io_in_c_bypass_regNext_9_3_is_stationary_26;
  reg        [15:0]   io_in_c_bypass_regNext_10_0_data_26;
  reg                 io_in_c_bypass_regNext_10_0_is_stationary_26;
  reg        [15:0]   io_in_c_bypass_regNext_10_1_data_26;
  reg                 io_in_c_bypass_regNext_10_1_is_stationary_26;
  reg        [15:0]   io_in_c_bypass_regNext_10_2_data_26;
  reg                 io_in_c_bypass_regNext_10_2_is_stationary_26;
  reg        [15:0]   io_in_c_bypass_regNext_10_3_data_26;
  reg                 io_in_c_bypass_regNext_10_3_is_stationary_26;
  reg        [15:0]   io_in_c_bypass_regNext_11_0_data_26;
  reg                 io_in_c_bypass_regNext_11_0_is_stationary_26;
  reg        [15:0]   io_in_c_bypass_regNext_11_1_data_26;
  reg                 io_in_c_bypass_regNext_11_1_is_stationary_26;
  reg        [15:0]   io_in_c_bypass_regNext_11_2_data_26;
  reg                 io_in_c_bypass_regNext_11_2_is_stationary_26;
  reg        [15:0]   io_in_c_bypass_regNext_11_3_data_26;
  reg                 io_in_c_bypass_regNext_11_3_is_stationary_26;
  reg        [15:0]   io_in_c_bypass_regNext_12_0_data_26;
  reg                 io_in_c_bypass_regNext_12_0_is_stationary_26;
  reg        [15:0]   io_in_c_bypass_regNext_12_1_data_26;
  reg                 io_in_c_bypass_regNext_12_1_is_stationary_26;
  reg        [15:0]   io_in_c_bypass_regNext_12_2_data_26;
  reg                 io_in_c_bypass_regNext_12_2_is_stationary_26;
  reg        [15:0]   io_in_c_bypass_regNext_12_3_data_26;
  reg                 io_in_c_bypass_regNext_12_3_is_stationary_26;
  reg        [15:0]   io_in_c_bypass_regNext_13_0_data_26;
  reg                 io_in_c_bypass_regNext_13_0_is_stationary_26;
  reg        [15:0]   io_in_c_bypass_regNext_13_1_data_26;
  reg                 io_in_c_bypass_regNext_13_1_is_stationary_26;
  reg        [15:0]   io_in_c_bypass_regNext_13_2_data_26;
  reg                 io_in_c_bypass_regNext_13_2_is_stationary_26;
  reg        [15:0]   io_in_c_bypass_regNext_13_3_data_26;
  reg                 io_in_c_bypass_regNext_13_3_is_stationary_26;
  reg        [15:0]   io_in_c_bypass_regNext_14_0_data_26;
  reg                 io_in_c_bypass_regNext_14_0_is_stationary_26;
  reg        [15:0]   io_in_c_bypass_regNext_14_1_data_26;
  reg                 io_in_c_bypass_regNext_14_1_is_stationary_26;
  reg        [15:0]   io_in_c_bypass_regNext_14_2_data_26;
  reg                 io_in_c_bypass_regNext_14_2_is_stationary_26;
  reg        [15:0]   io_in_c_bypass_regNext_14_3_data_26;
  reg                 io_in_c_bypass_regNext_14_3_is_stationary_26;
  reg        [15:0]   io_in_c_bypass_regNext_15_0_data_26;
  reg                 io_in_c_bypass_regNext_15_0_is_stationary_26;
  reg        [15:0]   io_in_c_bypass_regNext_15_1_data_26;
  reg                 io_in_c_bypass_regNext_15_1_is_stationary_26;
  reg        [15:0]   io_in_c_bypass_regNext_15_2_data_26;
  reg                 io_in_c_bypass_regNext_15_2_is_stationary_26;
  reg        [15:0]   io_in_c_bypass_regNext_15_3_data_26;
  reg                 io_in_c_bypass_regNext_15_3_is_stationary_26;
  reg        [15:0]   io_in_c_bypass_regNext_16_0_data_26;
  reg                 io_in_c_bypass_regNext_16_0_is_stationary_26;
  reg        [15:0]   io_in_c_bypass_regNext_16_1_data_26;
  reg                 io_in_c_bypass_regNext_16_1_is_stationary_26;
  reg        [15:0]   io_in_c_bypass_regNext_16_2_data_26;
  reg                 io_in_c_bypass_regNext_16_2_is_stationary_26;
  reg        [15:0]   io_in_c_bypass_regNext_16_3_data_26;
  reg                 io_in_c_bypass_regNext_16_3_is_stationary_26;
  reg        [15:0]   io_in_c_bypass_regNext_17_0_data_26;
  reg                 io_in_c_bypass_regNext_17_0_is_stationary_26;
  reg        [15:0]   io_in_c_bypass_regNext_17_1_data_26;
  reg                 io_in_c_bypass_regNext_17_1_is_stationary_26;
  reg        [15:0]   io_in_c_bypass_regNext_17_2_data_26;
  reg                 io_in_c_bypass_regNext_17_2_is_stationary_26;
  reg        [15:0]   io_in_c_bypass_regNext_17_3_data_26;
  reg                 io_in_c_bypass_regNext_17_3_is_stationary_26;
  reg        [15:0]   io_in_c_bypass_regNext_18_0_data_26;
  reg                 io_in_c_bypass_regNext_18_0_is_stationary_26;
  reg        [15:0]   io_in_c_bypass_regNext_18_1_data_26;
  reg                 io_in_c_bypass_regNext_18_1_is_stationary_26;
  reg        [15:0]   io_in_c_bypass_regNext_18_2_data_26;
  reg                 io_in_c_bypass_regNext_18_2_is_stationary_26;
  reg        [15:0]   io_in_c_bypass_regNext_18_3_data_26;
  reg                 io_in_c_bypass_regNext_18_3_is_stationary_26;
  reg        [15:0]   io_in_c_bypass_regNext_19_0_data_26;
  reg                 io_in_c_bypass_regNext_19_0_is_stationary_26;
  reg        [15:0]   io_in_c_bypass_regNext_19_1_data_26;
  reg                 io_in_c_bypass_regNext_19_1_is_stationary_26;
  reg        [15:0]   io_in_c_bypass_regNext_19_2_data_26;
  reg                 io_in_c_bypass_regNext_19_2_is_stationary_26;
  reg        [15:0]   io_in_c_bypass_regNext_19_3_data_26;
  reg                 io_in_c_bypass_regNext_19_3_is_stationary_26;
  reg        [15:0]   io_in_c_bypass_regNext_20_0_data_26;
  reg                 io_in_c_bypass_regNext_20_0_is_stationary_26;
  reg        [15:0]   io_in_c_bypass_regNext_20_1_data_26;
  reg                 io_in_c_bypass_regNext_20_1_is_stationary_26;
  reg        [15:0]   io_in_c_bypass_regNext_20_2_data_26;
  reg                 io_in_c_bypass_regNext_20_2_is_stationary_26;
  reg        [15:0]   io_in_c_bypass_regNext_20_3_data_26;
  reg                 io_in_c_bypass_regNext_20_3_is_stationary_26;
  reg        [15:0]   io_in_c_bypass_regNext_21_0_data_26;
  reg                 io_in_c_bypass_regNext_21_0_is_stationary_26;
  reg        [15:0]   io_in_c_bypass_regNext_21_1_data_26;
  reg                 io_in_c_bypass_regNext_21_1_is_stationary_26;
  reg        [15:0]   io_in_c_bypass_regNext_21_2_data_26;
  reg                 io_in_c_bypass_regNext_21_2_is_stationary_26;
  reg        [15:0]   io_in_c_bypass_regNext_21_3_data_26;
  reg                 io_in_c_bypass_regNext_21_3_is_stationary_26;
  reg        [15:0]   io_in_c_bypass_regNext_22_0_data_26;
  reg                 io_in_c_bypass_regNext_22_0_is_stationary_26;
  reg        [15:0]   io_in_c_bypass_regNext_22_1_data_26;
  reg                 io_in_c_bypass_regNext_22_1_is_stationary_26;
  reg        [15:0]   io_in_c_bypass_regNext_22_2_data_26;
  reg                 io_in_c_bypass_regNext_22_2_is_stationary_26;
  reg        [15:0]   io_in_c_bypass_regNext_22_3_data_26;
  reg                 io_in_c_bypass_regNext_22_3_is_stationary_26;
  reg        [15:0]   io_in_c_bypass_regNext_23_0_data_26;
  reg                 io_in_c_bypass_regNext_23_0_is_stationary_26;
  reg        [15:0]   io_in_c_bypass_regNext_23_1_data_26;
  reg                 io_in_c_bypass_regNext_23_1_is_stationary_26;
  reg        [15:0]   io_in_c_bypass_regNext_23_2_data_26;
  reg                 io_in_c_bypass_regNext_23_2_is_stationary_26;
  reg        [15:0]   io_in_c_bypass_regNext_23_3_data_26;
  reg                 io_in_c_bypass_regNext_23_3_is_stationary_26;
  reg        [15:0]   io_in_c_bypass_regNext_24_0_data_26;
  reg                 io_in_c_bypass_regNext_24_0_is_stationary_26;
  reg        [15:0]   io_in_c_bypass_regNext_24_1_data_26;
  reg                 io_in_c_bypass_regNext_24_1_is_stationary_26;
  reg        [15:0]   io_in_c_bypass_regNext_24_2_data_26;
  reg                 io_in_c_bypass_regNext_24_2_is_stationary_26;
  reg        [15:0]   io_in_c_bypass_regNext_24_3_data_26;
  reg                 io_in_c_bypass_regNext_24_3_is_stationary_26;
  reg        [15:0]   io_in_c_bypass_regNext_25_0_data_26;
  reg                 io_in_c_bypass_regNext_25_0_is_stationary_26;
  reg        [15:0]   io_in_c_bypass_regNext_25_1_data_26;
  reg                 io_in_c_bypass_regNext_25_1_is_stationary_26;
  reg        [15:0]   io_in_c_bypass_regNext_25_2_data_26;
  reg                 io_in_c_bypass_regNext_25_2_is_stationary_26;
  reg        [15:0]   io_in_c_bypass_regNext_25_3_data_26;
  reg                 io_in_c_bypass_regNext_25_3_is_stationary_26;
  reg        [15:0]   io_in_c_bypass_regNext_26_0_data_26;
  reg                 io_in_c_bypass_regNext_26_0_is_stationary_26;
  reg        [15:0]   io_in_c_bypass_regNext_26_1_data_26;
  reg                 io_in_c_bypass_regNext_26_1_is_stationary_26;
  reg        [15:0]   io_in_c_bypass_regNext_26_2_data_26;
  reg                 io_in_c_bypass_regNext_26_2_is_stationary_26;
  reg        [15:0]   io_in_c_bypass_regNext_26_3_data_26;
  reg                 io_in_c_bypass_regNext_26_3_is_stationary_26;
  reg        [15:0]   io_in_c_bypass_regNext_27_0_data_26;
  reg                 io_in_c_bypass_regNext_27_0_is_stationary_26;
  reg        [15:0]   io_in_c_bypass_regNext_27_1_data_26;
  reg                 io_in_c_bypass_regNext_27_1_is_stationary_26;
  reg        [15:0]   io_in_c_bypass_regNext_27_2_data_26;
  reg                 io_in_c_bypass_regNext_27_2_is_stationary_26;
  reg        [15:0]   io_in_c_bypass_regNext_27_3_data_26;
  reg                 io_in_c_bypass_regNext_27_3_is_stationary_26;
  reg        [15:0]   io_in_c_bypass_regNext_28_0_data_26;
  reg                 io_in_c_bypass_regNext_28_0_is_stationary_26;
  reg        [15:0]   io_in_c_bypass_regNext_28_1_data_26;
  reg                 io_in_c_bypass_regNext_28_1_is_stationary_26;
  reg        [15:0]   io_in_c_bypass_regNext_28_2_data_26;
  reg                 io_in_c_bypass_regNext_28_2_is_stationary_26;
  reg        [15:0]   io_in_c_bypass_regNext_28_3_data_26;
  reg                 io_in_c_bypass_regNext_28_3_is_stationary_26;
  reg        [15:0]   io_in_c_bypass_regNext_29_0_data_26;
  reg                 io_in_c_bypass_regNext_29_0_is_stationary_26;
  reg        [15:0]   io_in_c_bypass_regNext_29_1_data_26;
  reg                 io_in_c_bypass_regNext_29_1_is_stationary_26;
  reg        [15:0]   io_in_c_bypass_regNext_29_2_data_26;
  reg                 io_in_c_bypass_regNext_29_2_is_stationary_26;
  reg        [15:0]   io_in_c_bypass_regNext_29_3_data_26;
  reg                 io_in_c_bypass_regNext_29_3_is_stationary_26;
  reg        [15:0]   io_in_c_bypass_regNext_30_0_data_26;
  reg                 io_in_c_bypass_regNext_30_0_is_stationary_26;
  reg        [15:0]   io_in_c_bypass_regNext_30_1_data_26;
  reg                 io_in_c_bypass_regNext_30_1_is_stationary_26;
  reg        [15:0]   io_in_c_bypass_regNext_30_2_data_26;
  reg                 io_in_c_bypass_regNext_30_2_is_stationary_26;
  reg        [15:0]   io_in_c_bypass_regNext_30_3_data_26;
  reg                 io_in_c_bypass_regNext_30_3_is_stationary_26;
  reg        [15:0]   io_in_c_bypass_regNext_31_0_data_26;
  reg                 io_in_c_bypass_regNext_31_0_is_stationary_26;
  reg        [15:0]   io_in_c_bypass_regNext_31_1_data_26;
  reg                 io_in_c_bypass_regNext_31_1_is_stationary_26;
  reg        [15:0]   io_in_c_bypass_regNext_31_2_data_26;
  reg                 io_in_c_bypass_regNext_31_2_is_stationary_26;
  reg        [15:0]   io_in_c_bypass_regNext_31_3_data_26;
  reg                 io_in_c_bypass_regNext_31_3_is_stationary_26;
  reg        [15:0]   io_in_c_bypass_regNext_0_0_data_27;
  reg                 io_in_c_bypass_regNext_0_0_is_stationary_27;
  reg        [15:0]   io_in_c_bypass_regNext_0_1_data_27;
  reg                 io_in_c_bypass_regNext_0_1_is_stationary_27;
  reg        [15:0]   io_in_c_bypass_regNext_0_2_data_27;
  reg                 io_in_c_bypass_regNext_0_2_is_stationary_27;
  reg        [15:0]   io_in_c_bypass_regNext_0_3_data_27;
  reg                 io_in_c_bypass_regNext_0_3_is_stationary_27;
  reg        [15:0]   io_in_c_bypass_regNext_1_0_data_27;
  reg                 io_in_c_bypass_regNext_1_0_is_stationary_27;
  reg        [15:0]   io_in_c_bypass_regNext_1_1_data_27;
  reg                 io_in_c_bypass_regNext_1_1_is_stationary_27;
  reg        [15:0]   io_in_c_bypass_regNext_1_2_data_27;
  reg                 io_in_c_bypass_regNext_1_2_is_stationary_27;
  reg        [15:0]   io_in_c_bypass_regNext_1_3_data_27;
  reg                 io_in_c_bypass_regNext_1_3_is_stationary_27;
  reg        [15:0]   io_in_c_bypass_regNext_2_0_data_27;
  reg                 io_in_c_bypass_regNext_2_0_is_stationary_27;
  reg        [15:0]   io_in_c_bypass_regNext_2_1_data_27;
  reg                 io_in_c_bypass_regNext_2_1_is_stationary_27;
  reg        [15:0]   io_in_c_bypass_regNext_2_2_data_27;
  reg                 io_in_c_bypass_regNext_2_2_is_stationary_27;
  reg        [15:0]   io_in_c_bypass_regNext_2_3_data_27;
  reg                 io_in_c_bypass_regNext_2_3_is_stationary_27;
  reg        [15:0]   io_in_c_bypass_regNext_3_0_data_27;
  reg                 io_in_c_bypass_regNext_3_0_is_stationary_27;
  reg        [15:0]   io_in_c_bypass_regNext_3_1_data_27;
  reg                 io_in_c_bypass_regNext_3_1_is_stationary_27;
  reg        [15:0]   io_in_c_bypass_regNext_3_2_data_27;
  reg                 io_in_c_bypass_regNext_3_2_is_stationary_27;
  reg        [15:0]   io_in_c_bypass_regNext_3_3_data_27;
  reg                 io_in_c_bypass_regNext_3_3_is_stationary_27;
  reg        [15:0]   io_in_c_bypass_regNext_4_0_data_27;
  reg                 io_in_c_bypass_regNext_4_0_is_stationary_27;
  reg        [15:0]   io_in_c_bypass_regNext_4_1_data_27;
  reg                 io_in_c_bypass_regNext_4_1_is_stationary_27;
  reg        [15:0]   io_in_c_bypass_regNext_4_2_data_27;
  reg                 io_in_c_bypass_regNext_4_2_is_stationary_27;
  reg        [15:0]   io_in_c_bypass_regNext_4_3_data_27;
  reg                 io_in_c_bypass_regNext_4_3_is_stationary_27;
  reg        [15:0]   io_in_c_bypass_regNext_5_0_data_27;
  reg                 io_in_c_bypass_regNext_5_0_is_stationary_27;
  reg        [15:0]   io_in_c_bypass_regNext_5_1_data_27;
  reg                 io_in_c_bypass_regNext_5_1_is_stationary_27;
  reg        [15:0]   io_in_c_bypass_regNext_5_2_data_27;
  reg                 io_in_c_bypass_regNext_5_2_is_stationary_27;
  reg        [15:0]   io_in_c_bypass_regNext_5_3_data_27;
  reg                 io_in_c_bypass_regNext_5_3_is_stationary_27;
  reg        [15:0]   io_in_c_bypass_regNext_6_0_data_27;
  reg                 io_in_c_bypass_regNext_6_0_is_stationary_27;
  reg        [15:0]   io_in_c_bypass_regNext_6_1_data_27;
  reg                 io_in_c_bypass_regNext_6_1_is_stationary_27;
  reg        [15:0]   io_in_c_bypass_regNext_6_2_data_27;
  reg                 io_in_c_bypass_regNext_6_2_is_stationary_27;
  reg        [15:0]   io_in_c_bypass_regNext_6_3_data_27;
  reg                 io_in_c_bypass_regNext_6_3_is_stationary_27;
  reg        [15:0]   io_in_c_bypass_regNext_7_0_data_27;
  reg                 io_in_c_bypass_regNext_7_0_is_stationary_27;
  reg        [15:0]   io_in_c_bypass_regNext_7_1_data_27;
  reg                 io_in_c_bypass_regNext_7_1_is_stationary_27;
  reg        [15:0]   io_in_c_bypass_regNext_7_2_data_27;
  reg                 io_in_c_bypass_regNext_7_2_is_stationary_27;
  reg        [15:0]   io_in_c_bypass_regNext_7_3_data_27;
  reg                 io_in_c_bypass_regNext_7_3_is_stationary_27;
  reg        [15:0]   io_in_c_bypass_regNext_8_0_data_27;
  reg                 io_in_c_bypass_regNext_8_0_is_stationary_27;
  reg        [15:0]   io_in_c_bypass_regNext_8_1_data_27;
  reg                 io_in_c_bypass_regNext_8_1_is_stationary_27;
  reg        [15:0]   io_in_c_bypass_regNext_8_2_data_27;
  reg                 io_in_c_bypass_regNext_8_2_is_stationary_27;
  reg        [15:0]   io_in_c_bypass_regNext_8_3_data_27;
  reg                 io_in_c_bypass_regNext_8_3_is_stationary_27;
  reg        [15:0]   io_in_c_bypass_regNext_9_0_data_27;
  reg                 io_in_c_bypass_regNext_9_0_is_stationary_27;
  reg        [15:0]   io_in_c_bypass_regNext_9_1_data_27;
  reg                 io_in_c_bypass_regNext_9_1_is_stationary_27;
  reg        [15:0]   io_in_c_bypass_regNext_9_2_data_27;
  reg                 io_in_c_bypass_regNext_9_2_is_stationary_27;
  reg        [15:0]   io_in_c_bypass_regNext_9_3_data_27;
  reg                 io_in_c_bypass_regNext_9_3_is_stationary_27;
  reg        [15:0]   io_in_c_bypass_regNext_10_0_data_27;
  reg                 io_in_c_bypass_regNext_10_0_is_stationary_27;
  reg        [15:0]   io_in_c_bypass_regNext_10_1_data_27;
  reg                 io_in_c_bypass_regNext_10_1_is_stationary_27;
  reg        [15:0]   io_in_c_bypass_regNext_10_2_data_27;
  reg                 io_in_c_bypass_regNext_10_2_is_stationary_27;
  reg        [15:0]   io_in_c_bypass_regNext_10_3_data_27;
  reg                 io_in_c_bypass_regNext_10_3_is_stationary_27;
  reg        [15:0]   io_in_c_bypass_regNext_11_0_data_27;
  reg                 io_in_c_bypass_regNext_11_0_is_stationary_27;
  reg        [15:0]   io_in_c_bypass_regNext_11_1_data_27;
  reg                 io_in_c_bypass_regNext_11_1_is_stationary_27;
  reg        [15:0]   io_in_c_bypass_regNext_11_2_data_27;
  reg                 io_in_c_bypass_regNext_11_2_is_stationary_27;
  reg        [15:0]   io_in_c_bypass_regNext_11_3_data_27;
  reg                 io_in_c_bypass_regNext_11_3_is_stationary_27;
  reg        [15:0]   io_in_c_bypass_regNext_12_0_data_27;
  reg                 io_in_c_bypass_regNext_12_0_is_stationary_27;
  reg        [15:0]   io_in_c_bypass_regNext_12_1_data_27;
  reg                 io_in_c_bypass_regNext_12_1_is_stationary_27;
  reg        [15:0]   io_in_c_bypass_regNext_12_2_data_27;
  reg                 io_in_c_bypass_regNext_12_2_is_stationary_27;
  reg        [15:0]   io_in_c_bypass_regNext_12_3_data_27;
  reg                 io_in_c_bypass_regNext_12_3_is_stationary_27;
  reg        [15:0]   io_in_c_bypass_regNext_13_0_data_27;
  reg                 io_in_c_bypass_regNext_13_0_is_stationary_27;
  reg        [15:0]   io_in_c_bypass_regNext_13_1_data_27;
  reg                 io_in_c_bypass_regNext_13_1_is_stationary_27;
  reg        [15:0]   io_in_c_bypass_regNext_13_2_data_27;
  reg                 io_in_c_bypass_regNext_13_2_is_stationary_27;
  reg        [15:0]   io_in_c_bypass_regNext_13_3_data_27;
  reg                 io_in_c_bypass_regNext_13_3_is_stationary_27;
  reg        [15:0]   io_in_c_bypass_regNext_14_0_data_27;
  reg                 io_in_c_bypass_regNext_14_0_is_stationary_27;
  reg        [15:0]   io_in_c_bypass_regNext_14_1_data_27;
  reg                 io_in_c_bypass_regNext_14_1_is_stationary_27;
  reg        [15:0]   io_in_c_bypass_regNext_14_2_data_27;
  reg                 io_in_c_bypass_regNext_14_2_is_stationary_27;
  reg        [15:0]   io_in_c_bypass_regNext_14_3_data_27;
  reg                 io_in_c_bypass_regNext_14_3_is_stationary_27;
  reg        [15:0]   io_in_c_bypass_regNext_15_0_data_27;
  reg                 io_in_c_bypass_regNext_15_0_is_stationary_27;
  reg        [15:0]   io_in_c_bypass_regNext_15_1_data_27;
  reg                 io_in_c_bypass_regNext_15_1_is_stationary_27;
  reg        [15:0]   io_in_c_bypass_regNext_15_2_data_27;
  reg                 io_in_c_bypass_regNext_15_2_is_stationary_27;
  reg        [15:0]   io_in_c_bypass_regNext_15_3_data_27;
  reg                 io_in_c_bypass_regNext_15_3_is_stationary_27;
  reg        [15:0]   io_in_c_bypass_regNext_16_0_data_27;
  reg                 io_in_c_bypass_regNext_16_0_is_stationary_27;
  reg        [15:0]   io_in_c_bypass_regNext_16_1_data_27;
  reg                 io_in_c_bypass_regNext_16_1_is_stationary_27;
  reg        [15:0]   io_in_c_bypass_regNext_16_2_data_27;
  reg                 io_in_c_bypass_regNext_16_2_is_stationary_27;
  reg        [15:0]   io_in_c_bypass_regNext_16_3_data_27;
  reg                 io_in_c_bypass_regNext_16_3_is_stationary_27;
  reg        [15:0]   io_in_c_bypass_regNext_17_0_data_27;
  reg                 io_in_c_bypass_regNext_17_0_is_stationary_27;
  reg        [15:0]   io_in_c_bypass_regNext_17_1_data_27;
  reg                 io_in_c_bypass_regNext_17_1_is_stationary_27;
  reg        [15:0]   io_in_c_bypass_regNext_17_2_data_27;
  reg                 io_in_c_bypass_regNext_17_2_is_stationary_27;
  reg        [15:0]   io_in_c_bypass_regNext_17_3_data_27;
  reg                 io_in_c_bypass_regNext_17_3_is_stationary_27;
  reg        [15:0]   io_in_c_bypass_regNext_18_0_data_27;
  reg                 io_in_c_bypass_regNext_18_0_is_stationary_27;
  reg        [15:0]   io_in_c_bypass_regNext_18_1_data_27;
  reg                 io_in_c_bypass_regNext_18_1_is_stationary_27;
  reg        [15:0]   io_in_c_bypass_regNext_18_2_data_27;
  reg                 io_in_c_bypass_regNext_18_2_is_stationary_27;
  reg        [15:0]   io_in_c_bypass_regNext_18_3_data_27;
  reg                 io_in_c_bypass_regNext_18_3_is_stationary_27;
  reg        [15:0]   io_in_c_bypass_regNext_19_0_data_27;
  reg                 io_in_c_bypass_regNext_19_0_is_stationary_27;
  reg        [15:0]   io_in_c_bypass_regNext_19_1_data_27;
  reg                 io_in_c_bypass_regNext_19_1_is_stationary_27;
  reg        [15:0]   io_in_c_bypass_regNext_19_2_data_27;
  reg                 io_in_c_bypass_regNext_19_2_is_stationary_27;
  reg        [15:0]   io_in_c_bypass_regNext_19_3_data_27;
  reg                 io_in_c_bypass_regNext_19_3_is_stationary_27;
  reg        [15:0]   io_in_c_bypass_regNext_20_0_data_27;
  reg                 io_in_c_bypass_regNext_20_0_is_stationary_27;
  reg        [15:0]   io_in_c_bypass_regNext_20_1_data_27;
  reg                 io_in_c_bypass_regNext_20_1_is_stationary_27;
  reg        [15:0]   io_in_c_bypass_regNext_20_2_data_27;
  reg                 io_in_c_bypass_regNext_20_2_is_stationary_27;
  reg        [15:0]   io_in_c_bypass_regNext_20_3_data_27;
  reg                 io_in_c_bypass_regNext_20_3_is_stationary_27;
  reg        [15:0]   io_in_c_bypass_regNext_21_0_data_27;
  reg                 io_in_c_bypass_regNext_21_0_is_stationary_27;
  reg        [15:0]   io_in_c_bypass_regNext_21_1_data_27;
  reg                 io_in_c_bypass_regNext_21_1_is_stationary_27;
  reg        [15:0]   io_in_c_bypass_regNext_21_2_data_27;
  reg                 io_in_c_bypass_regNext_21_2_is_stationary_27;
  reg        [15:0]   io_in_c_bypass_regNext_21_3_data_27;
  reg                 io_in_c_bypass_regNext_21_3_is_stationary_27;
  reg        [15:0]   io_in_c_bypass_regNext_22_0_data_27;
  reg                 io_in_c_bypass_regNext_22_0_is_stationary_27;
  reg        [15:0]   io_in_c_bypass_regNext_22_1_data_27;
  reg                 io_in_c_bypass_regNext_22_1_is_stationary_27;
  reg        [15:0]   io_in_c_bypass_regNext_22_2_data_27;
  reg                 io_in_c_bypass_regNext_22_2_is_stationary_27;
  reg        [15:0]   io_in_c_bypass_regNext_22_3_data_27;
  reg                 io_in_c_bypass_regNext_22_3_is_stationary_27;
  reg        [15:0]   io_in_c_bypass_regNext_23_0_data_27;
  reg                 io_in_c_bypass_regNext_23_0_is_stationary_27;
  reg        [15:0]   io_in_c_bypass_regNext_23_1_data_27;
  reg                 io_in_c_bypass_regNext_23_1_is_stationary_27;
  reg        [15:0]   io_in_c_bypass_regNext_23_2_data_27;
  reg                 io_in_c_bypass_regNext_23_2_is_stationary_27;
  reg        [15:0]   io_in_c_bypass_regNext_23_3_data_27;
  reg                 io_in_c_bypass_regNext_23_3_is_stationary_27;
  reg        [15:0]   io_in_c_bypass_regNext_24_0_data_27;
  reg                 io_in_c_bypass_regNext_24_0_is_stationary_27;
  reg        [15:0]   io_in_c_bypass_regNext_24_1_data_27;
  reg                 io_in_c_bypass_regNext_24_1_is_stationary_27;
  reg        [15:0]   io_in_c_bypass_regNext_24_2_data_27;
  reg                 io_in_c_bypass_regNext_24_2_is_stationary_27;
  reg        [15:0]   io_in_c_bypass_regNext_24_3_data_27;
  reg                 io_in_c_bypass_regNext_24_3_is_stationary_27;
  reg        [15:0]   io_in_c_bypass_regNext_25_0_data_27;
  reg                 io_in_c_bypass_regNext_25_0_is_stationary_27;
  reg        [15:0]   io_in_c_bypass_regNext_25_1_data_27;
  reg                 io_in_c_bypass_regNext_25_1_is_stationary_27;
  reg        [15:0]   io_in_c_bypass_regNext_25_2_data_27;
  reg                 io_in_c_bypass_regNext_25_2_is_stationary_27;
  reg        [15:0]   io_in_c_bypass_regNext_25_3_data_27;
  reg                 io_in_c_bypass_regNext_25_3_is_stationary_27;
  reg        [15:0]   io_in_c_bypass_regNext_26_0_data_27;
  reg                 io_in_c_bypass_regNext_26_0_is_stationary_27;
  reg        [15:0]   io_in_c_bypass_regNext_26_1_data_27;
  reg                 io_in_c_bypass_regNext_26_1_is_stationary_27;
  reg        [15:0]   io_in_c_bypass_regNext_26_2_data_27;
  reg                 io_in_c_bypass_regNext_26_2_is_stationary_27;
  reg        [15:0]   io_in_c_bypass_regNext_26_3_data_27;
  reg                 io_in_c_bypass_regNext_26_3_is_stationary_27;
  reg        [15:0]   io_in_c_bypass_regNext_27_0_data_27;
  reg                 io_in_c_bypass_regNext_27_0_is_stationary_27;
  reg        [15:0]   io_in_c_bypass_regNext_27_1_data_27;
  reg                 io_in_c_bypass_regNext_27_1_is_stationary_27;
  reg        [15:0]   io_in_c_bypass_regNext_27_2_data_27;
  reg                 io_in_c_bypass_regNext_27_2_is_stationary_27;
  reg        [15:0]   io_in_c_bypass_regNext_27_3_data_27;
  reg                 io_in_c_bypass_regNext_27_3_is_stationary_27;
  reg        [15:0]   io_in_c_bypass_regNext_28_0_data_27;
  reg                 io_in_c_bypass_regNext_28_0_is_stationary_27;
  reg        [15:0]   io_in_c_bypass_regNext_28_1_data_27;
  reg                 io_in_c_bypass_regNext_28_1_is_stationary_27;
  reg        [15:0]   io_in_c_bypass_regNext_28_2_data_27;
  reg                 io_in_c_bypass_regNext_28_2_is_stationary_27;
  reg        [15:0]   io_in_c_bypass_regNext_28_3_data_27;
  reg                 io_in_c_bypass_regNext_28_3_is_stationary_27;
  reg        [15:0]   io_in_c_bypass_regNext_29_0_data_27;
  reg                 io_in_c_bypass_regNext_29_0_is_stationary_27;
  reg        [15:0]   io_in_c_bypass_regNext_29_1_data_27;
  reg                 io_in_c_bypass_regNext_29_1_is_stationary_27;
  reg        [15:0]   io_in_c_bypass_regNext_29_2_data_27;
  reg                 io_in_c_bypass_regNext_29_2_is_stationary_27;
  reg        [15:0]   io_in_c_bypass_regNext_29_3_data_27;
  reg                 io_in_c_bypass_regNext_29_3_is_stationary_27;
  reg        [15:0]   io_in_c_bypass_regNext_30_0_data_27;
  reg                 io_in_c_bypass_regNext_30_0_is_stationary_27;
  reg        [15:0]   io_in_c_bypass_regNext_30_1_data_27;
  reg                 io_in_c_bypass_regNext_30_1_is_stationary_27;
  reg        [15:0]   io_in_c_bypass_regNext_30_2_data_27;
  reg                 io_in_c_bypass_regNext_30_2_is_stationary_27;
  reg        [15:0]   io_in_c_bypass_regNext_30_3_data_27;
  reg                 io_in_c_bypass_regNext_30_3_is_stationary_27;
  reg        [15:0]   io_in_c_bypass_regNext_31_0_data_27;
  reg                 io_in_c_bypass_regNext_31_0_is_stationary_27;
  reg        [15:0]   io_in_c_bypass_regNext_31_1_data_27;
  reg                 io_in_c_bypass_regNext_31_1_is_stationary_27;
  reg        [15:0]   io_in_c_bypass_regNext_31_2_data_27;
  reg                 io_in_c_bypass_regNext_31_2_is_stationary_27;
  reg        [15:0]   io_in_c_bypass_regNext_31_3_data_27;
  reg                 io_in_c_bypass_regNext_31_3_is_stationary_27;
  reg        [15:0]   io_in_c_bypass_regNext_0_0_data_28;
  reg                 io_in_c_bypass_regNext_0_0_is_stationary_28;
  reg        [15:0]   io_in_c_bypass_regNext_0_1_data_28;
  reg                 io_in_c_bypass_regNext_0_1_is_stationary_28;
  reg        [15:0]   io_in_c_bypass_regNext_0_2_data_28;
  reg                 io_in_c_bypass_regNext_0_2_is_stationary_28;
  reg        [15:0]   io_in_c_bypass_regNext_0_3_data_28;
  reg                 io_in_c_bypass_regNext_0_3_is_stationary_28;
  reg        [15:0]   io_in_c_bypass_regNext_1_0_data_28;
  reg                 io_in_c_bypass_regNext_1_0_is_stationary_28;
  reg        [15:0]   io_in_c_bypass_regNext_1_1_data_28;
  reg                 io_in_c_bypass_regNext_1_1_is_stationary_28;
  reg        [15:0]   io_in_c_bypass_regNext_1_2_data_28;
  reg                 io_in_c_bypass_regNext_1_2_is_stationary_28;
  reg        [15:0]   io_in_c_bypass_regNext_1_3_data_28;
  reg                 io_in_c_bypass_regNext_1_3_is_stationary_28;
  reg        [15:0]   io_in_c_bypass_regNext_2_0_data_28;
  reg                 io_in_c_bypass_regNext_2_0_is_stationary_28;
  reg        [15:0]   io_in_c_bypass_regNext_2_1_data_28;
  reg                 io_in_c_bypass_regNext_2_1_is_stationary_28;
  reg        [15:0]   io_in_c_bypass_regNext_2_2_data_28;
  reg                 io_in_c_bypass_regNext_2_2_is_stationary_28;
  reg        [15:0]   io_in_c_bypass_regNext_2_3_data_28;
  reg                 io_in_c_bypass_regNext_2_3_is_stationary_28;
  reg        [15:0]   io_in_c_bypass_regNext_3_0_data_28;
  reg                 io_in_c_bypass_regNext_3_0_is_stationary_28;
  reg        [15:0]   io_in_c_bypass_regNext_3_1_data_28;
  reg                 io_in_c_bypass_regNext_3_1_is_stationary_28;
  reg        [15:0]   io_in_c_bypass_regNext_3_2_data_28;
  reg                 io_in_c_bypass_regNext_3_2_is_stationary_28;
  reg        [15:0]   io_in_c_bypass_regNext_3_3_data_28;
  reg                 io_in_c_bypass_regNext_3_3_is_stationary_28;
  reg        [15:0]   io_in_c_bypass_regNext_4_0_data_28;
  reg                 io_in_c_bypass_regNext_4_0_is_stationary_28;
  reg        [15:0]   io_in_c_bypass_regNext_4_1_data_28;
  reg                 io_in_c_bypass_regNext_4_1_is_stationary_28;
  reg        [15:0]   io_in_c_bypass_regNext_4_2_data_28;
  reg                 io_in_c_bypass_regNext_4_2_is_stationary_28;
  reg        [15:0]   io_in_c_bypass_regNext_4_3_data_28;
  reg                 io_in_c_bypass_regNext_4_3_is_stationary_28;
  reg        [15:0]   io_in_c_bypass_regNext_5_0_data_28;
  reg                 io_in_c_bypass_regNext_5_0_is_stationary_28;
  reg        [15:0]   io_in_c_bypass_regNext_5_1_data_28;
  reg                 io_in_c_bypass_regNext_5_1_is_stationary_28;
  reg        [15:0]   io_in_c_bypass_regNext_5_2_data_28;
  reg                 io_in_c_bypass_regNext_5_2_is_stationary_28;
  reg        [15:0]   io_in_c_bypass_regNext_5_3_data_28;
  reg                 io_in_c_bypass_regNext_5_3_is_stationary_28;
  reg        [15:0]   io_in_c_bypass_regNext_6_0_data_28;
  reg                 io_in_c_bypass_regNext_6_0_is_stationary_28;
  reg        [15:0]   io_in_c_bypass_regNext_6_1_data_28;
  reg                 io_in_c_bypass_regNext_6_1_is_stationary_28;
  reg        [15:0]   io_in_c_bypass_regNext_6_2_data_28;
  reg                 io_in_c_bypass_regNext_6_2_is_stationary_28;
  reg        [15:0]   io_in_c_bypass_regNext_6_3_data_28;
  reg                 io_in_c_bypass_regNext_6_3_is_stationary_28;
  reg        [15:0]   io_in_c_bypass_regNext_7_0_data_28;
  reg                 io_in_c_bypass_regNext_7_0_is_stationary_28;
  reg        [15:0]   io_in_c_bypass_regNext_7_1_data_28;
  reg                 io_in_c_bypass_regNext_7_1_is_stationary_28;
  reg        [15:0]   io_in_c_bypass_regNext_7_2_data_28;
  reg                 io_in_c_bypass_regNext_7_2_is_stationary_28;
  reg        [15:0]   io_in_c_bypass_regNext_7_3_data_28;
  reg                 io_in_c_bypass_regNext_7_3_is_stationary_28;
  reg        [15:0]   io_in_c_bypass_regNext_8_0_data_28;
  reg                 io_in_c_bypass_regNext_8_0_is_stationary_28;
  reg        [15:0]   io_in_c_bypass_regNext_8_1_data_28;
  reg                 io_in_c_bypass_regNext_8_1_is_stationary_28;
  reg        [15:0]   io_in_c_bypass_regNext_8_2_data_28;
  reg                 io_in_c_bypass_regNext_8_2_is_stationary_28;
  reg        [15:0]   io_in_c_bypass_regNext_8_3_data_28;
  reg                 io_in_c_bypass_regNext_8_3_is_stationary_28;
  reg        [15:0]   io_in_c_bypass_regNext_9_0_data_28;
  reg                 io_in_c_bypass_regNext_9_0_is_stationary_28;
  reg        [15:0]   io_in_c_bypass_regNext_9_1_data_28;
  reg                 io_in_c_bypass_regNext_9_1_is_stationary_28;
  reg        [15:0]   io_in_c_bypass_regNext_9_2_data_28;
  reg                 io_in_c_bypass_regNext_9_2_is_stationary_28;
  reg        [15:0]   io_in_c_bypass_regNext_9_3_data_28;
  reg                 io_in_c_bypass_regNext_9_3_is_stationary_28;
  reg        [15:0]   io_in_c_bypass_regNext_10_0_data_28;
  reg                 io_in_c_bypass_regNext_10_0_is_stationary_28;
  reg        [15:0]   io_in_c_bypass_regNext_10_1_data_28;
  reg                 io_in_c_bypass_regNext_10_1_is_stationary_28;
  reg        [15:0]   io_in_c_bypass_regNext_10_2_data_28;
  reg                 io_in_c_bypass_regNext_10_2_is_stationary_28;
  reg        [15:0]   io_in_c_bypass_regNext_10_3_data_28;
  reg                 io_in_c_bypass_regNext_10_3_is_stationary_28;
  reg        [15:0]   io_in_c_bypass_regNext_11_0_data_28;
  reg                 io_in_c_bypass_regNext_11_0_is_stationary_28;
  reg        [15:0]   io_in_c_bypass_regNext_11_1_data_28;
  reg                 io_in_c_bypass_regNext_11_1_is_stationary_28;
  reg        [15:0]   io_in_c_bypass_regNext_11_2_data_28;
  reg                 io_in_c_bypass_regNext_11_2_is_stationary_28;
  reg        [15:0]   io_in_c_bypass_regNext_11_3_data_28;
  reg                 io_in_c_bypass_regNext_11_3_is_stationary_28;
  reg        [15:0]   io_in_c_bypass_regNext_12_0_data_28;
  reg                 io_in_c_bypass_regNext_12_0_is_stationary_28;
  reg        [15:0]   io_in_c_bypass_regNext_12_1_data_28;
  reg                 io_in_c_bypass_regNext_12_1_is_stationary_28;
  reg        [15:0]   io_in_c_bypass_regNext_12_2_data_28;
  reg                 io_in_c_bypass_regNext_12_2_is_stationary_28;
  reg        [15:0]   io_in_c_bypass_regNext_12_3_data_28;
  reg                 io_in_c_bypass_regNext_12_3_is_stationary_28;
  reg        [15:0]   io_in_c_bypass_regNext_13_0_data_28;
  reg                 io_in_c_bypass_regNext_13_0_is_stationary_28;
  reg        [15:0]   io_in_c_bypass_regNext_13_1_data_28;
  reg                 io_in_c_bypass_regNext_13_1_is_stationary_28;
  reg        [15:0]   io_in_c_bypass_regNext_13_2_data_28;
  reg                 io_in_c_bypass_regNext_13_2_is_stationary_28;
  reg        [15:0]   io_in_c_bypass_regNext_13_3_data_28;
  reg                 io_in_c_bypass_regNext_13_3_is_stationary_28;
  reg        [15:0]   io_in_c_bypass_regNext_14_0_data_28;
  reg                 io_in_c_bypass_regNext_14_0_is_stationary_28;
  reg        [15:0]   io_in_c_bypass_regNext_14_1_data_28;
  reg                 io_in_c_bypass_regNext_14_1_is_stationary_28;
  reg        [15:0]   io_in_c_bypass_regNext_14_2_data_28;
  reg                 io_in_c_bypass_regNext_14_2_is_stationary_28;
  reg        [15:0]   io_in_c_bypass_regNext_14_3_data_28;
  reg                 io_in_c_bypass_regNext_14_3_is_stationary_28;
  reg        [15:0]   io_in_c_bypass_regNext_15_0_data_28;
  reg                 io_in_c_bypass_regNext_15_0_is_stationary_28;
  reg        [15:0]   io_in_c_bypass_regNext_15_1_data_28;
  reg                 io_in_c_bypass_regNext_15_1_is_stationary_28;
  reg        [15:0]   io_in_c_bypass_regNext_15_2_data_28;
  reg                 io_in_c_bypass_regNext_15_2_is_stationary_28;
  reg        [15:0]   io_in_c_bypass_regNext_15_3_data_28;
  reg                 io_in_c_bypass_regNext_15_3_is_stationary_28;
  reg        [15:0]   io_in_c_bypass_regNext_16_0_data_28;
  reg                 io_in_c_bypass_regNext_16_0_is_stationary_28;
  reg        [15:0]   io_in_c_bypass_regNext_16_1_data_28;
  reg                 io_in_c_bypass_regNext_16_1_is_stationary_28;
  reg        [15:0]   io_in_c_bypass_regNext_16_2_data_28;
  reg                 io_in_c_bypass_regNext_16_2_is_stationary_28;
  reg        [15:0]   io_in_c_bypass_regNext_16_3_data_28;
  reg                 io_in_c_bypass_regNext_16_3_is_stationary_28;
  reg        [15:0]   io_in_c_bypass_regNext_17_0_data_28;
  reg                 io_in_c_bypass_regNext_17_0_is_stationary_28;
  reg        [15:0]   io_in_c_bypass_regNext_17_1_data_28;
  reg                 io_in_c_bypass_regNext_17_1_is_stationary_28;
  reg        [15:0]   io_in_c_bypass_regNext_17_2_data_28;
  reg                 io_in_c_bypass_regNext_17_2_is_stationary_28;
  reg        [15:0]   io_in_c_bypass_regNext_17_3_data_28;
  reg                 io_in_c_bypass_regNext_17_3_is_stationary_28;
  reg        [15:0]   io_in_c_bypass_regNext_18_0_data_28;
  reg                 io_in_c_bypass_regNext_18_0_is_stationary_28;
  reg        [15:0]   io_in_c_bypass_regNext_18_1_data_28;
  reg                 io_in_c_bypass_regNext_18_1_is_stationary_28;
  reg        [15:0]   io_in_c_bypass_regNext_18_2_data_28;
  reg                 io_in_c_bypass_regNext_18_2_is_stationary_28;
  reg        [15:0]   io_in_c_bypass_regNext_18_3_data_28;
  reg                 io_in_c_bypass_regNext_18_3_is_stationary_28;
  reg        [15:0]   io_in_c_bypass_regNext_19_0_data_28;
  reg                 io_in_c_bypass_regNext_19_0_is_stationary_28;
  reg        [15:0]   io_in_c_bypass_regNext_19_1_data_28;
  reg                 io_in_c_bypass_regNext_19_1_is_stationary_28;
  reg        [15:0]   io_in_c_bypass_regNext_19_2_data_28;
  reg                 io_in_c_bypass_regNext_19_2_is_stationary_28;
  reg        [15:0]   io_in_c_bypass_regNext_19_3_data_28;
  reg                 io_in_c_bypass_regNext_19_3_is_stationary_28;
  reg        [15:0]   io_in_c_bypass_regNext_20_0_data_28;
  reg                 io_in_c_bypass_regNext_20_0_is_stationary_28;
  reg        [15:0]   io_in_c_bypass_regNext_20_1_data_28;
  reg                 io_in_c_bypass_regNext_20_1_is_stationary_28;
  reg        [15:0]   io_in_c_bypass_regNext_20_2_data_28;
  reg                 io_in_c_bypass_regNext_20_2_is_stationary_28;
  reg        [15:0]   io_in_c_bypass_regNext_20_3_data_28;
  reg                 io_in_c_bypass_regNext_20_3_is_stationary_28;
  reg        [15:0]   io_in_c_bypass_regNext_21_0_data_28;
  reg                 io_in_c_bypass_regNext_21_0_is_stationary_28;
  reg        [15:0]   io_in_c_bypass_regNext_21_1_data_28;
  reg                 io_in_c_bypass_regNext_21_1_is_stationary_28;
  reg        [15:0]   io_in_c_bypass_regNext_21_2_data_28;
  reg                 io_in_c_bypass_regNext_21_2_is_stationary_28;
  reg        [15:0]   io_in_c_bypass_regNext_21_3_data_28;
  reg                 io_in_c_bypass_regNext_21_3_is_stationary_28;
  reg        [15:0]   io_in_c_bypass_regNext_22_0_data_28;
  reg                 io_in_c_bypass_regNext_22_0_is_stationary_28;
  reg        [15:0]   io_in_c_bypass_regNext_22_1_data_28;
  reg                 io_in_c_bypass_regNext_22_1_is_stationary_28;
  reg        [15:0]   io_in_c_bypass_regNext_22_2_data_28;
  reg                 io_in_c_bypass_regNext_22_2_is_stationary_28;
  reg        [15:0]   io_in_c_bypass_regNext_22_3_data_28;
  reg                 io_in_c_bypass_regNext_22_3_is_stationary_28;
  reg        [15:0]   io_in_c_bypass_regNext_23_0_data_28;
  reg                 io_in_c_bypass_regNext_23_0_is_stationary_28;
  reg        [15:0]   io_in_c_bypass_regNext_23_1_data_28;
  reg                 io_in_c_bypass_regNext_23_1_is_stationary_28;
  reg        [15:0]   io_in_c_bypass_regNext_23_2_data_28;
  reg                 io_in_c_bypass_regNext_23_2_is_stationary_28;
  reg        [15:0]   io_in_c_bypass_regNext_23_3_data_28;
  reg                 io_in_c_bypass_regNext_23_3_is_stationary_28;
  reg        [15:0]   io_in_c_bypass_regNext_24_0_data_28;
  reg                 io_in_c_bypass_regNext_24_0_is_stationary_28;
  reg        [15:0]   io_in_c_bypass_regNext_24_1_data_28;
  reg                 io_in_c_bypass_regNext_24_1_is_stationary_28;
  reg        [15:0]   io_in_c_bypass_regNext_24_2_data_28;
  reg                 io_in_c_bypass_regNext_24_2_is_stationary_28;
  reg        [15:0]   io_in_c_bypass_regNext_24_3_data_28;
  reg                 io_in_c_bypass_regNext_24_3_is_stationary_28;
  reg        [15:0]   io_in_c_bypass_regNext_25_0_data_28;
  reg                 io_in_c_bypass_regNext_25_0_is_stationary_28;
  reg        [15:0]   io_in_c_bypass_regNext_25_1_data_28;
  reg                 io_in_c_bypass_regNext_25_1_is_stationary_28;
  reg        [15:0]   io_in_c_bypass_regNext_25_2_data_28;
  reg                 io_in_c_bypass_regNext_25_2_is_stationary_28;
  reg        [15:0]   io_in_c_bypass_regNext_25_3_data_28;
  reg                 io_in_c_bypass_regNext_25_3_is_stationary_28;
  reg        [15:0]   io_in_c_bypass_regNext_26_0_data_28;
  reg                 io_in_c_bypass_regNext_26_0_is_stationary_28;
  reg        [15:0]   io_in_c_bypass_regNext_26_1_data_28;
  reg                 io_in_c_bypass_regNext_26_1_is_stationary_28;
  reg        [15:0]   io_in_c_bypass_regNext_26_2_data_28;
  reg                 io_in_c_bypass_regNext_26_2_is_stationary_28;
  reg        [15:0]   io_in_c_bypass_regNext_26_3_data_28;
  reg                 io_in_c_bypass_regNext_26_3_is_stationary_28;
  reg        [15:0]   io_in_c_bypass_regNext_27_0_data_28;
  reg                 io_in_c_bypass_regNext_27_0_is_stationary_28;
  reg        [15:0]   io_in_c_bypass_regNext_27_1_data_28;
  reg                 io_in_c_bypass_regNext_27_1_is_stationary_28;
  reg        [15:0]   io_in_c_bypass_regNext_27_2_data_28;
  reg                 io_in_c_bypass_regNext_27_2_is_stationary_28;
  reg        [15:0]   io_in_c_bypass_regNext_27_3_data_28;
  reg                 io_in_c_bypass_regNext_27_3_is_stationary_28;
  reg        [15:0]   io_in_c_bypass_regNext_28_0_data_28;
  reg                 io_in_c_bypass_regNext_28_0_is_stationary_28;
  reg        [15:0]   io_in_c_bypass_regNext_28_1_data_28;
  reg                 io_in_c_bypass_regNext_28_1_is_stationary_28;
  reg        [15:0]   io_in_c_bypass_regNext_28_2_data_28;
  reg                 io_in_c_bypass_regNext_28_2_is_stationary_28;
  reg        [15:0]   io_in_c_bypass_regNext_28_3_data_28;
  reg                 io_in_c_bypass_regNext_28_3_is_stationary_28;
  reg        [15:0]   io_in_c_bypass_regNext_29_0_data_28;
  reg                 io_in_c_bypass_regNext_29_0_is_stationary_28;
  reg        [15:0]   io_in_c_bypass_regNext_29_1_data_28;
  reg                 io_in_c_bypass_regNext_29_1_is_stationary_28;
  reg        [15:0]   io_in_c_bypass_regNext_29_2_data_28;
  reg                 io_in_c_bypass_regNext_29_2_is_stationary_28;
  reg        [15:0]   io_in_c_bypass_regNext_29_3_data_28;
  reg                 io_in_c_bypass_regNext_29_3_is_stationary_28;
  reg        [15:0]   io_in_c_bypass_regNext_30_0_data_28;
  reg                 io_in_c_bypass_regNext_30_0_is_stationary_28;
  reg        [15:0]   io_in_c_bypass_regNext_30_1_data_28;
  reg                 io_in_c_bypass_regNext_30_1_is_stationary_28;
  reg        [15:0]   io_in_c_bypass_regNext_30_2_data_28;
  reg                 io_in_c_bypass_regNext_30_2_is_stationary_28;
  reg        [15:0]   io_in_c_bypass_regNext_30_3_data_28;
  reg                 io_in_c_bypass_regNext_30_3_is_stationary_28;
  reg        [15:0]   io_in_c_bypass_regNext_31_0_data_28;
  reg                 io_in_c_bypass_regNext_31_0_is_stationary_28;
  reg        [15:0]   io_in_c_bypass_regNext_31_1_data_28;
  reg                 io_in_c_bypass_regNext_31_1_is_stationary_28;
  reg        [15:0]   io_in_c_bypass_regNext_31_2_data_28;
  reg                 io_in_c_bypass_regNext_31_2_is_stationary_28;
  reg        [15:0]   io_in_c_bypass_regNext_31_3_data_28;
  reg                 io_in_c_bypass_regNext_31_3_is_stationary_28;
  reg        [15:0]   io_in_c_bypass_regNext_0_0_data_29;
  reg                 io_in_c_bypass_regNext_0_0_is_stationary_29;
  reg        [15:0]   io_in_c_bypass_regNext_0_1_data_29;
  reg                 io_in_c_bypass_regNext_0_1_is_stationary_29;
  reg        [15:0]   io_in_c_bypass_regNext_0_2_data_29;
  reg                 io_in_c_bypass_regNext_0_2_is_stationary_29;
  reg        [15:0]   io_in_c_bypass_regNext_0_3_data_29;
  reg                 io_in_c_bypass_regNext_0_3_is_stationary_29;
  reg        [15:0]   io_in_c_bypass_regNext_1_0_data_29;
  reg                 io_in_c_bypass_regNext_1_0_is_stationary_29;
  reg        [15:0]   io_in_c_bypass_regNext_1_1_data_29;
  reg                 io_in_c_bypass_regNext_1_1_is_stationary_29;
  reg        [15:0]   io_in_c_bypass_regNext_1_2_data_29;
  reg                 io_in_c_bypass_regNext_1_2_is_stationary_29;
  reg        [15:0]   io_in_c_bypass_regNext_1_3_data_29;
  reg                 io_in_c_bypass_regNext_1_3_is_stationary_29;
  reg        [15:0]   io_in_c_bypass_regNext_2_0_data_29;
  reg                 io_in_c_bypass_regNext_2_0_is_stationary_29;
  reg        [15:0]   io_in_c_bypass_regNext_2_1_data_29;
  reg                 io_in_c_bypass_regNext_2_1_is_stationary_29;
  reg        [15:0]   io_in_c_bypass_regNext_2_2_data_29;
  reg                 io_in_c_bypass_regNext_2_2_is_stationary_29;
  reg        [15:0]   io_in_c_bypass_regNext_2_3_data_29;
  reg                 io_in_c_bypass_regNext_2_3_is_stationary_29;
  reg        [15:0]   io_in_c_bypass_regNext_3_0_data_29;
  reg                 io_in_c_bypass_regNext_3_0_is_stationary_29;
  reg        [15:0]   io_in_c_bypass_regNext_3_1_data_29;
  reg                 io_in_c_bypass_regNext_3_1_is_stationary_29;
  reg        [15:0]   io_in_c_bypass_regNext_3_2_data_29;
  reg                 io_in_c_bypass_regNext_3_2_is_stationary_29;
  reg        [15:0]   io_in_c_bypass_regNext_3_3_data_29;
  reg                 io_in_c_bypass_regNext_3_3_is_stationary_29;
  reg        [15:0]   io_in_c_bypass_regNext_4_0_data_29;
  reg                 io_in_c_bypass_regNext_4_0_is_stationary_29;
  reg        [15:0]   io_in_c_bypass_regNext_4_1_data_29;
  reg                 io_in_c_bypass_regNext_4_1_is_stationary_29;
  reg        [15:0]   io_in_c_bypass_regNext_4_2_data_29;
  reg                 io_in_c_bypass_regNext_4_2_is_stationary_29;
  reg        [15:0]   io_in_c_bypass_regNext_4_3_data_29;
  reg                 io_in_c_bypass_regNext_4_3_is_stationary_29;
  reg        [15:0]   io_in_c_bypass_regNext_5_0_data_29;
  reg                 io_in_c_bypass_regNext_5_0_is_stationary_29;
  reg        [15:0]   io_in_c_bypass_regNext_5_1_data_29;
  reg                 io_in_c_bypass_regNext_5_1_is_stationary_29;
  reg        [15:0]   io_in_c_bypass_regNext_5_2_data_29;
  reg                 io_in_c_bypass_regNext_5_2_is_stationary_29;
  reg        [15:0]   io_in_c_bypass_regNext_5_3_data_29;
  reg                 io_in_c_bypass_regNext_5_3_is_stationary_29;
  reg        [15:0]   io_in_c_bypass_regNext_6_0_data_29;
  reg                 io_in_c_bypass_regNext_6_0_is_stationary_29;
  reg        [15:0]   io_in_c_bypass_regNext_6_1_data_29;
  reg                 io_in_c_bypass_regNext_6_1_is_stationary_29;
  reg        [15:0]   io_in_c_bypass_regNext_6_2_data_29;
  reg                 io_in_c_bypass_regNext_6_2_is_stationary_29;
  reg        [15:0]   io_in_c_bypass_regNext_6_3_data_29;
  reg                 io_in_c_bypass_regNext_6_3_is_stationary_29;
  reg        [15:0]   io_in_c_bypass_regNext_7_0_data_29;
  reg                 io_in_c_bypass_regNext_7_0_is_stationary_29;
  reg        [15:0]   io_in_c_bypass_regNext_7_1_data_29;
  reg                 io_in_c_bypass_regNext_7_1_is_stationary_29;
  reg        [15:0]   io_in_c_bypass_regNext_7_2_data_29;
  reg                 io_in_c_bypass_regNext_7_2_is_stationary_29;
  reg        [15:0]   io_in_c_bypass_regNext_7_3_data_29;
  reg                 io_in_c_bypass_regNext_7_3_is_stationary_29;
  reg        [15:0]   io_in_c_bypass_regNext_8_0_data_29;
  reg                 io_in_c_bypass_regNext_8_0_is_stationary_29;
  reg        [15:0]   io_in_c_bypass_regNext_8_1_data_29;
  reg                 io_in_c_bypass_regNext_8_1_is_stationary_29;
  reg        [15:0]   io_in_c_bypass_regNext_8_2_data_29;
  reg                 io_in_c_bypass_regNext_8_2_is_stationary_29;
  reg        [15:0]   io_in_c_bypass_regNext_8_3_data_29;
  reg                 io_in_c_bypass_regNext_8_3_is_stationary_29;
  reg        [15:0]   io_in_c_bypass_regNext_9_0_data_29;
  reg                 io_in_c_bypass_regNext_9_0_is_stationary_29;
  reg        [15:0]   io_in_c_bypass_regNext_9_1_data_29;
  reg                 io_in_c_bypass_regNext_9_1_is_stationary_29;
  reg        [15:0]   io_in_c_bypass_regNext_9_2_data_29;
  reg                 io_in_c_bypass_regNext_9_2_is_stationary_29;
  reg        [15:0]   io_in_c_bypass_regNext_9_3_data_29;
  reg                 io_in_c_bypass_regNext_9_3_is_stationary_29;
  reg        [15:0]   io_in_c_bypass_regNext_10_0_data_29;
  reg                 io_in_c_bypass_regNext_10_0_is_stationary_29;
  reg        [15:0]   io_in_c_bypass_regNext_10_1_data_29;
  reg                 io_in_c_bypass_regNext_10_1_is_stationary_29;
  reg        [15:0]   io_in_c_bypass_regNext_10_2_data_29;
  reg                 io_in_c_bypass_regNext_10_2_is_stationary_29;
  reg        [15:0]   io_in_c_bypass_regNext_10_3_data_29;
  reg                 io_in_c_bypass_regNext_10_3_is_stationary_29;
  reg        [15:0]   io_in_c_bypass_regNext_11_0_data_29;
  reg                 io_in_c_bypass_regNext_11_0_is_stationary_29;
  reg        [15:0]   io_in_c_bypass_regNext_11_1_data_29;
  reg                 io_in_c_bypass_regNext_11_1_is_stationary_29;
  reg        [15:0]   io_in_c_bypass_regNext_11_2_data_29;
  reg                 io_in_c_bypass_regNext_11_2_is_stationary_29;
  reg        [15:0]   io_in_c_bypass_regNext_11_3_data_29;
  reg                 io_in_c_bypass_regNext_11_3_is_stationary_29;
  reg        [15:0]   io_in_c_bypass_regNext_12_0_data_29;
  reg                 io_in_c_bypass_regNext_12_0_is_stationary_29;
  reg        [15:0]   io_in_c_bypass_regNext_12_1_data_29;
  reg                 io_in_c_bypass_regNext_12_1_is_stationary_29;
  reg        [15:0]   io_in_c_bypass_regNext_12_2_data_29;
  reg                 io_in_c_bypass_regNext_12_2_is_stationary_29;
  reg        [15:0]   io_in_c_bypass_regNext_12_3_data_29;
  reg                 io_in_c_bypass_regNext_12_3_is_stationary_29;
  reg        [15:0]   io_in_c_bypass_regNext_13_0_data_29;
  reg                 io_in_c_bypass_regNext_13_0_is_stationary_29;
  reg        [15:0]   io_in_c_bypass_regNext_13_1_data_29;
  reg                 io_in_c_bypass_regNext_13_1_is_stationary_29;
  reg        [15:0]   io_in_c_bypass_regNext_13_2_data_29;
  reg                 io_in_c_bypass_regNext_13_2_is_stationary_29;
  reg        [15:0]   io_in_c_bypass_regNext_13_3_data_29;
  reg                 io_in_c_bypass_regNext_13_3_is_stationary_29;
  reg        [15:0]   io_in_c_bypass_regNext_14_0_data_29;
  reg                 io_in_c_bypass_regNext_14_0_is_stationary_29;
  reg        [15:0]   io_in_c_bypass_regNext_14_1_data_29;
  reg                 io_in_c_bypass_regNext_14_1_is_stationary_29;
  reg        [15:0]   io_in_c_bypass_regNext_14_2_data_29;
  reg                 io_in_c_bypass_regNext_14_2_is_stationary_29;
  reg        [15:0]   io_in_c_bypass_regNext_14_3_data_29;
  reg                 io_in_c_bypass_regNext_14_3_is_stationary_29;
  reg        [15:0]   io_in_c_bypass_regNext_15_0_data_29;
  reg                 io_in_c_bypass_regNext_15_0_is_stationary_29;
  reg        [15:0]   io_in_c_bypass_regNext_15_1_data_29;
  reg                 io_in_c_bypass_regNext_15_1_is_stationary_29;
  reg        [15:0]   io_in_c_bypass_regNext_15_2_data_29;
  reg                 io_in_c_bypass_regNext_15_2_is_stationary_29;
  reg        [15:0]   io_in_c_bypass_regNext_15_3_data_29;
  reg                 io_in_c_bypass_regNext_15_3_is_stationary_29;
  reg        [15:0]   io_in_c_bypass_regNext_16_0_data_29;
  reg                 io_in_c_bypass_regNext_16_0_is_stationary_29;
  reg        [15:0]   io_in_c_bypass_regNext_16_1_data_29;
  reg                 io_in_c_bypass_regNext_16_1_is_stationary_29;
  reg        [15:0]   io_in_c_bypass_regNext_16_2_data_29;
  reg                 io_in_c_bypass_regNext_16_2_is_stationary_29;
  reg        [15:0]   io_in_c_bypass_regNext_16_3_data_29;
  reg                 io_in_c_bypass_regNext_16_3_is_stationary_29;
  reg        [15:0]   io_in_c_bypass_regNext_17_0_data_29;
  reg                 io_in_c_bypass_regNext_17_0_is_stationary_29;
  reg        [15:0]   io_in_c_bypass_regNext_17_1_data_29;
  reg                 io_in_c_bypass_regNext_17_1_is_stationary_29;
  reg        [15:0]   io_in_c_bypass_regNext_17_2_data_29;
  reg                 io_in_c_bypass_regNext_17_2_is_stationary_29;
  reg        [15:0]   io_in_c_bypass_regNext_17_3_data_29;
  reg                 io_in_c_bypass_regNext_17_3_is_stationary_29;
  reg        [15:0]   io_in_c_bypass_regNext_18_0_data_29;
  reg                 io_in_c_bypass_regNext_18_0_is_stationary_29;
  reg        [15:0]   io_in_c_bypass_regNext_18_1_data_29;
  reg                 io_in_c_bypass_regNext_18_1_is_stationary_29;
  reg        [15:0]   io_in_c_bypass_regNext_18_2_data_29;
  reg                 io_in_c_bypass_regNext_18_2_is_stationary_29;
  reg        [15:0]   io_in_c_bypass_regNext_18_3_data_29;
  reg                 io_in_c_bypass_regNext_18_3_is_stationary_29;
  reg        [15:0]   io_in_c_bypass_regNext_19_0_data_29;
  reg                 io_in_c_bypass_regNext_19_0_is_stationary_29;
  reg        [15:0]   io_in_c_bypass_regNext_19_1_data_29;
  reg                 io_in_c_bypass_regNext_19_1_is_stationary_29;
  reg        [15:0]   io_in_c_bypass_regNext_19_2_data_29;
  reg                 io_in_c_bypass_regNext_19_2_is_stationary_29;
  reg        [15:0]   io_in_c_bypass_regNext_19_3_data_29;
  reg                 io_in_c_bypass_regNext_19_3_is_stationary_29;
  reg        [15:0]   io_in_c_bypass_regNext_20_0_data_29;
  reg                 io_in_c_bypass_regNext_20_0_is_stationary_29;
  reg        [15:0]   io_in_c_bypass_regNext_20_1_data_29;
  reg                 io_in_c_bypass_regNext_20_1_is_stationary_29;
  reg        [15:0]   io_in_c_bypass_regNext_20_2_data_29;
  reg                 io_in_c_bypass_regNext_20_2_is_stationary_29;
  reg        [15:0]   io_in_c_bypass_regNext_20_3_data_29;
  reg                 io_in_c_bypass_regNext_20_3_is_stationary_29;
  reg        [15:0]   io_in_c_bypass_regNext_21_0_data_29;
  reg                 io_in_c_bypass_regNext_21_0_is_stationary_29;
  reg        [15:0]   io_in_c_bypass_regNext_21_1_data_29;
  reg                 io_in_c_bypass_regNext_21_1_is_stationary_29;
  reg        [15:0]   io_in_c_bypass_regNext_21_2_data_29;
  reg                 io_in_c_bypass_regNext_21_2_is_stationary_29;
  reg        [15:0]   io_in_c_bypass_regNext_21_3_data_29;
  reg                 io_in_c_bypass_regNext_21_3_is_stationary_29;
  reg        [15:0]   io_in_c_bypass_regNext_22_0_data_29;
  reg                 io_in_c_bypass_regNext_22_0_is_stationary_29;
  reg        [15:0]   io_in_c_bypass_regNext_22_1_data_29;
  reg                 io_in_c_bypass_regNext_22_1_is_stationary_29;
  reg        [15:0]   io_in_c_bypass_regNext_22_2_data_29;
  reg                 io_in_c_bypass_regNext_22_2_is_stationary_29;
  reg        [15:0]   io_in_c_bypass_regNext_22_3_data_29;
  reg                 io_in_c_bypass_regNext_22_3_is_stationary_29;
  reg        [15:0]   io_in_c_bypass_regNext_23_0_data_29;
  reg                 io_in_c_bypass_regNext_23_0_is_stationary_29;
  reg        [15:0]   io_in_c_bypass_regNext_23_1_data_29;
  reg                 io_in_c_bypass_regNext_23_1_is_stationary_29;
  reg        [15:0]   io_in_c_bypass_regNext_23_2_data_29;
  reg                 io_in_c_bypass_regNext_23_2_is_stationary_29;
  reg        [15:0]   io_in_c_bypass_regNext_23_3_data_29;
  reg                 io_in_c_bypass_regNext_23_3_is_stationary_29;
  reg        [15:0]   io_in_c_bypass_regNext_24_0_data_29;
  reg                 io_in_c_bypass_regNext_24_0_is_stationary_29;
  reg        [15:0]   io_in_c_bypass_regNext_24_1_data_29;
  reg                 io_in_c_bypass_regNext_24_1_is_stationary_29;
  reg        [15:0]   io_in_c_bypass_regNext_24_2_data_29;
  reg                 io_in_c_bypass_regNext_24_2_is_stationary_29;
  reg        [15:0]   io_in_c_bypass_regNext_24_3_data_29;
  reg                 io_in_c_bypass_regNext_24_3_is_stationary_29;
  reg        [15:0]   io_in_c_bypass_regNext_25_0_data_29;
  reg                 io_in_c_bypass_regNext_25_0_is_stationary_29;
  reg        [15:0]   io_in_c_bypass_regNext_25_1_data_29;
  reg                 io_in_c_bypass_regNext_25_1_is_stationary_29;
  reg        [15:0]   io_in_c_bypass_regNext_25_2_data_29;
  reg                 io_in_c_bypass_regNext_25_2_is_stationary_29;
  reg        [15:0]   io_in_c_bypass_regNext_25_3_data_29;
  reg                 io_in_c_bypass_regNext_25_3_is_stationary_29;
  reg        [15:0]   io_in_c_bypass_regNext_26_0_data_29;
  reg                 io_in_c_bypass_regNext_26_0_is_stationary_29;
  reg        [15:0]   io_in_c_bypass_regNext_26_1_data_29;
  reg                 io_in_c_bypass_regNext_26_1_is_stationary_29;
  reg        [15:0]   io_in_c_bypass_regNext_26_2_data_29;
  reg                 io_in_c_bypass_regNext_26_2_is_stationary_29;
  reg        [15:0]   io_in_c_bypass_regNext_26_3_data_29;
  reg                 io_in_c_bypass_regNext_26_3_is_stationary_29;
  reg        [15:0]   io_in_c_bypass_regNext_27_0_data_29;
  reg                 io_in_c_bypass_regNext_27_0_is_stationary_29;
  reg        [15:0]   io_in_c_bypass_regNext_27_1_data_29;
  reg                 io_in_c_bypass_regNext_27_1_is_stationary_29;
  reg        [15:0]   io_in_c_bypass_regNext_27_2_data_29;
  reg                 io_in_c_bypass_regNext_27_2_is_stationary_29;
  reg        [15:0]   io_in_c_bypass_regNext_27_3_data_29;
  reg                 io_in_c_bypass_regNext_27_3_is_stationary_29;
  reg        [15:0]   io_in_c_bypass_regNext_28_0_data_29;
  reg                 io_in_c_bypass_regNext_28_0_is_stationary_29;
  reg        [15:0]   io_in_c_bypass_regNext_28_1_data_29;
  reg                 io_in_c_bypass_regNext_28_1_is_stationary_29;
  reg        [15:0]   io_in_c_bypass_regNext_28_2_data_29;
  reg                 io_in_c_bypass_regNext_28_2_is_stationary_29;
  reg        [15:0]   io_in_c_bypass_regNext_28_3_data_29;
  reg                 io_in_c_bypass_regNext_28_3_is_stationary_29;
  reg        [15:0]   io_in_c_bypass_regNext_29_0_data_29;
  reg                 io_in_c_bypass_regNext_29_0_is_stationary_29;
  reg        [15:0]   io_in_c_bypass_regNext_29_1_data_29;
  reg                 io_in_c_bypass_regNext_29_1_is_stationary_29;
  reg        [15:0]   io_in_c_bypass_regNext_29_2_data_29;
  reg                 io_in_c_bypass_regNext_29_2_is_stationary_29;
  reg        [15:0]   io_in_c_bypass_regNext_29_3_data_29;
  reg                 io_in_c_bypass_regNext_29_3_is_stationary_29;
  reg        [15:0]   io_in_c_bypass_regNext_30_0_data_29;
  reg                 io_in_c_bypass_regNext_30_0_is_stationary_29;
  reg        [15:0]   io_in_c_bypass_regNext_30_1_data_29;
  reg                 io_in_c_bypass_regNext_30_1_is_stationary_29;
  reg        [15:0]   io_in_c_bypass_regNext_30_2_data_29;
  reg                 io_in_c_bypass_regNext_30_2_is_stationary_29;
  reg        [15:0]   io_in_c_bypass_regNext_30_3_data_29;
  reg                 io_in_c_bypass_regNext_30_3_is_stationary_29;
  reg        [15:0]   io_in_c_bypass_regNext_31_0_data_29;
  reg                 io_in_c_bypass_regNext_31_0_is_stationary_29;
  reg        [15:0]   io_in_c_bypass_regNext_31_1_data_29;
  reg                 io_in_c_bypass_regNext_31_1_is_stationary_29;
  reg        [15:0]   io_in_c_bypass_regNext_31_2_data_29;
  reg                 io_in_c_bypass_regNext_31_2_is_stationary_29;
  reg        [15:0]   io_in_c_bypass_regNext_31_3_data_29;
  reg                 io_in_c_bypass_regNext_31_3_is_stationary_29;
  reg        [15:0]   io_in_c_bypass_regNext_0_0_data_30;
  reg                 io_in_c_bypass_regNext_0_0_is_stationary_30;
  reg        [15:0]   io_in_c_bypass_regNext_0_1_data_30;
  reg                 io_in_c_bypass_regNext_0_1_is_stationary_30;
  reg        [15:0]   io_in_c_bypass_regNext_0_2_data_30;
  reg                 io_in_c_bypass_regNext_0_2_is_stationary_30;
  reg        [15:0]   io_in_c_bypass_regNext_0_3_data_30;
  reg                 io_in_c_bypass_regNext_0_3_is_stationary_30;
  reg        [15:0]   io_in_c_bypass_regNext_1_0_data_30;
  reg                 io_in_c_bypass_regNext_1_0_is_stationary_30;
  reg        [15:0]   io_in_c_bypass_regNext_1_1_data_30;
  reg                 io_in_c_bypass_regNext_1_1_is_stationary_30;
  reg        [15:0]   io_in_c_bypass_regNext_1_2_data_30;
  reg                 io_in_c_bypass_regNext_1_2_is_stationary_30;
  reg        [15:0]   io_in_c_bypass_regNext_1_3_data_30;
  reg                 io_in_c_bypass_regNext_1_3_is_stationary_30;
  reg        [15:0]   io_in_c_bypass_regNext_2_0_data_30;
  reg                 io_in_c_bypass_regNext_2_0_is_stationary_30;
  reg        [15:0]   io_in_c_bypass_regNext_2_1_data_30;
  reg                 io_in_c_bypass_regNext_2_1_is_stationary_30;
  reg        [15:0]   io_in_c_bypass_regNext_2_2_data_30;
  reg                 io_in_c_bypass_regNext_2_2_is_stationary_30;
  reg        [15:0]   io_in_c_bypass_regNext_2_3_data_30;
  reg                 io_in_c_bypass_regNext_2_3_is_stationary_30;
  reg        [15:0]   io_in_c_bypass_regNext_3_0_data_30;
  reg                 io_in_c_bypass_regNext_3_0_is_stationary_30;
  reg        [15:0]   io_in_c_bypass_regNext_3_1_data_30;
  reg                 io_in_c_bypass_regNext_3_1_is_stationary_30;
  reg        [15:0]   io_in_c_bypass_regNext_3_2_data_30;
  reg                 io_in_c_bypass_regNext_3_2_is_stationary_30;
  reg        [15:0]   io_in_c_bypass_regNext_3_3_data_30;
  reg                 io_in_c_bypass_regNext_3_3_is_stationary_30;
  reg        [15:0]   io_in_c_bypass_regNext_4_0_data_30;
  reg                 io_in_c_bypass_regNext_4_0_is_stationary_30;
  reg        [15:0]   io_in_c_bypass_regNext_4_1_data_30;
  reg                 io_in_c_bypass_regNext_4_1_is_stationary_30;
  reg        [15:0]   io_in_c_bypass_regNext_4_2_data_30;
  reg                 io_in_c_bypass_regNext_4_2_is_stationary_30;
  reg        [15:0]   io_in_c_bypass_regNext_4_3_data_30;
  reg                 io_in_c_bypass_regNext_4_3_is_stationary_30;
  reg        [15:0]   io_in_c_bypass_regNext_5_0_data_30;
  reg                 io_in_c_bypass_regNext_5_0_is_stationary_30;
  reg        [15:0]   io_in_c_bypass_regNext_5_1_data_30;
  reg                 io_in_c_bypass_regNext_5_1_is_stationary_30;
  reg        [15:0]   io_in_c_bypass_regNext_5_2_data_30;
  reg                 io_in_c_bypass_regNext_5_2_is_stationary_30;
  reg        [15:0]   io_in_c_bypass_regNext_5_3_data_30;
  reg                 io_in_c_bypass_regNext_5_3_is_stationary_30;
  reg        [15:0]   io_in_c_bypass_regNext_6_0_data_30;
  reg                 io_in_c_bypass_regNext_6_0_is_stationary_30;
  reg        [15:0]   io_in_c_bypass_regNext_6_1_data_30;
  reg                 io_in_c_bypass_regNext_6_1_is_stationary_30;
  reg        [15:0]   io_in_c_bypass_regNext_6_2_data_30;
  reg                 io_in_c_bypass_regNext_6_2_is_stationary_30;
  reg        [15:0]   io_in_c_bypass_regNext_6_3_data_30;
  reg                 io_in_c_bypass_regNext_6_3_is_stationary_30;
  reg        [15:0]   io_in_c_bypass_regNext_7_0_data_30;
  reg                 io_in_c_bypass_regNext_7_0_is_stationary_30;
  reg        [15:0]   io_in_c_bypass_regNext_7_1_data_30;
  reg                 io_in_c_bypass_regNext_7_1_is_stationary_30;
  reg        [15:0]   io_in_c_bypass_regNext_7_2_data_30;
  reg                 io_in_c_bypass_regNext_7_2_is_stationary_30;
  reg        [15:0]   io_in_c_bypass_regNext_7_3_data_30;
  reg                 io_in_c_bypass_regNext_7_3_is_stationary_30;
  reg        [15:0]   io_in_c_bypass_regNext_8_0_data_30;
  reg                 io_in_c_bypass_regNext_8_0_is_stationary_30;
  reg        [15:0]   io_in_c_bypass_regNext_8_1_data_30;
  reg                 io_in_c_bypass_regNext_8_1_is_stationary_30;
  reg        [15:0]   io_in_c_bypass_regNext_8_2_data_30;
  reg                 io_in_c_bypass_regNext_8_2_is_stationary_30;
  reg        [15:0]   io_in_c_bypass_regNext_8_3_data_30;
  reg                 io_in_c_bypass_regNext_8_3_is_stationary_30;
  reg        [15:0]   io_in_c_bypass_regNext_9_0_data_30;
  reg                 io_in_c_bypass_regNext_9_0_is_stationary_30;
  reg        [15:0]   io_in_c_bypass_regNext_9_1_data_30;
  reg                 io_in_c_bypass_regNext_9_1_is_stationary_30;
  reg        [15:0]   io_in_c_bypass_regNext_9_2_data_30;
  reg                 io_in_c_bypass_regNext_9_2_is_stationary_30;
  reg        [15:0]   io_in_c_bypass_regNext_9_3_data_30;
  reg                 io_in_c_bypass_regNext_9_3_is_stationary_30;
  reg        [15:0]   io_in_c_bypass_regNext_10_0_data_30;
  reg                 io_in_c_bypass_regNext_10_0_is_stationary_30;
  reg        [15:0]   io_in_c_bypass_regNext_10_1_data_30;
  reg                 io_in_c_bypass_regNext_10_1_is_stationary_30;
  reg        [15:0]   io_in_c_bypass_regNext_10_2_data_30;
  reg                 io_in_c_bypass_regNext_10_2_is_stationary_30;
  reg        [15:0]   io_in_c_bypass_regNext_10_3_data_30;
  reg                 io_in_c_bypass_regNext_10_3_is_stationary_30;
  reg        [15:0]   io_in_c_bypass_regNext_11_0_data_30;
  reg                 io_in_c_bypass_regNext_11_0_is_stationary_30;
  reg        [15:0]   io_in_c_bypass_regNext_11_1_data_30;
  reg                 io_in_c_bypass_regNext_11_1_is_stationary_30;
  reg        [15:0]   io_in_c_bypass_regNext_11_2_data_30;
  reg                 io_in_c_bypass_regNext_11_2_is_stationary_30;
  reg        [15:0]   io_in_c_bypass_regNext_11_3_data_30;
  reg                 io_in_c_bypass_regNext_11_3_is_stationary_30;
  reg        [15:0]   io_in_c_bypass_regNext_12_0_data_30;
  reg                 io_in_c_bypass_regNext_12_0_is_stationary_30;
  reg        [15:0]   io_in_c_bypass_regNext_12_1_data_30;
  reg                 io_in_c_bypass_regNext_12_1_is_stationary_30;
  reg        [15:0]   io_in_c_bypass_regNext_12_2_data_30;
  reg                 io_in_c_bypass_regNext_12_2_is_stationary_30;
  reg        [15:0]   io_in_c_bypass_regNext_12_3_data_30;
  reg                 io_in_c_bypass_regNext_12_3_is_stationary_30;
  reg        [15:0]   io_in_c_bypass_regNext_13_0_data_30;
  reg                 io_in_c_bypass_regNext_13_0_is_stationary_30;
  reg        [15:0]   io_in_c_bypass_regNext_13_1_data_30;
  reg                 io_in_c_bypass_regNext_13_1_is_stationary_30;
  reg        [15:0]   io_in_c_bypass_regNext_13_2_data_30;
  reg                 io_in_c_bypass_regNext_13_2_is_stationary_30;
  reg        [15:0]   io_in_c_bypass_regNext_13_3_data_30;
  reg                 io_in_c_bypass_regNext_13_3_is_stationary_30;
  reg        [15:0]   io_in_c_bypass_regNext_14_0_data_30;
  reg                 io_in_c_bypass_regNext_14_0_is_stationary_30;
  reg        [15:0]   io_in_c_bypass_regNext_14_1_data_30;
  reg                 io_in_c_bypass_regNext_14_1_is_stationary_30;
  reg        [15:0]   io_in_c_bypass_regNext_14_2_data_30;
  reg                 io_in_c_bypass_regNext_14_2_is_stationary_30;
  reg        [15:0]   io_in_c_bypass_regNext_14_3_data_30;
  reg                 io_in_c_bypass_regNext_14_3_is_stationary_30;
  reg        [15:0]   io_in_c_bypass_regNext_15_0_data_30;
  reg                 io_in_c_bypass_regNext_15_0_is_stationary_30;
  reg        [15:0]   io_in_c_bypass_regNext_15_1_data_30;
  reg                 io_in_c_bypass_regNext_15_1_is_stationary_30;
  reg        [15:0]   io_in_c_bypass_regNext_15_2_data_30;
  reg                 io_in_c_bypass_regNext_15_2_is_stationary_30;
  reg        [15:0]   io_in_c_bypass_regNext_15_3_data_30;
  reg                 io_in_c_bypass_regNext_15_3_is_stationary_30;
  reg        [15:0]   io_in_c_bypass_regNext_16_0_data_30;
  reg                 io_in_c_bypass_regNext_16_0_is_stationary_30;
  reg        [15:0]   io_in_c_bypass_regNext_16_1_data_30;
  reg                 io_in_c_bypass_regNext_16_1_is_stationary_30;
  reg        [15:0]   io_in_c_bypass_regNext_16_2_data_30;
  reg                 io_in_c_bypass_regNext_16_2_is_stationary_30;
  reg        [15:0]   io_in_c_bypass_regNext_16_3_data_30;
  reg                 io_in_c_bypass_regNext_16_3_is_stationary_30;
  reg        [15:0]   io_in_c_bypass_regNext_17_0_data_30;
  reg                 io_in_c_bypass_regNext_17_0_is_stationary_30;
  reg        [15:0]   io_in_c_bypass_regNext_17_1_data_30;
  reg                 io_in_c_bypass_regNext_17_1_is_stationary_30;
  reg        [15:0]   io_in_c_bypass_regNext_17_2_data_30;
  reg                 io_in_c_bypass_regNext_17_2_is_stationary_30;
  reg        [15:0]   io_in_c_bypass_regNext_17_3_data_30;
  reg                 io_in_c_bypass_regNext_17_3_is_stationary_30;
  reg        [15:0]   io_in_c_bypass_regNext_18_0_data_30;
  reg                 io_in_c_bypass_regNext_18_0_is_stationary_30;
  reg        [15:0]   io_in_c_bypass_regNext_18_1_data_30;
  reg                 io_in_c_bypass_regNext_18_1_is_stationary_30;
  reg        [15:0]   io_in_c_bypass_regNext_18_2_data_30;
  reg                 io_in_c_bypass_regNext_18_2_is_stationary_30;
  reg        [15:0]   io_in_c_bypass_regNext_18_3_data_30;
  reg                 io_in_c_bypass_regNext_18_3_is_stationary_30;
  reg        [15:0]   io_in_c_bypass_regNext_19_0_data_30;
  reg                 io_in_c_bypass_regNext_19_0_is_stationary_30;
  reg        [15:0]   io_in_c_bypass_regNext_19_1_data_30;
  reg                 io_in_c_bypass_regNext_19_1_is_stationary_30;
  reg        [15:0]   io_in_c_bypass_regNext_19_2_data_30;
  reg                 io_in_c_bypass_regNext_19_2_is_stationary_30;
  reg        [15:0]   io_in_c_bypass_regNext_19_3_data_30;
  reg                 io_in_c_bypass_regNext_19_3_is_stationary_30;
  reg        [15:0]   io_in_c_bypass_regNext_20_0_data_30;
  reg                 io_in_c_bypass_regNext_20_0_is_stationary_30;
  reg        [15:0]   io_in_c_bypass_regNext_20_1_data_30;
  reg                 io_in_c_bypass_regNext_20_1_is_stationary_30;
  reg        [15:0]   io_in_c_bypass_regNext_20_2_data_30;
  reg                 io_in_c_bypass_regNext_20_2_is_stationary_30;
  reg        [15:0]   io_in_c_bypass_regNext_20_3_data_30;
  reg                 io_in_c_bypass_regNext_20_3_is_stationary_30;
  reg        [15:0]   io_in_c_bypass_regNext_21_0_data_30;
  reg                 io_in_c_bypass_regNext_21_0_is_stationary_30;
  reg        [15:0]   io_in_c_bypass_regNext_21_1_data_30;
  reg                 io_in_c_bypass_regNext_21_1_is_stationary_30;
  reg        [15:0]   io_in_c_bypass_regNext_21_2_data_30;
  reg                 io_in_c_bypass_regNext_21_2_is_stationary_30;
  reg        [15:0]   io_in_c_bypass_regNext_21_3_data_30;
  reg                 io_in_c_bypass_regNext_21_3_is_stationary_30;
  reg        [15:0]   io_in_c_bypass_regNext_22_0_data_30;
  reg                 io_in_c_bypass_regNext_22_0_is_stationary_30;
  reg        [15:0]   io_in_c_bypass_regNext_22_1_data_30;
  reg                 io_in_c_bypass_regNext_22_1_is_stationary_30;
  reg        [15:0]   io_in_c_bypass_regNext_22_2_data_30;
  reg                 io_in_c_bypass_regNext_22_2_is_stationary_30;
  reg        [15:0]   io_in_c_bypass_regNext_22_3_data_30;
  reg                 io_in_c_bypass_regNext_22_3_is_stationary_30;
  reg        [15:0]   io_in_c_bypass_regNext_23_0_data_30;
  reg                 io_in_c_bypass_regNext_23_0_is_stationary_30;
  reg        [15:0]   io_in_c_bypass_regNext_23_1_data_30;
  reg                 io_in_c_bypass_regNext_23_1_is_stationary_30;
  reg        [15:0]   io_in_c_bypass_regNext_23_2_data_30;
  reg                 io_in_c_bypass_regNext_23_2_is_stationary_30;
  reg        [15:0]   io_in_c_bypass_regNext_23_3_data_30;
  reg                 io_in_c_bypass_regNext_23_3_is_stationary_30;
  reg        [15:0]   io_in_c_bypass_regNext_24_0_data_30;
  reg                 io_in_c_bypass_regNext_24_0_is_stationary_30;
  reg        [15:0]   io_in_c_bypass_regNext_24_1_data_30;
  reg                 io_in_c_bypass_regNext_24_1_is_stationary_30;
  reg        [15:0]   io_in_c_bypass_regNext_24_2_data_30;
  reg                 io_in_c_bypass_regNext_24_2_is_stationary_30;
  reg        [15:0]   io_in_c_bypass_regNext_24_3_data_30;
  reg                 io_in_c_bypass_regNext_24_3_is_stationary_30;
  reg        [15:0]   io_in_c_bypass_regNext_25_0_data_30;
  reg                 io_in_c_bypass_regNext_25_0_is_stationary_30;
  reg        [15:0]   io_in_c_bypass_regNext_25_1_data_30;
  reg                 io_in_c_bypass_regNext_25_1_is_stationary_30;
  reg        [15:0]   io_in_c_bypass_regNext_25_2_data_30;
  reg                 io_in_c_bypass_regNext_25_2_is_stationary_30;
  reg        [15:0]   io_in_c_bypass_regNext_25_3_data_30;
  reg                 io_in_c_bypass_regNext_25_3_is_stationary_30;
  reg        [15:0]   io_in_c_bypass_regNext_26_0_data_30;
  reg                 io_in_c_bypass_regNext_26_0_is_stationary_30;
  reg        [15:0]   io_in_c_bypass_regNext_26_1_data_30;
  reg                 io_in_c_bypass_regNext_26_1_is_stationary_30;
  reg        [15:0]   io_in_c_bypass_regNext_26_2_data_30;
  reg                 io_in_c_bypass_regNext_26_2_is_stationary_30;
  reg        [15:0]   io_in_c_bypass_regNext_26_3_data_30;
  reg                 io_in_c_bypass_regNext_26_3_is_stationary_30;
  reg        [15:0]   io_in_c_bypass_regNext_27_0_data_30;
  reg                 io_in_c_bypass_regNext_27_0_is_stationary_30;
  reg        [15:0]   io_in_c_bypass_regNext_27_1_data_30;
  reg                 io_in_c_bypass_regNext_27_1_is_stationary_30;
  reg        [15:0]   io_in_c_bypass_regNext_27_2_data_30;
  reg                 io_in_c_bypass_regNext_27_2_is_stationary_30;
  reg        [15:0]   io_in_c_bypass_regNext_27_3_data_30;
  reg                 io_in_c_bypass_regNext_27_3_is_stationary_30;
  reg        [15:0]   io_in_c_bypass_regNext_28_0_data_30;
  reg                 io_in_c_bypass_regNext_28_0_is_stationary_30;
  reg        [15:0]   io_in_c_bypass_regNext_28_1_data_30;
  reg                 io_in_c_bypass_regNext_28_1_is_stationary_30;
  reg        [15:0]   io_in_c_bypass_regNext_28_2_data_30;
  reg                 io_in_c_bypass_regNext_28_2_is_stationary_30;
  reg        [15:0]   io_in_c_bypass_regNext_28_3_data_30;
  reg                 io_in_c_bypass_regNext_28_3_is_stationary_30;
  reg        [15:0]   io_in_c_bypass_regNext_29_0_data_30;
  reg                 io_in_c_bypass_regNext_29_0_is_stationary_30;
  reg        [15:0]   io_in_c_bypass_regNext_29_1_data_30;
  reg                 io_in_c_bypass_regNext_29_1_is_stationary_30;
  reg        [15:0]   io_in_c_bypass_regNext_29_2_data_30;
  reg                 io_in_c_bypass_regNext_29_2_is_stationary_30;
  reg        [15:0]   io_in_c_bypass_regNext_29_3_data_30;
  reg                 io_in_c_bypass_regNext_29_3_is_stationary_30;
  reg        [15:0]   io_in_c_bypass_regNext_30_0_data_30;
  reg                 io_in_c_bypass_regNext_30_0_is_stationary_30;
  reg        [15:0]   io_in_c_bypass_regNext_30_1_data_30;
  reg                 io_in_c_bypass_regNext_30_1_is_stationary_30;
  reg        [15:0]   io_in_c_bypass_regNext_30_2_data_30;
  reg                 io_in_c_bypass_regNext_30_2_is_stationary_30;
  reg        [15:0]   io_in_c_bypass_regNext_30_3_data_30;
  reg                 io_in_c_bypass_regNext_30_3_is_stationary_30;
  reg        [15:0]   io_in_c_bypass_regNext_31_0_data_30;
  reg                 io_in_c_bypass_regNext_31_0_is_stationary_30;
  reg        [15:0]   io_in_c_bypass_regNext_31_1_data_30;
  reg                 io_in_c_bypass_regNext_31_1_is_stationary_30;
  reg        [15:0]   io_in_c_bypass_regNext_31_2_data_30;
  reg                 io_in_c_bypass_regNext_31_2_is_stationary_30;
  reg        [15:0]   io_in_c_bypass_regNext_31_3_data_30;
  reg                 io_in_c_bypass_regNext_31_3_is_stationary_30;
  reg                 io_in_r_input_from_bypass_regNext_0;
  reg                 io_in_r_input_from_bypass_regNext_1;
  reg                 io_in_r_input_from_bypass_regNext_2;
  reg                 io_in_r_input_from_bypass_regNext_3;
  reg                 io_in_r_input_from_bypass_regNext_4;
  reg                 io_in_r_input_from_bypass_regNext_5;
  reg                 io_in_r_input_from_bypass_regNext_6;
  reg                 io_in_r_input_from_bypass_regNext_7;
  reg                 io_in_r_input_from_bypass_regNext_8;
  reg                 io_in_r_input_from_bypass_regNext_9;
  reg                 io_in_r_input_from_bypass_regNext_10;
  reg                 io_in_r_input_from_bypass_regNext_11;
  reg                 io_in_r_input_from_bypass_regNext_12;
  reg                 io_in_r_input_from_bypass_regNext_13;
  reg                 io_in_r_input_from_bypass_regNext_14;
  reg                 io_in_r_input_from_bypass_regNext_15;
  reg                 io_in_r_input_from_bypass_regNext_16;
  reg                 io_in_r_input_from_bypass_regNext_17;
  reg                 io_in_r_input_from_bypass_regNext_18;
  reg                 io_in_r_input_from_bypass_regNext_19;
  reg                 io_in_r_input_from_bypass_regNext_20;
  reg                 io_in_r_input_from_bypass_regNext_21;
  reg                 io_in_r_input_from_bypass_regNext_22;
  reg                 io_in_r_input_from_bypass_regNext_23;
  reg                 io_in_r_input_from_bypass_regNext_24;
  reg                 io_in_r_input_from_bypass_regNext_25;
  reg                 io_in_r_input_from_bypass_regNext_26;
  reg                 io_in_r_input_from_bypass_regNext_27;
  reg                 io_in_r_input_from_bypass_regNext_28;
  reg                 io_in_r_input_from_bypass_regNext_29;
  reg                 io_in_r_input_from_bypass_regNext_30;
  reg                 io_in_r_input_from_bypass_regNext_31;
  reg                 io_in_c_input_from_bypass_regNext_0;
  reg                 io_in_c_input_from_bypass_regNext_1;
  reg                 io_in_c_input_from_bypass_regNext_2;
  reg                 io_in_c_input_from_bypass_regNext_3;
  reg                 io_in_c_input_from_bypass_regNext_4;
  reg                 io_in_c_input_from_bypass_regNext_5;
  reg                 io_in_c_input_from_bypass_regNext_6;
  reg                 io_in_c_input_from_bypass_regNext_7;
  reg                 io_in_c_input_from_bypass_regNext_8;
  reg                 io_in_c_input_from_bypass_regNext_9;
  reg                 io_in_c_input_from_bypass_regNext_10;
  reg                 io_in_c_input_from_bypass_regNext_11;
  reg                 io_in_c_input_from_bypass_regNext_12;
  reg                 io_in_c_input_from_bypass_regNext_13;
  reg                 io_in_c_input_from_bypass_regNext_14;
  reg                 io_in_c_input_from_bypass_regNext_15;
  reg                 io_in_c_input_from_bypass_regNext_16;
  reg                 io_in_c_input_from_bypass_regNext_17;
  reg                 io_in_c_input_from_bypass_regNext_18;
  reg                 io_in_c_input_from_bypass_regNext_19;
  reg                 io_in_c_input_from_bypass_regNext_20;
  reg                 io_in_c_input_from_bypass_regNext_21;
  reg                 io_in_c_input_from_bypass_regNext_22;
  reg                 io_in_c_input_from_bypass_regNext_23;
  reg                 io_in_c_input_from_bypass_regNext_24;
  reg                 io_in_c_input_from_bypass_regNext_25;
  reg                 io_in_c_input_from_bypass_regNext_26;
  reg                 io_in_c_input_from_bypass_regNext_27;
  reg                 io_in_c_input_from_bypass_regNext_28;
  reg                 io_in_c_input_from_bypass_regNext_29;
  reg                 io_in_c_input_from_bypass_regNext_30;
  reg                 io_in_c_input_from_bypass_regNext_31;

  PEWSOS_15 pes_0_0 (
    .io_in_r_data           (in_r_0_data[15:0]             ), //i
    .io_in_r_load_store     (in_r_0_load_store             ), //i
    .io_in_r_df_is_ws       (in_r_0_df_is_ws               ), //i
    .io_in_r_stall          (in_r_0_stall                  ), //i
    .io_out_r_data          (pes_0_0_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pes_0_0_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pes_0_0_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pes_0_0_io_out_r_stall        ), //o
    .io_in_c_data           (in_c_0_data[15:0]             ), //i
    .io_in_c_is_stationary  (in_c_0_is_stationary          ), //i
    .io_out_c_data          (pes_0_0_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pes_0_0_io_out_c_is_stationary), //o
    .clk                    (clk                           ), //i
    .reset                  (reset                         )  //i
  );
  PEWSOS_15 pes_0_1 (
    .io_in_r_data           (pes_0_0_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pes_0_0_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pes_0_0_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pes_0_0_io_out_r_stall        ), //i
    .io_out_r_data          (pes_0_1_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pes_0_1_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pes_0_1_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pes_0_1_io_out_r_stall        ), //o
    .io_in_c_data           (in_c_1_data[15:0]             ), //i
    .io_in_c_is_stationary  (in_c_1_is_stationary          ), //i
    .io_out_c_data          (pes_0_1_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pes_0_1_io_out_c_is_stationary), //o
    .clk                    (clk                           ), //i
    .reset                  (reset                         )  //i
  );
  PEWSOS_15 pes_0_2 (
    .io_in_r_data           (pes_0_1_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pes_0_1_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pes_0_1_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pes_0_1_io_out_r_stall        ), //i
    .io_out_r_data          (pes_0_2_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pes_0_2_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pes_0_2_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pes_0_2_io_out_r_stall        ), //o
    .io_in_c_data           (in_c_2_data[15:0]             ), //i
    .io_in_c_is_stationary  (in_c_2_is_stationary          ), //i
    .io_out_c_data          (pes_0_2_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pes_0_2_io_out_c_is_stationary), //o
    .clk                    (clk                           ), //i
    .reset                  (reset                         )  //i
  );
  PEWSOS_15 pes_0_3 (
    .io_in_r_data           (pes_0_2_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pes_0_2_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pes_0_2_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pes_0_2_io_out_r_stall        ), //i
    .io_out_r_data          (pes_0_3_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pes_0_3_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pes_0_3_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pes_0_3_io_out_r_stall        ), //o
    .io_in_c_data           (in_c_3_data[15:0]             ), //i
    .io_in_c_is_stationary  (in_c_3_is_stationary          ), //i
    .io_out_c_data          (pes_0_3_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pes_0_3_io_out_c_is_stationary), //o
    .clk                    (clk                           ), //i
    .reset                  (reset                         )  //i
  );
  PEWSOS_15 pes_1_0 (
    .io_in_r_data           (in_r_1_data[15:0]             ), //i
    .io_in_r_load_store     (in_r_1_load_store             ), //i
    .io_in_r_df_is_ws       (in_r_1_df_is_ws               ), //i
    .io_in_r_stall          (in_r_1_stall                  ), //i
    .io_out_r_data          (pes_1_0_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pes_1_0_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pes_1_0_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pes_1_0_io_out_r_stall        ), //o
    .io_in_c_data           (pes_0_0_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pes_0_0_io_out_c_is_stationary), //i
    .io_out_c_data          (pes_1_0_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pes_1_0_io_out_c_is_stationary), //o
    .clk                    (clk                           ), //i
    .reset                  (reset                         )  //i
  );
  PEWSOS_15 pes_1_1 (
    .io_in_r_data           (pes_1_0_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pes_1_0_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pes_1_0_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pes_1_0_io_out_r_stall        ), //i
    .io_out_r_data          (pes_1_1_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pes_1_1_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pes_1_1_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pes_1_1_io_out_r_stall        ), //o
    .io_in_c_data           (pes_0_1_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pes_0_1_io_out_c_is_stationary), //i
    .io_out_c_data          (pes_1_1_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pes_1_1_io_out_c_is_stationary), //o
    .clk                    (clk                           ), //i
    .reset                  (reset                         )  //i
  );
  PEWSOS_15 pes_1_2 (
    .io_in_r_data           (pes_1_1_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pes_1_1_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pes_1_1_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pes_1_1_io_out_r_stall        ), //i
    .io_out_r_data          (pes_1_2_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pes_1_2_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pes_1_2_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pes_1_2_io_out_r_stall        ), //o
    .io_in_c_data           (pes_0_2_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pes_0_2_io_out_c_is_stationary), //i
    .io_out_c_data          (pes_1_2_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pes_1_2_io_out_c_is_stationary), //o
    .clk                    (clk                           ), //i
    .reset                  (reset                         )  //i
  );
  PEWSOS_15 pes_1_3 (
    .io_in_r_data           (pes_1_2_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pes_1_2_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pes_1_2_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pes_1_2_io_out_r_stall        ), //i
    .io_out_r_data          (pes_1_3_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pes_1_3_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pes_1_3_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pes_1_3_io_out_r_stall        ), //o
    .io_in_c_data           (pes_0_3_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pes_0_3_io_out_c_is_stationary), //i
    .io_out_c_data          (pes_1_3_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pes_1_3_io_out_c_is_stationary), //o
    .clk                    (clk                           ), //i
    .reset                  (reset                         )  //i
  );
  PEWSOS_15 pes_2_0 (
    .io_in_r_data           (in_r_2_data[15:0]             ), //i
    .io_in_r_load_store     (in_r_2_load_store             ), //i
    .io_in_r_df_is_ws       (in_r_2_df_is_ws               ), //i
    .io_in_r_stall          (in_r_2_stall                  ), //i
    .io_out_r_data          (pes_2_0_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pes_2_0_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pes_2_0_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pes_2_0_io_out_r_stall        ), //o
    .io_in_c_data           (pes_1_0_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pes_1_0_io_out_c_is_stationary), //i
    .io_out_c_data          (pes_2_0_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pes_2_0_io_out_c_is_stationary), //o
    .clk                    (clk                           ), //i
    .reset                  (reset                         )  //i
  );
  PEWSOS_15 pes_2_1 (
    .io_in_r_data           (pes_2_0_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pes_2_0_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pes_2_0_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pes_2_0_io_out_r_stall        ), //i
    .io_out_r_data          (pes_2_1_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pes_2_1_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pes_2_1_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pes_2_1_io_out_r_stall        ), //o
    .io_in_c_data           (pes_1_1_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pes_1_1_io_out_c_is_stationary), //i
    .io_out_c_data          (pes_2_1_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pes_2_1_io_out_c_is_stationary), //o
    .clk                    (clk                           ), //i
    .reset                  (reset                         )  //i
  );
  PEWSOS_15 pes_2_2 (
    .io_in_r_data           (pes_2_1_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pes_2_1_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pes_2_1_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pes_2_1_io_out_r_stall        ), //i
    .io_out_r_data          (pes_2_2_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pes_2_2_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pes_2_2_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pes_2_2_io_out_r_stall        ), //o
    .io_in_c_data           (pes_1_2_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pes_1_2_io_out_c_is_stationary), //i
    .io_out_c_data          (pes_2_2_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pes_2_2_io_out_c_is_stationary), //o
    .clk                    (clk                           ), //i
    .reset                  (reset                         )  //i
  );
  PEWSOS_15 pes_2_3 (
    .io_in_r_data           (pes_2_2_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pes_2_2_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pes_2_2_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pes_2_2_io_out_r_stall        ), //i
    .io_out_r_data          (pes_2_3_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pes_2_3_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pes_2_3_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pes_2_3_io_out_r_stall        ), //o
    .io_in_c_data           (pes_1_3_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pes_1_3_io_out_c_is_stationary), //i
    .io_out_c_data          (pes_2_3_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pes_2_3_io_out_c_is_stationary), //o
    .clk                    (clk                           ), //i
    .reset                  (reset                         )  //i
  );
  PEWSOS_15 pes_3_0 (
    .io_in_r_data           (in_r_3_data[15:0]             ), //i
    .io_in_r_load_store     (in_r_3_load_store             ), //i
    .io_in_r_df_is_ws       (in_r_3_df_is_ws               ), //i
    .io_in_r_stall          (in_r_3_stall                  ), //i
    .io_out_r_data          (pes_3_0_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pes_3_0_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pes_3_0_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pes_3_0_io_out_r_stall        ), //o
    .io_in_c_data           (pes_2_0_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pes_2_0_io_out_c_is_stationary), //i
    .io_out_c_data          (pes_3_0_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pes_3_0_io_out_c_is_stationary), //o
    .clk                    (clk                           ), //i
    .reset                  (reset                         )  //i
  );
  PEWSOS_15 pes_3_1 (
    .io_in_r_data           (pes_3_0_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pes_3_0_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pes_3_0_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pes_3_0_io_out_r_stall        ), //i
    .io_out_r_data          (pes_3_1_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pes_3_1_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pes_3_1_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pes_3_1_io_out_r_stall        ), //o
    .io_in_c_data           (pes_2_1_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pes_2_1_io_out_c_is_stationary), //i
    .io_out_c_data          (pes_3_1_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pes_3_1_io_out_c_is_stationary), //o
    .clk                    (clk                           ), //i
    .reset                  (reset                         )  //i
  );
  PEWSOS_15 pes_3_2 (
    .io_in_r_data           (pes_3_1_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pes_3_1_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pes_3_1_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pes_3_1_io_out_r_stall        ), //i
    .io_out_r_data          (pes_3_2_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pes_3_2_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pes_3_2_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pes_3_2_io_out_r_stall        ), //o
    .io_in_c_data           (pes_2_2_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pes_2_2_io_out_c_is_stationary), //i
    .io_out_c_data          (pes_3_2_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pes_3_2_io_out_c_is_stationary), //o
    .clk                    (clk                           ), //i
    .reset                  (reset                         )  //i
  );
  PEWSOS_15 pes_3_3 (
    .io_in_r_data           (pes_3_2_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pes_3_2_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pes_3_2_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pes_3_2_io_out_r_stall        ), //i
    .io_out_r_data          (pes_3_3_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pes_3_3_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pes_3_3_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pes_3_3_io_out_r_stall        ), //o
    .io_in_c_data           (pes_2_3_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pes_2_3_io_out_c_is_stationary), //i
    .io_out_c_data          (pes_3_3_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pes_3_3_io_out_c_is_stationary), //o
    .clk                    (clk                           ), //i
    .reset                  (reset                         )  //i
  );
  assign in_r_0_data = (io_in_r_input_from_bypass_0 ? io_in_r_bypass_0_0_data : io_in_r_data_0_data); // @[Expression.scala 1420:25]
  assign in_r_0_load_store = (io_in_r_input_from_bypass_0 ? io_in_r_bypass_0_0_load_store : io_in_r_data_0_load_store); // @[Expression.scala 1420:25]
  assign in_r_0_df_is_ws = (io_in_r_input_from_bypass_0 ? io_in_r_bypass_0_0_df_is_ws : io_in_r_data_0_df_is_ws); // @[Expression.scala 1420:25]
  assign in_r_0_stall = (io_in_r_input_from_bypass_0 ? io_in_r_bypass_0_0_stall : io_in_r_data_0_stall); // @[Expression.scala 1420:25]
  assign in_r_1_data = (io_in_r_input_from_bypass_0 ? io_in_r_bypass_0_1_data : io_in_r_data_1_data); // @[Expression.scala 1420:25]
  assign in_r_1_load_store = (io_in_r_input_from_bypass_0 ? io_in_r_bypass_0_1_load_store : io_in_r_data_1_load_store); // @[Expression.scala 1420:25]
  assign in_r_1_df_is_ws = (io_in_r_input_from_bypass_0 ? io_in_r_bypass_0_1_df_is_ws : io_in_r_data_1_df_is_ws); // @[Expression.scala 1420:25]
  assign in_r_1_stall = (io_in_r_input_from_bypass_0 ? io_in_r_bypass_0_1_stall : io_in_r_data_1_stall); // @[Expression.scala 1420:25]
  assign in_r_2_data = (io_in_r_input_from_bypass_0 ? io_in_r_bypass_0_2_data : io_in_r_data_2_data); // @[Expression.scala 1420:25]
  assign in_r_2_load_store = (io_in_r_input_from_bypass_0 ? io_in_r_bypass_0_2_load_store : io_in_r_data_2_load_store); // @[Expression.scala 1420:25]
  assign in_r_2_df_is_ws = (io_in_r_input_from_bypass_0 ? io_in_r_bypass_0_2_df_is_ws : io_in_r_data_2_df_is_ws); // @[Expression.scala 1420:25]
  assign in_r_2_stall = (io_in_r_input_from_bypass_0 ? io_in_r_bypass_0_2_stall : io_in_r_data_2_stall); // @[Expression.scala 1420:25]
  assign in_r_3_data = (io_in_r_input_from_bypass_0 ? io_in_r_bypass_0_3_data : io_in_r_data_3_data); // @[Expression.scala 1420:25]
  assign in_r_3_load_store = (io_in_r_input_from_bypass_0 ? io_in_r_bypass_0_3_load_store : io_in_r_data_3_load_store); // @[Expression.scala 1420:25]
  assign in_r_3_df_is_ws = (io_in_r_input_from_bypass_0 ? io_in_r_bypass_0_3_df_is_ws : io_in_r_data_3_df_is_ws); // @[Expression.scala 1420:25]
  assign in_r_3_stall = (io_in_r_input_from_bypass_0 ? io_in_r_bypass_0_3_stall : io_in_r_data_3_stall); // @[Expression.scala 1420:25]
  assign in_c_0_data = (io_in_c_input_from_bypass_0 ? io_in_c_bypass_0_0_data : io_in_c_data_0_data); // @[Expression.scala 1420:25]
  assign in_c_0_is_stationary = (io_in_c_input_from_bypass_0 ? io_in_c_bypass_0_0_is_stationary : io_in_c_data_0_is_stationary); // @[Expression.scala 1420:25]
  assign in_c_1_data = (io_in_c_input_from_bypass_0 ? io_in_c_bypass_0_1_data : io_in_c_data_1_data); // @[Expression.scala 1420:25]
  assign in_c_1_is_stationary = (io_in_c_input_from_bypass_0 ? io_in_c_bypass_0_1_is_stationary : io_in_c_data_1_is_stationary); // @[Expression.scala 1420:25]
  assign in_c_2_data = (io_in_c_input_from_bypass_0 ? io_in_c_bypass_0_2_data : io_in_c_data_2_data); // @[Expression.scala 1420:25]
  assign in_c_2_is_stationary = (io_in_c_input_from_bypass_0 ? io_in_c_bypass_0_2_is_stationary : io_in_c_data_2_is_stationary); // @[Expression.scala 1420:25]
  assign in_c_3_data = (io_in_c_input_from_bypass_0 ? io_in_c_bypass_0_3_data : io_in_c_data_3_data); // @[Expression.scala 1420:25]
  assign in_c_3_is_stationary = (io_in_c_input_from_bypass_0 ? io_in_c_bypass_0_3_is_stationary : io_in_c_data_3_is_stationary); // @[Expression.scala 1420:25]
  assign out_r_0_data = pes_0_3_io_out_r_data; // @[SystolicConnect.scala 50:16]
  assign out_r_0_load_store = pes_0_3_io_out_r_load_store; // @[SystolicConnect.scala 50:16]
  assign out_r_0_df_is_ws = pes_0_3_io_out_r_df_is_ws; // @[SystolicConnect.scala 50:16]
  assign out_r_0_stall = pes_0_3_io_out_r_stall; // @[SystolicConnect.scala 50:16]
  assign out_r_1_data = pes_1_3_io_out_r_data; // @[SystolicConnect.scala 50:16]
  assign out_r_1_load_store = pes_1_3_io_out_r_load_store; // @[SystolicConnect.scala 50:16]
  assign out_r_1_df_is_ws = pes_1_3_io_out_r_df_is_ws; // @[SystolicConnect.scala 50:16]
  assign out_r_1_stall = pes_1_3_io_out_r_stall; // @[SystolicConnect.scala 50:16]
  assign out_r_2_data = pes_2_3_io_out_r_data; // @[SystolicConnect.scala 50:16]
  assign out_r_2_load_store = pes_2_3_io_out_r_load_store; // @[SystolicConnect.scala 50:16]
  assign out_r_2_df_is_ws = pes_2_3_io_out_r_df_is_ws; // @[SystolicConnect.scala 50:16]
  assign out_r_2_stall = pes_2_3_io_out_r_stall; // @[SystolicConnect.scala 50:16]
  assign out_r_3_data = pes_3_3_io_out_r_data; // @[SystolicConnect.scala 50:16]
  assign out_r_3_load_store = pes_3_3_io_out_r_load_store; // @[SystolicConnect.scala 50:16]
  assign out_r_3_df_is_ws = pes_3_3_io_out_r_df_is_ws; // @[SystolicConnect.scala 50:16]
  assign out_r_3_stall = pes_3_3_io_out_r_stall; // @[SystolicConnect.scala 50:16]
  assign out_c_0_data = pes_3_0_io_out_c_data; // @[SystolicConnect.scala 56:16]
  assign out_c_0_is_stationary = pes_3_0_io_out_c_is_stationary; // @[SystolicConnect.scala 56:16]
  assign out_c_1_data = pes_3_1_io_out_c_data; // @[SystolicConnect.scala 56:16]
  assign out_c_1_is_stationary = pes_3_1_io_out_c_is_stationary; // @[SystolicConnect.scala 56:16]
  assign out_c_2_data = pes_3_2_io_out_c_data; // @[SystolicConnect.scala 56:16]
  assign out_c_2_is_stationary = pes_3_2_io_out_c_is_stationary; // @[SystolicConnect.scala 56:16]
  assign out_c_3_data = pes_3_3_io_out_c_data; // @[SystolicConnect.scala 56:16]
  assign out_c_3_is_stationary = pes_3_3_io_out_c_is_stationary; // @[SystolicConnect.scala 56:16]
  assign io_out_r_data_0_data = out_r_0_data; // @[ArraySARA.scala 90:17]
  assign io_out_r_data_0_load_store = out_r_0_load_store; // @[ArraySARA.scala 90:17]
  assign io_out_r_data_0_df_is_ws = out_r_0_df_is_ws; // @[ArraySARA.scala 90:17]
  assign io_out_r_data_0_stall = out_r_0_stall; // @[ArraySARA.scala 90:17]
  assign io_out_r_data_1_data = out_r_1_data; // @[ArraySARA.scala 90:17]
  assign io_out_r_data_1_load_store = out_r_1_load_store; // @[ArraySARA.scala 90:17]
  assign io_out_r_data_1_df_is_ws = out_r_1_df_is_ws; // @[ArraySARA.scala 90:17]
  assign io_out_r_data_1_stall = out_r_1_stall; // @[ArraySARA.scala 90:17]
  assign io_out_r_data_2_data = out_r_2_data; // @[ArraySARA.scala 90:17]
  assign io_out_r_data_2_load_store = out_r_2_load_store; // @[ArraySARA.scala 90:17]
  assign io_out_r_data_2_df_is_ws = out_r_2_df_is_ws; // @[ArraySARA.scala 90:17]
  assign io_out_r_data_2_stall = out_r_2_stall; // @[ArraySARA.scala 90:17]
  assign io_out_r_data_3_data = out_r_3_data; // @[ArraySARA.scala 90:17]
  assign io_out_r_data_3_load_store = out_r_3_load_store; // @[ArraySARA.scala 90:17]
  assign io_out_r_data_3_df_is_ws = out_r_3_df_is_ws; // @[ArraySARA.scala 90:17]
  assign io_out_r_data_3_stall = out_r_3_stall; // @[ArraySARA.scala 90:17]
  assign io_out_c_data_0_data = out_c_0_data; // @[ArraySARA.scala 91:17]
  assign io_out_c_data_0_is_stationary = out_c_0_is_stationary; // @[ArraySARA.scala 91:17]
  assign io_out_c_data_1_data = out_c_1_data; // @[ArraySARA.scala 91:17]
  assign io_out_c_data_1_is_stationary = out_c_1_is_stationary; // @[ArraySARA.scala 91:17]
  assign io_out_c_data_2_data = out_c_2_data; // @[ArraySARA.scala 91:17]
  assign io_out_c_data_2_is_stationary = out_c_2_is_stationary; // @[ArraySARA.scala 91:17]
  assign io_out_c_data_3_data = out_c_3_data; // @[ArraySARA.scala 91:17]
  assign io_out_c_data_3_is_stationary = out_c_3_is_stationary; // @[ArraySARA.scala 91:17]
  assign io_out_r_bypass_0_0_data = out_r_regNext_0_data; // @[ArraySARA.scala 92:31]
  assign io_out_r_bypass_0_0_load_store = out_r_regNext_0_load_store; // @[ArraySARA.scala 92:31]
  assign io_out_r_bypass_0_0_df_is_ws = out_r_regNext_0_df_is_ws; // @[ArraySARA.scala 92:31]
  assign io_out_r_bypass_0_0_stall = out_r_regNext_0_stall; // @[ArraySARA.scala 92:31]
  assign io_out_r_bypass_0_1_data = out_r_regNext_1_data; // @[ArraySARA.scala 92:31]
  assign io_out_r_bypass_0_1_load_store = out_r_regNext_1_load_store; // @[ArraySARA.scala 92:31]
  assign io_out_r_bypass_0_1_df_is_ws = out_r_regNext_1_df_is_ws; // @[ArraySARA.scala 92:31]
  assign io_out_r_bypass_0_1_stall = out_r_regNext_1_stall; // @[ArraySARA.scala 92:31]
  assign io_out_r_bypass_0_2_data = out_r_regNext_2_data; // @[ArraySARA.scala 92:31]
  assign io_out_r_bypass_0_2_load_store = out_r_regNext_2_load_store; // @[ArraySARA.scala 92:31]
  assign io_out_r_bypass_0_2_df_is_ws = out_r_regNext_2_df_is_ws; // @[ArraySARA.scala 92:31]
  assign io_out_r_bypass_0_2_stall = out_r_regNext_2_stall; // @[ArraySARA.scala 92:31]
  assign io_out_r_bypass_0_3_data = out_r_regNext_3_data; // @[ArraySARA.scala 92:31]
  assign io_out_r_bypass_0_3_load_store = out_r_regNext_3_load_store; // @[ArraySARA.scala 92:31]
  assign io_out_r_bypass_0_3_df_is_ws = out_r_regNext_3_df_is_ws; // @[ArraySARA.scala 92:31]
  assign io_out_r_bypass_0_3_stall = out_r_regNext_3_stall; // @[ArraySARA.scala 92:31]
  assign io_out_c_bypass_0_0_data = out_c_regNext_0_data; // @[ArraySARA.scala 93:31]
  assign io_out_c_bypass_0_0_is_stationary = out_c_regNext_0_is_stationary; // @[ArraySARA.scala 93:31]
  assign io_out_c_bypass_0_1_data = out_c_regNext_1_data; // @[ArraySARA.scala 93:31]
  assign io_out_c_bypass_0_1_is_stationary = out_c_regNext_1_is_stationary; // @[ArraySARA.scala 93:31]
  assign io_out_c_bypass_0_2_data = out_c_regNext_2_data; // @[ArraySARA.scala 93:31]
  assign io_out_c_bypass_0_2_is_stationary = out_c_regNext_2_is_stationary; // @[ArraySARA.scala 93:31]
  assign io_out_c_bypass_0_3_data = out_c_regNext_3_data; // @[ArraySARA.scala 93:31]
  assign io_out_c_bypass_0_3_is_stationary = out_c_regNext_3_is_stationary; // @[ArraySARA.scala 93:31]
  assign io_out_r_bypass_1_0_data = io_in_r_bypass_regNext_1_0_data; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_1_0_load_store = io_in_r_bypass_regNext_1_0_load_store; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_1_0_df_is_ws = io_in_r_bypass_regNext_1_0_df_is_ws; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_1_0_stall = io_in_r_bypass_regNext_1_0_stall; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_1_1_data = io_in_r_bypass_regNext_1_1_data; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_1_1_load_store = io_in_r_bypass_regNext_1_1_load_store; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_1_1_df_is_ws = io_in_r_bypass_regNext_1_1_df_is_ws; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_1_1_stall = io_in_r_bypass_regNext_1_1_stall; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_1_2_data = io_in_r_bypass_regNext_1_2_data; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_1_2_load_store = io_in_r_bypass_regNext_1_2_load_store; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_1_2_df_is_ws = io_in_r_bypass_regNext_1_2_df_is_ws; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_1_2_stall = io_in_r_bypass_regNext_1_2_stall; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_1_3_data = io_in_r_bypass_regNext_1_3_data; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_1_3_load_store = io_in_r_bypass_regNext_1_3_load_store; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_1_3_df_is_ws = io_in_r_bypass_regNext_1_3_df_is_ws; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_1_3_stall = io_in_r_bypass_regNext_1_3_stall; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_2_0_data = io_in_r_bypass_regNext_2_0_data_1; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_2_0_load_store = io_in_r_bypass_regNext_2_0_load_store_1; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_2_0_df_is_ws = io_in_r_bypass_regNext_2_0_df_is_ws_1; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_2_0_stall = io_in_r_bypass_regNext_2_0_stall_1; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_2_1_data = io_in_r_bypass_regNext_2_1_data_1; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_2_1_load_store = io_in_r_bypass_regNext_2_1_load_store_1; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_2_1_df_is_ws = io_in_r_bypass_regNext_2_1_df_is_ws_1; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_2_1_stall = io_in_r_bypass_regNext_2_1_stall_1; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_2_2_data = io_in_r_bypass_regNext_2_2_data_1; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_2_2_load_store = io_in_r_bypass_regNext_2_2_load_store_1; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_2_2_df_is_ws = io_in_r_bypass_regNext_2_2_df_is_ws_1; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_2_2_stall = io_in_r_bypass_regNext_2_2_stall_1; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_2_3_data = io_in_r_bypass_regNext_2_3_data_1; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_2_3_load_store = io_in_r_bypass_regNext_2_3_load_store_1; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_2_3_df_is_ws = io_in_r_bypass_regNext_2_3_df_is_ws_1; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_2_3_stall = io_in_r_bypass_regNext_2_3_stall_1; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_3_0_data = io_in_r_bypass_regNext_3_0_data_2; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_3_0_load_store = io_in_r_bypass_regNext_3_0_load_store_2; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_3_0_df_is_ws = io_in_r_bypass_regNext_3_0_df_is_ws_2; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_3_0_stall = io_in_r_bypass_regNext_3_0_stall_2; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_3_1_data = io_in_r_bypass_regNext_3_1_data_2; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_3_1_load_store = io_in_r_bypass_regNext_3_1_load_store_2; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_3_1_df_is_ws = io_in_r_bypass_regNext_3_1_df_is_ws_2; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_3_1_stall = io_in_r_bypass_regNext_3_1_stall_2; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_3_2_data = io_in_r_bypass_regNext_3_2_data_2; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_3_2_load_store = io_in_r_bypass_regNext_3_2_load_store_2; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_3_2_df_is_ws = io_in_r_bypass_regNext_3_2_df_is_ws_2; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_3_2_stall = io_in_r_bypass_regNext_3_2_stall_2; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_3_3_data = io_in_r_bypass_regNext_3_3_data_2; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_3_3_load_store = io_in_r_bypass_regNext_3_3_load_store_2; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_3_3_df_is_ws = io_in_r_bypass_regNext_3_3_df_is_ws_2; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_3_3_stall = io_in_r_bypass_regNext_3_3_stall_2; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_4_0_data = io_in_r_bypass_regNext_4_0_data_3; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_4_0_load_store = io_in_r_bypass_regNext_4_0_load_store_3; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_4_0_df_is_ws = io_in_r_bypass_regNext_4_0_df_is_ws_3; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_4_0_stall = io_in_r_bypass_regNext_4_0_stall_3; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_4_1_data = io_in_r_bypass_regNext_4_1_data_3; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_4_1_load_store = io_in_r_bypass_regNext_4_1_load_store_3; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_4_1_df_is_ws = io_in_r_bypass_regNext_4_1_df_is_ws_3; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_4_1_stall = io_in_r_bypass_regNext_4_1_stall_3; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_4_2_data = io_in_r_bypass_regNext_4_2_data_3; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_4_2_load_store = io_in_r_bypass_regNext_4_2_load_store_3; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_4_2_df_is_ws = io_in_r_bypass_regNext_4_2_df_is_ws_3; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_4_2_stall = io_in_r_bypass_regNext_4_2_stall_3; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_4_3_data = io_in_r_bypass_regNext_4_3_data_3; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_4_3_load_store = io_in_r_bypass_regNext_4_3_load_store_3; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_4_3_df_is_ws = io_in_r_bypass_regNext_4_3_df_is_ws_3; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_4_3_stall = io_in_r_bypass_regNext_4_3_stall_3; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_5_0_data = io_in_r_bypass_regNext_5_0_data_4; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_5_0_load_store = io_in_r_bypass_regNext_5_0_load_store_4; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_5_0_df_is_ws = io_in_r_bypass_regNext_5_0_df_is_ws_4; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_5_0_stall = io_in_r_bypass_regNext_5_0_stall_4; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_5_1_data = io_in_r_bypass_regNext_5_1_data_4; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_5_1_load_store = io_in_r_bypass_regNext_5_1_load_store_4; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_5_1_df_is_ws = io_in_r_bypass_regNext_5_1_df_is_ws_4; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_5_1_stall = io_in_r_bypass_regNext_5_1_stall_4; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_5_2_data = io_in_r_bypass_regNext_5_2_data_4; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_5_2_load_store = io_in_r_bypass_regNext_5_2_load_store_4; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_5_2_df_is_ws = io_in_r_bypass_regNext_5_2_df_is_ws_4; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_5_2_stall = io_in_r_bypass_regNext_5_2_stall_4; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_5_3_data = io_in_r_bypass_regNext_5_3_data_4; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_5_3_load_store = io_in_r_bypass_regNext_5_3_load_store_4; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_5_3_df_is_ws = io_in_r_bypass_regNext_5_3_df_is_ws_4; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_5_3_stall = io_in_r_bypass_regNext_5_3_stall_4; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_6_0_data = io_in_r_bypass_regNext_6_0_data_5; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_6_0_load_store = io_in_r_bypass_regNext_6_0_load_store_5; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_6_0_df_is_ws = io_in_r_bypass_regNext_6_0_df_is_ws_5; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_6_0_stall = io_in_r_bypass_regNext_6_0_stall_5; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_6_1_data = io_in_r_bypass_regNext_6_1_data_5; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_6_1_load_store = io_in_r_bypass_regNext_6_1_load_store_5; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_6_1_df_is_ws = io_in_r_bypass_regNext_6_1_df_is_ws_5; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_6_1_stall = io_in_r_bypass_regNext_6_1_stall_5; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_6_2_data = io_in_r_bypass_regNext_6_2_data_5; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_6_2_load_store = io_in_r_bypass_regNext_6_2_load_store_5; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_6_2_df_is_ws = io_in_r_bypass_regNext_6_2_df_is_ws_5; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_6_2_stall = io_in_r_bypass_regNext_6_2_stall_5; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_6_3_data = io_in_r_bypass_regNext_6_3_data_5; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_6_3_load_store = io_in_r_bypass_regNext_6_3_load_store_5; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_6_3_df_is_ws = io_in_r_bypass_regNext_6_3_df_is_ws_5; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_6_3_stall = io_in_r_bypass_regNext_6_3_stall_5; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_7_0_data = io_in_r_bypass_regNext_7_0_data_6; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_7_0_load_store = io_in_r_bypass_regNext_7_0_load_store_6; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_7_0_df_is_ws = io_in_r_bypass_regNext_7_0_df_is_ws_6; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_7_0_stall = io_in_r_bypass_regNext_7_0_stall_6; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_7_1_data = io_in_r_bypass_regNext_7_1_data_6; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_7_1_load_store = io_in_r_bypass_regNext_7_1_load_store_6; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_7_1_df_is_ws = io_in_r_bypass_regNext_7_1_df_is_ws_6; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_7_1_stall = io_in_r_bypass_regNext_7_1_stall_6; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_7_2_data = io_in_r_bypass_regNext_7_2_data_6; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_7_2_load_store = io_in_r_bypass_regNext_7_2_load_store_6; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_7_2_df_is_ws = io_in_r_bypass_regNext_7_2_df_is_ws_6; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_7_2_stall = io_in_r_bypass_regNext_7_2_stall_6; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_7_3_data = io_in_r_bypass_regNext_7_3_data_6; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_7_3_load_store = io_in_r_bypass_regNext_7_3_load_store_6; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_7_3_df_is_ws = io_in_r_bypass_regNext_7_3_df_is_ws_6; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_7_3_stall = io_in_r_bypass_regNext_7_3_stall_6; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_8_0_data = io_in_r_bypass_regNext_8_0_data_7; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_8_0_load_store = io_in_r_bypass_regNext_8_0_load_store_7; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_8_0_df_is_ws = io_in_r_bypass_regNext_8_0_df_is_ws_7; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_8_0_stall = io_in_r_bypass_regNext_8_0_stall_7; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_8_1_data = io_in_r_bypass_regNext_8_1_data_7; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_8_1_load_store = io_in_r_bypass_regNext_8_1_load_store_7; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_8_1_df_is_ws = io_in_r_bypass_regNext_8_1_df_is_ws_7; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_8_1_stall = io_in_r_bypass_regNext_8_1_stall_7; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_8_2_data = io_in_r_bypass_regNext_8_2_data_7; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_8_2_load_store = io_in_r_bypass_regNext_8_2_load_store_7; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_8_2_df_is_ws = io_in_r_bypass_regNext_8_2_df_is_ws_7; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_8_2_stall = io_in_r_bypass_regNext_8_2_stall_7; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_8_3_data = io_in_r_bypass_regNext_8_3_data_7; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_8_3_load_store = io_in_r_bypass_regNext_8_3_load_store_7; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_8_3_df_is_ws = io_in_r_bypass_regNext_8_3_df_is_ws_7; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_8_3_stall = io_in_r_bypass_regNext_8_3_stall_7; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_9_0_data = io_in_r_bypass_regNext_9_0_data_8; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_9_0_load_store = io_in_r_bypass_regNext_9_0_load_store_8; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_9_0_df_is_ws = io_in_r_bypass_regNext_9_0_df_is_ws_8; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_9_0_stall = io_in_r_bypass_regNext_9_0_stall_8; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_9_1_data = io_in_r_bypass_regNext_9_1_data_8; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_9_1_load_store = io_in_r_bypass_regNext_9_1_load_store_8; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_9_1_df_is_ws = io_in_r_bypass_regNext_9_1_df_is_ws_8; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_9_1_stall = io_in_r_bypass_regNext_9_1_stall_8; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_9_2_data = io_in_r_bypass_regNext_9_2_data_8; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_9_2_load_store = io_in_r_bypass_regNext_9_2_load_store_8; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_9_2_df_is_ws = io_in_r_bypass_regNext_9_2_df_is_ws_8; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_9_2_stall = io_in_r_bypass_regNext_9_2_stall_8; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_9_3_data = io_in_r_bypass_regNext_9_3_data_8; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_9_3_load_store = io_in_r_bypass_regNext_9_3_load_store_8; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_9_3_df_is_ws = io_in_r_bypass_regNext_9_3_df_is_ws_8; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_9_3_stall = io_in_r_bypass_regNext_9_3_stall_8; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_10_0_data = io_in_r_bypass_regNext_10_0_data_9; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_10_0_load_store = io_in_r_bypass_regNext_10_0_load_store_9; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_10_0_df_is_ws = io_in_r_bypass_regNext_10_0_df_is_ws_9; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_10_0_stall = io_in_r_bypass_regNext_10_0_stall_9; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_10_1_data = io_in_r_bypass_regNext_10_1_data_9; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_10_1_load_store = io_in_r_bypass_regNext_10_1_load_store_9; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_10_1_df_is_ws = io_in_r_bypass_regNext_10_1_df_is_ws_9; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_10_1_stall = io_in_r_bypass_regNext_10_1_stall_9; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_10_2_data = io_in_r_bypass_regNext_10_2_data_9; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_10_2_load_store = io_in_r_bypass_regNext_10_2_load_store_9; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_10_2_df_is_ws = io_in_r_bypass_regNext_10_2_df_is_ws_9; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_10_2_stall = io_in_r_bypass_regNext_10_2_stall_9; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_10_3_data = io_in_r_bypass_regNext_10_3_data_9; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_10_3_load_store = io_in_r_bypass_regNext_10_3_load_store_9; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_10_3_df_is_ws = io_in_r_bypass_regNext_10_3_df_is_ws_9; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_10_3_stall = io_in_r_bypass_regNext_10_3_stall_9; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_11_0_data = io_in_r_bypass_regNext_11_0_data_10; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_11_0_load_store = io_in_r_bypass_regNext_11_0_load_store_10; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_11_0_df_is_ws = io_in_r_bypass_regNext_11_0_df_is_ws_10; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_11_0_stall = io_in_r_bypass_regNext_11_0_stall_10; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_11_1_data = io_in_r_bypass_regNext_11_1_data_10; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_11_1_load_store = io_in_r_bypass_regNext_11_1_load_store_10; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_11_1_df_is_ws = io_in_r_bypass_regNext_11_1_df_is_ws_10; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_11_1_stall = io_in_r_bypass_regNext_11_1_stall_10; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_11_2_data = io_in_r_bypass_regNext_11_2_data_10; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_11_2_load_store = io_in_r_bypass_regNext_11_2_load_store_10; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_11_2_df_is_ws = io_in_r_bypass_regNext_11_2_df_is_ws_10; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_11_2_stall = io_in_r_bypass_regNext_11_2_stall_10; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_11_3_data = io_in_r_bypass_regNext_11_3_data_10; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_11_3_load_store = io_in_r_bypass_regNext_11_3_load_store_10; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_11_3_df_is_ws = io_in_r_bypass_regNext_11_3_df_is_ws_10; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_11_3_stall = io_in_r_bypass_regNext_11_3_stall_10; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_12_0_data = io_in_r_bypass_regNext_12_0_data_11; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_12_0_load_store = io_in_r_bypass_regNext_12_0_load_store_11; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_12_0_df_is_ws = io_in_r_bypass_regNext_12_0_df_is_ws_11; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_12_0_stall = io_in_r_bypass_regNext_12_0_stall_11; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_12_1_data = io_in_r_bypass_regNext_12_1_data_11; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_12_1_load_store = io_in_r_bypass_regNext_12_1_load_store_11; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_12_1_df_is_ws = io_in_r_bypass_regNext_12_1_df_is_ws_11; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_12_1_stall = io_in_r_bypass_regNext_12_1_stall_11; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_12_2_data = io_in_r_bypass_regNext_12_2_data_11; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_12_2_load_store = io_in_r_bypass_regNext_12_2_load_store_11; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_12_2_df_is_ws = io_in_r_bypass_regNext_12_2_df_is_ws_11; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_12_2_stall = io_in_r_bypass_regNext_12_2_stall_11; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_12_3_data = io_in_r_bypass_regNext_12_3_data_11; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_12_3_load_store = io_in_r_bypass_regNext_12_3_load_store_11; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_12_3_df_is_ws = io_in_r_bypass_regNext_12_3_df_is_ws_11; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_12_3_stall = io_in_r_bypass_regNext_12_3_stall_11; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_13_0_data = io_in_r_bypass_regNext_13_0_data_12; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_13_0_load_store = io_in_r_bypass_regNext_13_0_load_store_12; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_13_0_df_is_ws = io_in_r_bypass_regNext_13_0_df_is_ws_12; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_13_0_stall = io_in_r_bypass_regNext_13_0_stall_12; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_13_1_data = io_in_r_bypass_regNext_13_1_data_12; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_13_1_load_store = io_in_r_bypass_regNext_13_1_load_store_12; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_13_1_df_is_ws = io_in_r_bypass_regNext_13_1_df_is_ws_12; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_13_1_stall = io_in_r_bypass_regNext_13_1_stall_12; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_13_2_data = io_in_r_bypass_regNext_13_2_data_12; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_13_2_load_store = io_in_r_bypass_regNext_13_2_load_store_12; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_13_2_df_is_ws = io_in_r_bypass_regNext_13_2_df_is_ws_12; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_13_2_stall = io_in_r_bypass_regNext_13_2_stall_12; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_13_3_data = io_in_r_bypass_regNext_13_3_data_12; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_13_3_load_store = io_in_r_bypass_regNext_13_3_load_store_12; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_13_3_df_is_ws = io_in_r_bypass_regNext_13_3_df_is_ws_12; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_13_3_stall = io_in_r_bypass_regNext_13_3_stall_12; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_14_0_data = io_in_r_bypass_regNext_14_0_data_13; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_14_0_load_store = io_in_r_bypass_regNext_14_0_load_store_13; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_14_0_df_is_ws = io_in_r_bypass_regNext_14_0_df_is_ws_13; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_14_0_stall = io_in_r_bypass_regNext_14_0_stall_13; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_14_1_data = io_in_r_bypass_regNext_14_1_data_13; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_14_1_load_store = io_in_r_bypass_regNext_14_1_load_store_13; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_14_1_df_is_ws = io_in_r_bypass_regNext_14_1_df_is_ws_13; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_14_1_stall = io_in_r_bypass_regNext_14_1_stall_13; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_14_2_data = io_in_r_bypass_regNext_14_2_data_13; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_14_2_load_store = io_in_r_bypass_regNext_14_2_load_store_13; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_14_2_df_is_ws = io_in_r_bypass_regNext_14_2_df_is_ws_13; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_14_2_stall = io_in_r_bypass_regNext_14_2_stall_13; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_14_3_data = io_in_r_bypass_regNext_14_3_data_13; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_14_3_load_store = io_in_r_bypass_regNext_14_3_load_store_13; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_14_3_df_is_ws = io_in_r_bypass_regNext_14_3_df_is_ws_13; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_14_3_stall = io_in_r_bypass_regNext_14_3_stall_13; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_15_0_data = io_in_r_bypass_regNext_15_0_data_14; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_15_0_load_store = io_in_r_bypass_regNext_15_0_load_store_14; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_15_0_df_is_ws = io_in_r_bypass_regNext_15_0_df_is_ws_14; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_15_0_stall = io_in_r_bypass_regNext_15_0_stall_14; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_15_1_data = io_in_r_bypass_regNext_15_1_data_14; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_15_1_load_store = io_in_r_bypass_regNext_15_1_load_store_14; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_15_1_df_is_ws = io_in_r_bypass_regNext_15_1_df_is_ws_14; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_15_1_stall = io_in_r_bypass_regNext_15_1_stall_14; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_15_2_data = io_in_r_bypass_regNext_15_2_data_14; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_15_2_load_store = io_in_r_bypass_regNext_15_2_load_store_14; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_15_2_df_is_ws = io_in_r_bypass_regNext_15_2_df_is_ws_14; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_15_2_stall = io_in_r_bypass_regNext_15_2_stall_14; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_15_3_data = io_in_r_bypass_regNext_15_3_data_14; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_15_3_load_store = io_in_r_bypass_regNext_15_3_load_store_14; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_15_3_df_is_ws = io_in_r_bypass_regNext_15_3_df_is_ws_14; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_15_3_stall = io_in_r_bypass_regNext_15_3_stall_14; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_16_0_data = io_in_r_bypass_regNext_16_0_data_15; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_16_0_load_store = io_in_r_bypass_regNext_16_0_load_store_15; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_16_0_df_is_ws = io_in_r_bypass_regNext_16_0_df_is_ws_15; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_16_0_stall = io_in_r_bypass_regNext_16_0_stall_15; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_16_1_data = io_in_r_bypass_regNext_16_1_data_15; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_16_1_load_store = io_in_r_bypass_regNext_16_1_load_store_15; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_16_1_df_is_ws = io_in_r_bypass_regNext_16_1_df_is_ws_15; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_16_1_stall = io_in_r_bypass_regNext_16_1_stall_15; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_16_2_data = io_in_r_bypass_regNext_16_2_data_15; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_16_2_load_store = io_in_r_bypass_regNext_16_2_load_store_15; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_16_2_df_is_ws = io_in_r_bypass_regNext_16_2_df_is_ws_15; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_16_2_stall = io_in_r_bypass_regNext_16_2_stall_15; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_16_3_data = io_in_r_bypass_regNext_16_3_data_15; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_16_3_load_store = io_in_r_bypass_regNext_16_3_load_store_15; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_16_3_df_is_ws = io_in_r_bypass_regNext_16_3_df_is_ws_15; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_16_3_stall = io_in_r_bypass_regNext_16_3_stall_15; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_17_0_data = io_in_r_bypass_regNext_17_0_data_16; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_17_0_load_store = io_in_r_bypass_regNext_17_0_load_store_16; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_17_0_df_is_ws = io_in_r_bypass_regNext_17_0_df_is_ws_16; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_17_0_stall = io_in_r_bypass_regNext_17_0_stall_16; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_17_1_data = io_in_r_bypass_regNext_17_1_data_16; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_17_1_load_store = io_in_r_bypass_regNext_17_1_load_store_16; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_17_1_df_is_ws = io_in_r_bypass_regNext_17_1_df_is_ws_16; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_17_1_stall = io_in_r_bypass_regNext_17_1_stall_16; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_17_2_data = io_in_r_bypass_regNext_17_2_data_16; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_17_2_load_store = io_in_r_bypass_regNext_17_2_load_store_16; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_17_2_df_is_ws = io_in_r_bypass_regNext_17_2_df_is_ws_16; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_17_2_stall = io_in_r_bypass_regNext_17_2_stall_16; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_17_3_data = io_in_r_bypass_regNext_17_3_data_16; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_17_3_load_store = io_in_r_bypass_regNext_17_3_load_store_16; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_17_3_df_is_ws = io_in_r_bypass_regNext_17_3_df_is_ws_16; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_17_3_stall = io_in_r_bypass_regNext_17_3_stall_16; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_18_0_data = io_in_r_bypass_regNext_18_0_data_17; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_18_0_load_store = io_in_r_bypass_regNext_18_0_load_store_17; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_18_0_df_is_ws = io_in_r_bypass_regNext_18_0_df_is_ws_17; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_18_0_stall = io_in_r_bypass_regNext_18_0_stall_17; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_18_1_data = io_in_r_bypass_regNext_18_1_data_17; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_18_1_load_store = io_in_r_bypass_regNext_18_1_load_store_17; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_18_1_df_is_ws = io_in_r_bypass_regNext_18_1_df_is_ws_17; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_18_1_stall = io_in_r_bypass_regNext_18_1_stall_17; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_18_2_data = io_in_r_bypass_regNext_18_2_data_17; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_18_2_load_store = io_in_r_bypass_regNext_18_2_load_store_17; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_18_2_df_is_ws = io_in_r_bypass_regNext_18_2_df_is_ws_17; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_18_2_stall = io_in_r_bypass_regNext_18_2_stall_17; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_18_3_data = io_in_r_bypass_regNext_18_3_data_17; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_18_3_load_store = io_in_r_bypass_regNext_18_3_load_store_17; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_18_3_df_is_ws = io_in_r_bypass_regNext_18_3_df_is_ws_17; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_18_3_stall = io_in_r_bypass_regNext_18_3_stall_17; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_19_0_data = io_in_r_bypass_regNext_19_0_data_18; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_19_0_load_store = io_in_r_bypass_regNext_19_0_load_store_18; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_19_0_df_is_ws = io_in_r_bypass_regNext_19_0_df_is_ws_18; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_19_0_stall = io_in_r_bypass_regNext_19_0_stall_18; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_19_1_data = io_in_r_bypass_regNext_19_1_data_18; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_19_1_load_store = io_in_r_bypass_regNext_19_1_load_store_18; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_19_1_df_is_ws = io_in_r_bypass_regNext_19_1_df_is_ws_18; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_19_1_stall = io_in_r_bypass_regNext_19_1_stall_18; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_19_2_data = io_in_r_bypass_regNext_19_2_data_18; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_19_2_load_store = io_in_r_bypass_regNext_19_2_load_store_18; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_19_2_df_is_ws = io_in_r_bypass_regNext_19_2_df_is_ws_18; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_19_2_stall = io_in_r_bypass_regNext_19_2_stall_18; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_19_3_data = io_in_r_bypass_regNext_19_3_data_18; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_19_3_load_store = io_in_r_bypass_regNext_19_3_load_store_18; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_19_3_df_is_ws = io_in_r_bypass_regNext_19_3_df_is_ws_18; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_19_3_stall = io_in_r_bypass_regNext_19_3_stall_18; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_20_0_data = io_in_r_bypass_regNext_20_0_data_19; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_20_0_load_store = io_in_r_bypass_regNext_20_0_load_store_19; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_20_0_df_is_ws = io_in_r_bypass_regNext_20_0_df_is_ws_19; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_20_0_stall = io_in_r_bypass_regNext_20_0_stall_19; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_20_1_data = io_in_r_bypass_regNext_20_1_data_19; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_20_1_load_store = io_in_r_bypass_regNext_20_1_load_store_19; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_20_1_df_is_ws = io_in_r_bypass_regNext_20_1_df_is_ws_19; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_20_1_stall = io_in_r_bypass_regNext_20_1_stall_19; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_20_2_data = io_in_r_bypass_regNext_20_2_data_19; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_20_2_load_store = io_in_r_bypass_regNext_20_2_load_store_19; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_20_2_df_is_ws = io_in_r_bypass_regNext_20_2_df_is_ws_19; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_20_2_stall = io_in_r_bypass_regNext_20_2_stall_19; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_20_3_data = io_in_r_bypass_regNext_20_3_data_19; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_20_3_load_store = io_in_r_bypass_regNext_20_3_load_store_19; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_20_3_df_is_ws = io_in_r_bypass_regNext_20_3_df_is_ws_19; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_20_3_stall = io_in_r_bypass_regNext_20_3_stall_19; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_21_0_data = io_in_r_bypass_regNext_21_0_data_20; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_21_0_load_store = io_in_r_bypass_regNext_21_0_load_store_20; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_21_0_df_is_ws = io_in_r_bypass_regNext_21_0_df_is_ws_20; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_21_0_stall = io_in_r_bypass_regNext_21_0_stall_20; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_21_1_data = io_in_r_bypass_regNext_21_1_data_20; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_21_1_load_store = io_in_r_bypass_regNext_21_1_load_store_20; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_21_1_df_is_ws = io_in_r_bypass_regNext_21_1_df_is_ws_20; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_21_1_stall = io_in_r_bypass_regNext_21_1_stall_20; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_21_2_data = io_in_r_bypass_regNext_21_2_data_20; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_21_2_load_store = io_in_r_bypass_regNext_21_2_load_store_20; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_21_2_df_is_ws = io_in_r_bypass_regNext_21_2_df_is_ws_20; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_21_2_stall = io_in_r_bypass_regNext_21_2_stall_20; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_21_3_data = io_in_r_bypass_regNext_21_3_data_20; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_21_3_load_store = io_in_r_bypass_regNext_21_3_load_store_20; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_21_3_df_is_ws = io_in_r_bypass_regNext_21_3_df_is_ws_20; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_21_3_stall = io_in_r_bypass_regNext_21_3_stall_20; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_22_0_data = io_in_r_bypass_regNext_22_0_data_21; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_22_0_load_store = io_in_r_bypass_regNext_22_0_load_store_21; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_22_0_df_is_ws = io_in_r_bypass_regNext_22_0_df_is_ws_21; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_22_0_stall = io_in_r_bypass_regNext_22_0_stall_21; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_22_1_data = io_in_r_bypass_regNext_22_1_data_21; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_22_1_load_store = io_in_r_bypass_regNext_22_1_load_store_21; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_22_1_df_is_ws = io_in_r_bypass_regNext_22_1_df_is_ws_21; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_22_1_stall = io_in_r_bypass_regNext_22_1_stall_21; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_22_2_data = io_in_r_bypass_regNext_22_2_data_21; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_22_2_load_store = io_in_r_bypass_regNext_22_2_load_store_21; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_22_2_df_is_ws = io_in_r_bypass_regNext_22_2_df_is_ws_21; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_22_2_stall = io_in_r_bypass_regNext_22_2_stall_21; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_22_3_data = io_in_r_bypass_regNext_22_3_data_21; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_22_3_load_store = io_in_r_bypass_regNext_22_3_load_store_21; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_22_3_df_is_ws = io_in_r_bypass_regNext_22_3_df_is_ws_21; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_22_3_stall = io_in_r_bypass_regNext_22_3_stall_21; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_23_0_data = io_in_r_bypass_regNext_23_0_data_22; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_23_0_load_store = io_in_r_bypass_regNext_23_0_load_store_22; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_23_0_df_is_ws = io_in_r_bypass_regNext_23_0_df_is_ws_22; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_23_0_stall = io_in_r_bypass_regNext_23_0_stall_22; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_23_1_data = io_in_r_bypass_regNext_23_1_data_22; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_23_1_load_store = io_in_r_bypass_regNext_23_1_load_store_22; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_23_1_df_is_ws = io_in_r_bypass_regNext_23_1_df_is_ws_22; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_23_1_stall = io_in_r_bypass_regNext_23_1_stall_22; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_23_2_data = io_in_r_bypass_regNext_23_2_data_22; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_23_2_load_store = io_in_r_bypass_regNext_23_2_load_store_22; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_23_2_df_is_ws = io_in_r_bypass_regNext_23_2_df_is_ws_22; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_23_2_stall = io_in_r_bypass_regNext_23_2_stall_22; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_23_3_data = io_in_r_bypass_regNext_23_3_data_22; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_23_3_load_store = io_in_r_bypass_regNext_23_3_load_store_22; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_23_3_df_is_ws = io_in_r_bypass_regNext_23_3_df_is_ws_22; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_23_3_stall = io_in_r_bypass_regNext_23_3_stall_22; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_24_0_data = io_in_r_bypass_regNext_24_0_data_23; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_24_0_load_store = io_in_r_bypass_regNext_24_0_load_store_23; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_24_0_df_is_ws = io_in_r_bypass_regNext_24_0_df_is_ws_23; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_24_0_stall = io_in_r_bypass_regNext_24_0_stall_23; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_24_1_data = io_in_r_bypass_regNext_24_1_data_23; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_24_1_load_store = io_in_r_bypass_regNext_24_1_load_store_23; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_24_1_df_is_ws = io_in_r_bypass_regNext_24_1_df_is_ws_23; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_24_1_stall = io_in_r_bypass_regNext_24_1_stall_23; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_24_2_data = io_in_r_bypass_regNext_24_2_data_23; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_24_2_load_store = io_in_r_bypass_regNext_24_2_load_store_23; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_24_2_df_is_ws = io_in_r_bypass_regNext_24_2_df_is_ws_23; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_24_2_stall = io_in_r_bypass_regNext_24_2_stall_23; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_24_3_data = io_in_r_bypass_regNext_24_3_data_23; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_24_3_load_store = io_in_r_bypass_regNext_24_3_load_store_23; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_24_3_df_is_ws = io_in_r_bypass_regNext_24_3_df_is_ws_23; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_24_3_stall = io_in_r_bypass_regNext_24_3_stall_23; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_25_0_data = io_in_r_bypass_regNext_25_0_data_24; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_25_0_load_store = io_in_r_bypass_regNext_25_0_load_store_24; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_25_0_df_is_ws = io_in_r_bypass_regNext_25_0_df_is_ws_24; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_25_0_stall = io_in_r_bypass_regNext_25_0_stall_24; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_25_1_data = io_in_r_bypass_regNext_25_1_data_24; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_25_1_load_store = io_in_r_bypass_regNext_25_1_load_store_24; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_25_1_df_is_ws = io_in_r_bypass_regNext_25_1_df_is_ws_24; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_25_1_stall = io_in_r_bypass_regNext_25_1_stall_24; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_25_2_data = io_in_r_bypass_regNext_25_2_data_24; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_25_2_load_store = io_in_r_bypass_regNext_25_2_load_store_24; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_25_2_df_is_ws = io_in_r_bypass_regNext_25_2_df_is_ws_24; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_25_2_stall = io_in_r_bypass_regNext_25_2_stall_24; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_25_3_data = io_in_r_bypass_regNext_25_3_data_24; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_25_3_load_store = io_in_r_bypass_regNext_25_3_load_store_24; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_25_3_df_is_ws = io_in_r_bypass_regNext_25_3_df_is_ws_24; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_25_3_stall = io_in_r_bypass_regNext_25_3_stall_24; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_26_0_data = io_in_r_bypass_regNext_26_0_data_25; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_26_0_load_store = io_in_r_bypass_regNext_26_0_load_store_25; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_26_0_df_is_ws = io_in_r_bypass_regNext_26_0_df_is_ws_25; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_26_0_stall = io_in_r_bypass_regNext_26_0_stall_25; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_26_1_data = io_in_r_bypass_regNext_26_1_data_25; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_26_1_load_store = io_in_r_bypass_regNext_26_1_load_store_25; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_26_1_df_is_ws = io_in_r_bypass_regNext_26_1_df_is_ws_25; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_26_1_stall = io_in_r_bypass_regNext_26_1_stall_25; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_26_2_data = io_in_r_bypass_regNext_26_2_data_25; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_26_2_load_store = io_in_r_bypass_regNext_26_2_load_store_25; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_26_2_df_is_ws = io_in_r_bypass_regNext_26_2_df_is_ws_25; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_26_2_stall = io_in_r_bypass_regNext_26_2_stall_25; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_26_3_data = io_in_r_bypass_regNext_26_3_data_25; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_26_3_load_store = io_in_r_bypass_regNext_26_3_load_store_25; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_26_3_df_is_ws = io_in_r_bypass_regNext_26_3_df_is_ws_25; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_26_3_stall = io_in_r_bypass_regNext_26_3_stall_25; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_27_0_data = io_in_r_bypass_regNext_27_0_data_26; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_27_0_load_store = io_in_r_bypass_regNext_27_0_load_store_26; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_27_0_df_is_ws = io_in_r_bypass_regNext_27_0_df_is_ws_26; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_27_0_stall = io_in_r_bypass_regNext_27_0_stall_26; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_27_1_data = io_in_r_bypass_regNext_27_1_data_26; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_27_1_load_store = io_in_r_bypass_regNext_27_1_load_store_26; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_27_1_df_is_ws = io_in_r_bypass_regNext_27_1_df_is_ws_26; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_27_1_stall = io_in_r_bypass_regNext_27_1_stall_26; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_27_2_data = io_in_r_bypass_regNext_27_2_data_26; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_27_2_load_store = io_in_r_bypass_regNext_27_2_load_store_26; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_27_2_df_is_ws = io_in_r_bypass_regNext_27_2_df_is_ws_26; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_27_2_stall = io_in_r_bypass_regNext_27_2_stall_26; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_27_3_data = io_in_r_bypass_regNext_27_3_data_26; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_27_3_load_store = io_in_r_bypass_regNext_27_3_load_store_26; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_27_3_df_is_ws = io_in_r_bypass_regNext_27_3_df_is_ws_26; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_27_3_stall = io_in_r_bypass_regNext_27_3_stall_26; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_28_0_data = io_in_r_bypass_regNext_28_0_data_27; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_28_0_load_store = io_in_r_bypass_regNext_28_0_load_store_27; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_28_0_df_is_ws = io_in_r_bypass_regNext_28_0_df_is_ws_27; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_28_0_stall = io_in_r_bypass_regNext_28_0_stall_27; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_28_1_data = io_in_r_bypass_regNext_28_1_data_27; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_28_1_load_store = io_in_r_bypass_regNext_28_1_load_store_27; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_28_1_df_is_ws = io_in_r_bypass_regNext_28_1_df_is_ws_27; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_28_1_stall = io_in_r_bypass_regNext_28_1_stall_27; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_28_2_data = io_in_r_bypass_regNext_28_2_data_27; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_28_2_load_store = io_in_r_bypass_regNext_28_2_load_store_27; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_28_2_df_is_ws = io_in_r_bypass_regNext_28_2_df_is_ws_27; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_28_2_stall = io_in_r_bypass_regNext_28_2_stall_27; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_28_3_data = io_in_r_bypass_regNext_28_3_data_27; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_28_3_load_store = io_in_r_bypass_regNext_28_3_load_store_27; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_28_3_df_is_ws = io_in_r_bypass_regNext_28_3_df_is_ws_27; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_28_3_stall = io_in_r_bypass_regNext_28_3_stall_27; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_29_0_data = io_in_r_bypass_regNext_29_0_data_28; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_29_0_load_store = io_in_r_bypass_regNext_29_0_load_store_28; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_29_0_df_is_ws = io_in_r_bypass_regNext_29_0_df_is_ws_28; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_29_0_stall = io_in_r_bypass_regNext_29_0_stall_28; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_29_1_data = io_in_r_bypass_regNext_29_1_data_28; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_29_1_load_store = io_in_r_bypass_regNext_29_1_load_store_28; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_29_1_df_is_ws = io_in_r_bypass_regNext_29_1_df_is_ws_28; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_29_1_stall = io_in_r_bypass_regNext_29_1_stall_28; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_29_2_data = io_in_r_bypass_regNext_29_2_data_28; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_29_2_load_store = io_in_r_bypass_regNext_29_2_load_store_28; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_29_2_df_is_ws = io_in_r_bypass_regNext_29_2_df_is_ws_28; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_29_2_stall = io_in_r_bypass_regNext_29_2_stall_28; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_29_3_data = io_in_r_bypass_regNext_29_3_data_28; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_29_3_load_store = io_in_r_bypass_regNext_29_3_load_store_28; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_29_3_df_is_ws = io_in_r_bypass_regNext_29_3_df_is_ws_28; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_29_3_stall = io_in_r_bypass_regNext_29_3_stall_28; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_30_0_data = io_in_r_bypass_regNext_30_0_data_29; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_30_0_load_store = io_in_r_bypass_regNext_30_0_load_store_29; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_30_0_df_is_ws = io_in_r_bypass_regNext_30_0_df_is_ws_29; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_30_0_stall = io_in_r_bypass_regNext_30_0_stall_29; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_30_1_data = io_in_r_bypass_regNext_30_1_data_29; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_30_1_load_store = io_in_r_bypass_regNext_30_1_load_store_29; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_30_1_df_is_ws = io_in_r_bypass_regNext_30_1_df_is_ws_29; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_30_1_stall = io_in_r_bypass_regNext_30_1_stall_29; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_30_2_data = io_in_r_bypass_regNext_30_2_data_29; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_30_2_load_store = io_in_r_bypass_regNext_30_2_load_store_29; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_30_2_df_is_ws = io_in_r_bypass_regNext_30_2_df_is_ws_29; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_30_2_stall = io_in_r_bypass_regNext_30_2_stall_29; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_30_3_data = io_in_r_bypass_regNext_30_3_data_29; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_30_3_load_store = io_in_r_bypass_regNext_30_3_load_store_29; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_30_3_df_is_ws = io_in_r_bypass_regNext_30_3_df_is_ws_29; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_30_3_stall = io_in_r_bypass_regNext_30_3_stall_29; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_31_0_data = io_in_r_bypass_regNext_31_0_data_30; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_31_0_load_store = io_in_r_bypass_regNext_31_0_load_store_30; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_31_0_df_is_ws = io_in_r_bypass_regNext_31_0_df_is_ws_30; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_31_0_stall = io_in_r_bypass_regNext_31_0_stall_30; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_31_1_data = io_in_r_bypass_regNext_31_1_data_30; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_31_1_load_store = io_in_r_bypass_regNext_31_1_load_store_30; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_31_1_df_is_ws = io_in_r_bypass_regNext_31_1_df_is_ws_30; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_31_1_stall = io_in_r_bypass_regNext_31_1_stall_30; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_31_2_data = io_in_r_bypass_regNext_31_2_data_30; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_31_2_load_store = io_in_r_bypass_regNext_31_2_load_store_30; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_31_2_df_is_ws = io_in_r_bypass_regNext_31_2_df_is_ws_30; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_31_2_stall = io_in_r_bypass_regNext_31_2_stall_30; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_31_3_data = io_in_r_bypass_regNext_31_3_data_30; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_31_3_load_store = io_in_r_bypass_regNext_31_3_load_store_30; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_31_3_df_is_ws = io_in_r_bypass_regNext_31_3_df_is_ws_30; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_31_3_stall = io_in_r_bypass_regNext_31_3_stall_30; // @[ArraySARA.scala 97:26]
  assign io_out_c_bypass_1_0_data = io_in_c_bypass_regNext_1_0_data; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_1_0_is_stationary = io_in_c_bypass_regNext_1_0_is_stationary; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_1_1_data = io_in_c_bypass_regNext_1_1_data; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_1_1_is_stationary = io_in_c_bypass_regNext_1_1_is_stationary; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_1_2_data = io_in_c_bypass_regNext_1_2_data; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_1_2_is_stationary = io_in_c_bypass_regNext_1_2_is_stationary; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_1_3_data = io_in_c_bypass_regNext_1_3_data; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_1_3_is_stationary = io_in_c_bypass_regNext_1_3_is_stationary; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_2_0_data = io_in_c_bypass_regNext_2_0_data_1; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_2_0_is_stationary = io_in_c_bypass_regNext_2_0_is_stationary_1; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_2_1_data = io_in_c_bypass_regNext_2_1_data_1; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_2_1_is_stationary = io_in_c_bypass_regNext_2_1_is_stationary_1; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_2_2_data = io_in_c_bypass_regNext_2_2_data_1; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_2_2_is_stationary = io_in_c_bypass_regNext_2_2_is_stationary_1; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_2_3_data = io_in_c_bypass_regNext_2_3_data_1; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_2_3_is_stationary = io_in_c_bypass_regNext_2_3_is_stationary_1; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_3_0_data = io_in_c_bypass_regNext_3_0_data_2; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_3_0_is_stationary = io_in_c_bypass_regNext_3_0_is_stationary_2; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_3_1_data = io_in_c_bypass_regNext_3_1_data_2; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_3_1_is_stationary = io_in_c_bypass_regNext_3_1_is_stationary_2; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_3_2_data = io_in_c_bypass_regNext_3_2_data_2; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_3_2_is_stationary = io_in_c_bypass_regNext_3_2_is_stationary_2; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_3_3_data = io_in_c_bypass_regNext_3_3_data_2; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_3_3_is_stationary = io_in_c_bypass_regNext_3_3_is_stationary_2; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_4_0_data = io_in_c_bypass_regNext_4_0_data_3; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_4_0_is_stationary = io_in_c_bypass_regNext_4_0_is_stationary_3; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_4_1_data = io_in_c_bypass_regNext_4_1_data_3; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_4_1_is_stationary = io_in_c_bypass_regNext_4_1_is_stationary_3; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_4_2_data = io_in_c_bypass_regNext_4_2_data_3; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_4_2_is_stationary = io_in_c_bypass_regNext_4_2_is_stationary_3; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_4_3_data = io_in_c_bypass_regNext_4_3_data_3; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_4_3_is_stationary = io_in_c_bypass_regNext_4_3_is_stationary_3; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_5_0_data = io_in_c_bypass_regNext_5_0_data_4; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_5_0_is_stationary = io_in_c_bypass_regNext_5_0_is_stationary_4; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_5_1_data = io_in_c_bypass_regNext_5_1_data_4; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_5_1_is_stationary = io_in_c_bypass_regNext_5_1_is_stationary_4; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_5_2_data = io_in_c_bypass_regNext_5_2_data_4; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_5_2_is_stationary = io_in_c_bypass_regNext_5_2_is_stationary_4; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_5_3_data = io_in_c_bypass_regNext_5_3_data_4; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_5_3_is_stationary = io_in_c_bypass_regNext_5_3_is_stationary_4; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_6_0_data = io_in_c_bypass_regNext_6_0_data_5; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_6_0_is_stationary = io_in_c_bypass_regNext_6_0_is_stationary_5; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_6_1_data = io_in_c_bypass_regNext_6_1_data_5; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_6_1_is_stationary = io_in_c_bypass_regNext_6_1_is_stationary_5; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_6_2_data = io_in_c_bypass_regNext_6_2_data_5; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_6_2_is_stationary = io_in_c_bypass_regNext_6_2_is_stationary_5; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_6_3_data = io_in_c_bypass_regNext_6_3_data_5; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_6_3_is_stationary = io_in_c_bypass_regNext_6_3_is_stationary_5; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_7_0_data = io_in_c_bypass_regNext_7_0_data_6; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_7_0_is_stationary = io_in_c_bypass_regNext_7_0_is_stationary_6; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_7_1_data = io_in_c_bypass_regNext_7_1_data_6; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_7_1_is_stationary = io_in_c_bypass_regNext_7_1_is_stationary_6; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_7_2_data = io_in_c_bypass_regNext_7_2_data_6; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_7_2_is_stationary = io_in_c_bypass_regNext_7_2_is_stationary_6; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_7_3_data = io_in_c_bypass_regNext_7_3_data_6; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_7_3_is_stationary = io_in_c_bypass_regNext_7_3_is_stationary_6; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_8_0_data = io_in_c_bypass_regNext_8_0_data_7; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_8_0_is_stationary = io_in_c_bypass_regNext_8_0_is_stationary_7; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_8_1_data = io_in_c_bypass_regNext_8_1_data_7; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_8_1_is_stationary = io_in_c_bypass_regNext_8_1_is_stationary_7; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_8_2_data = io_in_c_bypass_regNext_8_2_data_7; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_8_2_is_stationary = io_in_c_bypass_regNext_8_2_is_stationary_7; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_8_3_data = io_in_c_bypass_regNext_8_3_data_7; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_8_3_is_stationary = io_in_c_bypass_regNext_8_3_is_stationary_7; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_9_0_data = io_in_c_bypass_regNext_9_0_data_8; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_9_0_is_stationary = io_in_c_bypass_regNext_9_0_is_stationary_8; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_9_1_data = io_in_c_bypass_regNext_9_1_data_8; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_9_1_is_stationary = io_in_c_bypass_regNext_9_1_is_stationary_8; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_9_2_data = io_in_c_bypass_regNext_9_2_data_8; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_9_2_is_stationary = io_in_c_bypass_regNext_9_2_is_stationary_8; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_9_3_data = io_in_c_bypass_regNext_9_3_data_8; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_9_3_is_stationary = io_in_c_bypass_regNext_9_3_is_stationary_8; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_10_0_data = io_in_c_bypass_regNext_10_0_data_9; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_10_0_is_stationary = io_in_c_bypass_regNext_10_0_is_stationary_9; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_10_1_data = io_in_c_bypass_regNext_10_1_data_9; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_10_1_is_stationary = io_in_c_bypass_regNext_10_1_is_stationary_9; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_10_2_data = io_in_c_bypass_regNext_10_2_data_9; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_10_2_is_stationary = io_in_c_bypass_regNext_10_2_is_stationary_9; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_10_3_data = io_in_c_bypass_regNext_10_3_data_9; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_10_3_is_stationary = io_in_c_bypass_regNext_10_3_is_stationary_9; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_11_0_data = io_in_c_bypass_regNext_11_0_data_10; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_11_0_is_stationary = io_in_c_bypass_regNext_11_0_is_stationary_10; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_11_1_data = io_in_c_bypass_regNext_11_1_data_10; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_11_1_is_stationary = io_in_c_bypass_regNext_11_1_is_stationary_10; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_11_2_data = io_in_c_bypass_regNext_11_2_data_10; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_11_2_is_stationary = io_in_c_bypass_regNext_11_2_is_stationary_10; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_11_3_data = io_in_c_bypass_regNext_11_3_data_10; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_11_3_is_stationary = io_in_c_bypass_regNext_11_3_is_stationary_10; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_12_0_data = io_in_c_bypass_regNext_12_0_data_11; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_12_0_is_stationary = io_in_c_bypass_regNext_12_0_is_stationary_11; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_12_1_data = io_in_c_bypass_regNext_12_1_data_11; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_12_1_is_stationary = io_in_c_bypass_regNext_12_1_is_stationary_11; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_12_2_data = io_in_c_bypass_regNext_12_2_data_11; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_12_2_is_stationary = io_in_c_bypass_regNext_12_2_is_stationary_11; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_12_3_data = io_in_c_bypass_regNext_12_3_data_11; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_12_3_is_stationary = io_in_c_bypass_regNext_12_3_is_stationary_11; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_13_0_data = io_in_c_bypass_regNext_13_0_data_12; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_13_0_is_stationary = io_in_c_bypass_regNext_13_0_is_stationary_12; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_13_1_data = io_in_c_bypass_regNext_13_1_data_12; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_13_1_is_stationary = io_in_c_bypass_regNext_13_1_is_stationary_12; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_13_2_data = io_in_c_bypass_regNext_13_2_data_12; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_13_2_is_stationary = io_in_c_bypass_regNext_13_2_is_stationary_12; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_13_3_data = io_in_c_bypass_regNext_13_3_data_12; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_13_3_is_stationary = io_in_c_bypass_regNext_13_3_is_stationary_12; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_14_0_data = io_in_c_bypass_regNext_14_0_data_13; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_14_0_is_stationary = io_in_c_bypass_regNext_14_0_is_stationary_13; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_14_1_data = io_in_c_bypass_regNext_14_1_data_13; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_14_1_is_stationary = io_in_c_bypass_regNext_14_1_is_stationary_13; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_14_2_data = io_in_c_bypass_regNext_14_2_data_13; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_14_2_is_stationary = io_in_c_bypass_regNext_14_2_is_stationary_13; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_14_3_data = io_in_c_bypass_regNext_14_3_data_13; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_14_3_is_stationary = io_in_c_bypass_regNext_14_3_is_stationary_13; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_15_0_data = io_in_c_bypass_regNext_15_0_data_14; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_15_0_is_stationary = io_in_c_bypass_regNext_15_0_is_stationary_14; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_15_1_data = io_in_c_bypass_regNext_15_1_data_14; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_15_1_is_stationary = io_in_c_bypass_regNext_15_1_is_stationary_14; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_15_2_data = io_in_c_bypass_regNext_15_2_data_14; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_15_2_is_stationary = io_in_c_bypass_regNext_15_2_is_stationary_14; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_15_3_data = io_in_c_bypass_regNext_15_3_data_14; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_15_3_is_stationary = io_in_c_bypass_regNext_15_3_is_stationary_14; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_16_0_data = io_in_c_bypass_regNext_16_0_data_15; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_16_0_is_stationary = io_in_c_bypass_regNext_16_0_is_stationary_15; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_16_1_data = io_in_c_bypass_regNext_16_1_data_15; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_16_1_is_stationary = io_in_c_bypass_regNext_16_1_is_stationary_15; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_16_2_data = io_in_c_bypass_regNext_16_2_data_15; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_16_2_is_stationary = io_in_c_bypass_regNext_16_2_is_stationary_15; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_16_3_data = io_in_c_bypass_regNext_16_3_data_15; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_16_3_is_stationary = io_in_c_bypass_regNext_16_3_is_stationary_15; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_17_0_data = io_in_c_bypass_regNext_17_0_data_16; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_17_0_is_stationary = io_in_c_bypass_regNext_17_0_is_stationary_16; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_17_1_data = io_in_c_bypass_regNext_17_1_data_16; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_17_1_is_stationary = io_in_c_bypass_regNext_17_1_is_stationary_16; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_17_2_data = io_in_c_bypass_regNext_17_2_data_16; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_17_2_is_stationary = io_in_c_bypass_regNext_17_2_is_stationary_16; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_17_3_data = io_in_c_bypass_regNext_17_3_data_16; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_17_3_is_stationary = io_in_c_bypass_regNext_17_3_is_stationary_16; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_18_0_data = io_in_c_bypass_regNext_18_0_data_17; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_18_0_is_stationary = io_in_c_bypass_regNext_18_0_is_stationary_17; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_18_1_data = io_in_c_bypass_regNext_18_1_data_17; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_18_1_is_stationary = io_in_c_bypass_regNext_18_1_is_stationary_17; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_18_2_data = io_in_c_bypass_regNext_18_2_data_17; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_18_2_is_stationary = io_in_c_bypass_regNext_18_2_is_stationary_17; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_18_3_data = io_in_c_bypass_regNext_18_3_data_17; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_18_3_is_stationary = io_in_c_bypass_regNext_18_3_is_stationary_17; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_19_0_data = io_in_c_bypass_regNext_19_0_data_18; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_19_0_is_stationary = io_in_c_bypass_regNext_19_0_is_stationary_18; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_19_1_data = io_in_c_bypass_regNext_19_1_data_18; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_19_1_is_stationary = io_in_c_bypass_regNext_19_1_is_stationary_18; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_19_2_data = io_in_c_bypass_regNext_19_2_data_18; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_19_2_is_stationary = io_in_c_bypass_regNext_19_2_is_stationary_18; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_19_3_data = io_in_c_bypass_regNext_19_3_data_18; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_19_3_is_stationary = io_in_c_bypass_regNext_19_3_is_stationary_18; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_20_0_data = io_in_c_bypass_regNext_20_0_data_19; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_20_0_is_stationary = io_in_c_bypass_regNext_20_0_is_stationary_19; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_20_1_data = io_in_c_bypass_regNext_20_1_data_19; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_20_1_is_stationary = io_in_c_bypass_regNext_20_1_is_stationary_19; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_20_2_data = io_in_c_bypass_regNext_20_2_data_19; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_20_2_is_stationary = io_in_c_bypass_regNext_20_2_is_stationary_19; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_20_3_data = io_in_c_bypass_regNext_20_3_data_19; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_20_3_is_stationary = io_in_c_bypass_regNext_20_3_is_stationary_19; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_21_0_data = io_in_c_bypass_regNext_21_0_data_20; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_21_0_is_stationary = io_in_c_bypass_regNext_21_0_is_stationary_20; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_21_1_data = io_in_c_bypass_regNext_21_1_data_20; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_21_1_is_stationary = io_in_c_bypass_regNext_21_1_is_stationary_20; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_21_2_data = io_in_c_bypass_regNext_21_2_data_20; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_21_2_is_stationary = io_in_c_bypass_regNext_21_2_is_stationary_20; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_21_3_data = io_in_c_bypass_regNext_21_3_data_20; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_21_3_is_stationary = io_in_c_bypass_regNext_21_3_is_stationary_20; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_22_0_data = io_in_c_bypass_regNext_22_0_data_21; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_22_0_is_stationary = io_in_c_bypass_regNext_22_0_is_stationary_21; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_22_1_data = io_in_c_bypass_regNext_22_1_data_21; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_22_1_is_stationary = io_in_c_bypass_regNext_22_1_is_stationary_21; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_22_2_data = io_in_c_bypass_regNext_22_2_data_21; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_22_2_is_stationary = io_in_c_bypass_regNext_22_2_is_stationary_21; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_22_3_data = io_in_c_bypass_regNext_22_3_data_21; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_22_3_is_stationary = io_in_c_bypass_regNext_22_3_is_stationary_21; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_23_0_data = io_in_c_bypass_regNext_23_0_data_22; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_23_0_is_stationary = io_in_c_bypass_regNext_23_0_is_stationary_22; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_23_1_data = io_in_c_bypass_regNext_23_1_data_22; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_23_1_is_stationary = io_in_c_bypass_regNext_23_1_is_stationary_22; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_23_2_data = io_in_c_bypass_regNext_23_2_data_22; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_23_2_is_stationary = io_in_c_bypass_regNext_23_2_is_stationary_22; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_23_3_data = io_in_c_bypass_regNext_23_3_data_22; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_23_3_is_stationary = io_in_c_bypass_regNext_23_3_is_stationary_22; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_24_0_data = io_in_c_bypass_regNext_24_0_data_23; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_24_0_is_stationary = io_in_c_bypass_regNext_24_0_is_stationary_23; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_24_1_data = io_in_c_bypass_regNext_24_1_data_23; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_24_1_is_stationary = io_in_c_bypass_regNext_24_1_is_stationary_23; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_24_2_data = io_in_c_bypass_regNext_24_2_data_23; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_24_2_is_stationary = io_in_c_bypass_regNext_24_2_is_stationary_23; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_24_3_data = io_in_c_bypass_regNext_24_3_data_23; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_24_3_is_stationary = io_in_c_bypass_regNext_24_3_is_stationary_23; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_25_0_data = io_in_c_bypass_regNext_25_0_data_24; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_25_0_is_stationary = io_in_c_bypass_regNext_25_0_is_stationary_24; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_25_1_data = io_in_c_bypass_regNext_25_1_data_24; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_25_1_is_stationary = io_in_c_bypass_regNext_25_1_is_stationary_24; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_25_2_data = io_in_c_bypass_regNext_25_2_data_24; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_25_2_is_stationary = io_in_c_bypass_regNext_25_2_is_stationary_24; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_25_3_data = io_in_c_bypass_regNext_25_3_data_24; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_25_3_is_stationary = io_in_c_bypass_regNext_25_3_is_stationary_24; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_26_0_data = io_in_c_bypass_regNext_26_0_data_25; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_26_0_is_stationary = io_in_c_bypass_regNext_26_0_is_stationary_25; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_26_1_data = io_in_c_bypass_regNext_26_1_data_25; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_26_1_is_stationary = io_in_c_bypass_regNext_26_1_is_stationary_25; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_26_2_data = io_in_c_bypass_regNext_26_2_data_25; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_26_2_is_stationary = io_in_c_bypass_regNext_26_2_is_stationary_25; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_26_3_data = io_in_c_bypass_regNext_26_3_data_25; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_26_3_is_stationary = io_in_c_bypass_regNext_26_3_is_stationary_25; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_27_0_data = io_in_c_bypass_regNext_27_0_data_26; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_27_0_is_stationary = io_in_c_bypass_regNext_27_0_is_stationary_26; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_27_1_data = io_in_c_bypass_regNext_27_1_data_26; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_27_1_is_stationary = io_in_c_bypass_regNext_27_1_is_stationary_26; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_27_2_data = io_in_c_bypass_regNext_27_2_data_26; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_27_2_is_stationary = io_in_c_bypass_regNext_27_2_is_stationary_26; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_27_3_data = io_in_c_bypass_regNext_27_3_data_26; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_27_3_is_stationary = io_in_c_bypass_regNext_27_3_is_stationary_26; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_28_0_data = io_in_c_bypass_regNext_28_0_data_27; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_28_0_is_stationary = io_in_c_bypass_regNext_28_0_is_stationary_27; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_28_1_data = io_in_c_bypass_regNext_28_1_data_27; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_28_1_is_stationary = io_in_c_bypass_regNext_28_1_is_stationary_27; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_28_2_data = io_in_c_bypass_regNext_28_2_data_27; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_28_2_is_stationary = io_in_c_bypass_regNext_28_2_is_stationary_27; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_28_3_data = io_in_c_bypass_regNext_28_3_data_27; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_28_3_is_stationary = io_in_c_bypass_regNext_28_3_is_stationary_27; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_29_0_data = io_in_c_bypass_regNext_29_0_data_28; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_29_0_is_stationary = io_in_c_bypass_regNext_29_0_is_stationary_28; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_29_1_data = io_in_c_bypass_regNext_29_1_data_28; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_29_1_is_stationary = io_in_c_bypass_regNext_29_1_is_stationary_28; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_29_2_data = io_in_c_bypass_regNext_29_2_data_28; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_29_2_is_stationary = io_in_c_bypass_regNext_29_2_is_stationary_28; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_29_3_data = io_in_c_bypass_regNext_29_3_data_28; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_29_3_is_stationary = io_in_c_bypass_regNext_29_3_is_stationary_28; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_30_0_data = io_in_c_bypass_regNext_30_0_data_29; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_30_0_is_stationary = io_in_c_bypass_regNext_30_0_is_stationary_29; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_30_1_data = io_in_c_bypass_regNext_30_1_data_29; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_30_1_is_stationary = io_in_c_bypass_regNext_30_1_is_stationary_29; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_30_2_data = io_in_c_bypass_regNext_30_2_data_29; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_30_2_is_stationary = io_in_c_bypass_regNext_30_2_is_stationary_29; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_30_3_data = io_in_c_bypass_regNext_30_3_data_29; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_30_3_is_stationary = io_in_c_bypass_regNext_30_3_is_stationary_29; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_31_0_data = io_in_c_bypass_regNext_31_0_data_30; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_31_0_is_stationary = io_in_c_bypass_regNext_31_0_is_stationary_30; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_31_1_data = io_in_c_bypass_regNext_31_1_data_30; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_31_1_is_stationary = io_in_c_bypass_regNext_31_1_is_stationary_30; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_31_2_data = io_in_c_bypass_regNext_31_2_data_30; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_31_2_is_stationary = io_in_c_bypass_regNext_31_2_is_stationary_30; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_31_3_data = io_in_c_bypass_regNext_31_3_data_30; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_31_3_is_stationary = io_in_c_bypass_regNext_31_3_is_stationary_30; // @[ArraySARA.scala 101:26]
  assign io_out_r_input_from_bypass_0 = io_in_r_input_from_bypass_regNext_0; // @[ArraySARA.scala 103:30]
  assign io_out_r_input_from_bypass_1 = io_in_r_input_from_bypass_regNext_1; // @[ArraySARA.scala 103:30]
  assign io_out_r_input_from_bypass_2 = io_in_r_input_from_bypass_regNext_2; // @[ArraySARA.scala 103:30]
  assign io_out_r_input_from_bypass_3 = io_in_r_input_from_bypass_regNext_3; // @[ArraySARA.scala 103:30]
  assign io_out_r_input_from_bypass_4 = io_in_r_input_from_bypass_regNext_4; // @[ArraySARA.scala 103:30]
  assign io_out_r_input_from_bypass_5 = io_in_r_input_from_bypass_regNext_5; // @[ArraySARA.scala 103:30]
  assign io_out_r_input_from_bypass_6 = io_in_r_input_from_bypass_regNext_6; // @[ArraySARA.scala 103:30]
  assign io_out_r_input_from_bypass_7 = io_in_r_input_from_bypass_regNext_7; // @[ArraySARA.scala 103:30]
  assign io_out_r_input_from_bypass_8 = io_in_r_input_from_bypass_regNext_8; // @[ArraySARA.scala 103:30]
  assign io_out_r_input_from_bypass_9 = io_in_r_input_from_bypass_regNext_9; // @[ArraySARA.scala 103:30]
  assign io_out_r_input_from_bypass_10 = io_in_r_input_from_bypass_regNext_10; // @[ArraySARA.scala 103:30]
  assign io_out_r_input_from_bypass_11 = io_in_r_input_from_bypass_regNext_11; // @[ArraySARA.scala 103:30]
  assign io_out_r_input_from_bypass_12 = io_in_r_input_from_bypass_regNext_12; // @[ArraySARA.scala 103:30]
  assign io_out_r_input_from_bypass_13 = io_in_r_input_from_bypass_regNext_13; // @[ArraySARA.scala 103:30]
  assign io_out_r_input_from_bypass_14 = io_in_r_input_from_bypass_regNext_14; // @[ArraySARA.scala 103:30]
  assign io_out_r_input_from_bypass_15 = io_in_r_input_from_bypass_regNext_15; // @[ArraySARA.scala 103:30]
  assign io_out_r_input_from_bypass_16 = io_in_r_input_from_bypass_regNext_16; // @[ArraySARA.scala 103:30]
  assign io_out_r_input_from_bypass_17 = io_in_r_input_from_bypass_regNext_17; // @[ArraySARA.scala 103:30]
  assign io_out_r_input_from_bypass_18 = io_in_r_input_from_bypass_regNext_18; // @[ArraySARA.scala 103:30]
  assign io_out_r_input_from_bypass_19 = io_in_r_input_from_bypass_regNext_19; // @[ArraySARA.scala 103:30]
  assign io_out_r_input_from_bypass_20 = io_in_r_input_from_bypass_regNext_20; // @[ArraySARA.scala 103:30]
  assign io_out_r_input_from_bypass_21 = io_in_r_input_from_bypass_regNext_21; // @[ArraySARA.scala 103:30]
  assign io_out_r_input_from_bypass_22 = io_in_r_input_from_bypass_regNext_22; // @[ArraySARA.scala 103:30]
  assign io_out_r_input_from_bypass_23 = io_in_r_input_from_bypass_regNext_23; // @[ArraySARA.scala 103:30]
  assign io_out_r_input_from_bypass_24 = io_in_r_input_from_bypass_regNext_24; // @[ArraySARA.scala 103:30]
  assign io_out_r_input_from_bypass_25 = io_in_r_input_from_bypass_regNext_25; // @[ArraySARA.scala 103:30]
  assign io_out_r_input_from_bypass_26 = io_in_r_input_from_bypass_regNext_26; // @[ArraySARA.scala 103:30]
  assign io_out_r_input_from_bypass_27 = io_in_r_input_from_bypass_regNext_27; // @[ArraySARA.scala 103:30]
  assign io_out_r_input_from_bypass_28 = io_in_r_input_from_bypass_regNext_28; // @[ArraySARA.scala 103:30]
  assign io_out_r_input_from_bypass_29 = io_in_r_input_from_bypass_regNext_29; // @[ArraySARA.scala 103:30]
  assign io_out_r_input_from_bypass_30 = io_in_r_input_from_bypass_regNext_30; // @[ArraySARA.scala 103:30]
  assign io_out_r_input_from_bypass_31 = io_in_r_input_from_bypass_regNext_31; // @[ArraySARA.scala 103:30]
  assign io_out_c_input_from_bypass_0 = io_in_c_input_from_bypass_regNext_0; // @[ArraySARA.scala 104:30]
  assign io_out_c_input_from_bypass_1 = io_in_c_input_from_bypass_regNext_1; // @[ArraySARA.scala 104:30]
  assign io_out_c_input_from_bypass_2 = io_in_c_input_from_bypass_regNext_2; // @[ArraySARA.scala 104:30]
  assign io_out_c_input_from_bypass_3 = io_in_c_input_from_bypass_regNext_3; // @[ArraySARA.scala 104:30]
  assign io_out_c_input_from_bypass_4 = io_in_c_input_from_bypass_regNext_4; // @[ArraySARA.scala 104:30]
  assign io_out_c_input_from_bypass_5 = io_in_c_input_from_bypass_regNext_5; // @[ArraySARA.scala 104:30]
  assign io_out_c_input_from_bypass_6 = io_in_c_input_from_bypass_regNext_6; // @[ArraySARA.scala 104:30]
  assign io_out_c_input_from_bypass_7 = io_in_c_input_from_bypass_regNext_7; // @[ArraySARA.scala 104:30]
  assign io_out_c_input_from_bypass_8 = io_in_c_input_from_bypass_regNext_8; // @[ArraySARA.scala 104:30]
  assign io_out_c_input_from_bypass_9 = io_in_c_input_from_bypass_regNext_9; // @[ArraySARA.scala 104:30]
  assign io_out_c_input_from_bypass_10 = io_in_c_input_from_bypass_regNext_10; // @[ArraySARA.scala 104:30]
  assign io_out_c_input_from_bypass_11 = io_in_c_input_from_bypass_regNext_11; // @[ArraySARA.scala 104:30]
  assign io_out_c_input_from_bypass_12 = io_in_c_input_from_bypass_regNext_12; // @[ArraySARA.scala 104:30]
  assign io_out_c_input_from_bypass_13 = io_in_c_input_from_bypass_regNext_13; // @[ArraySARA.scala 104:30]
  assign io_out_c_input_from_bypass_14 = io_in_c_input_from_bypass_regNext_14; // @[ArraySARA.scala 104:30]
  assign io_out_c_input_from_bypass_15 = io_in_c_input_from_bypass_regNext_15; // @[ArraySARA.scala 104:30]
  assign io_out_c_input_from_bypass_16 = io_in_c_input_from_bypass_regNext_16; // @[ArraySARA.scala 104:30]
  assign io_out_c_input_from_bypass_17 = io_in_c_input_from_bypass_regNext_17; // @[ArraySARA.scala 104:30]
  assign io_out_c_input_from_bypass_18 = io_in_c_input_from_bypass_regNext_18; // @[ArraySARA.scala 104:30]
  assign io_out_c_input_from_bypass_19 = io_in_c_input_from_bypass_regNext_19; // @[ArraySARA.scala 104:30]
  assign io_out_c_input_from_bypass_20 = io_in_c_input_from_bypass_regNext_20; // @[ArraySARA.scala 104:30]
  assign io_out_c_input_from_bypass_21 = io_in_c_input_from_bypass_regNext_21; // @[ArraySARA.scala 104:30]
  assign io_out_c_input_from_bypass_22 = io_in_c_input_from_bypass_regNext_22; // @[ArraySARA.scala 104:30]
  assign io_out_c_input_from_bypass_23 = io_in_c_input_from_bypass_regNext_23; // @[ArraySARA.scala 104:30]
  assign io_out_c_input_from_bypass_24 = io_in_c_input_from_bypass_regNext_24; // @[ArraySARA.scala 104:30]
  assign io_out_c_input_from_bypass_25 = io_in_c_input_from_bypass_regNext_25; // @[ArraySARA.scala 104:30]
  assign io_out_c_input_from_bypass_26 = io_in_c_input_from_bypass_regNext_26; // @[ArraySARA.scala 104:30]
  assign io_out_c_input_from_bypass_27 = io_in_c_input_from_bypass_regNext_27; // @[ArraySARA.scala 104:30]
  assign io_out_c_input_from_bypass_28 = io_in_c_input_from_bypass_regNext_28; // @[ArraySARA.scala 104:30]
  assign io_out_c_input_from_bypass_29 = io_in_c_input_from_bypass_regNext_29; // @[ArraySARA.scala 104:30]
  assign io_out_c_input_from_bypass_30 = io_in_c_input_from_bypass_regNext_30; // @[ArraySARA.scala 104:30]
  assign io_out_c_input_from_bypass_31 = io_in_c_input_from_bypass_regNext_31; // @[ArraySARA.scala 104:30]
  always @(posedge clk) begin
    out_r_regNext_0_data <= out_r_0_data; // @[Reg.scala 39:30]
    out_r_regNext_0_load_store <= out_r_0_load_store; // @[Reg.scala 39:30]
    out_r_regNext_0_df_is_ws <= out_r_0_df_is_ws; // @[Reg.scala 39:30]
    out_r_regNext_0_stall <= out_r_0_stall; // @[Reg.scala 39:30]
    out_r_regNext_1_data <= out_r_1_data; // @[Reg.scala 39:30]
    out_r_regNext_1_load_store <= out_r_1_load_store; // @[Reg.scala 39:30]
    out_r_regNext_1_df_is_ws <= out_r_1_df_is_ws; // @[Reg.scala 39:30]
    out_r_regNext_1_stall <= out_r_1_stall; // @[Reg.scala 39:30]
    out_r_regNext_2_data <= out_r_2_data; // @[Reg.scala 39:30]
    out_r_regNext_2_load_store <= out_r_2_load_store; // @[Reg.scala 39:30]
    out_r_regNext_2_df_is_ws <= out_r_2_df_is_ws; // @[Reg.scala 39:30]
    out_r_regNext_2_stall <= out_r_2_stall; // @[Reg.scala 39:30]
    out_r_regNext_3_data <= out_r_3_data; // @[Reg.scala 39:30]
    out_r_regNext_3_load_store <= out_r_3_load_store; // @[Reg.scala 39:30]
    out_r_regNext_3_df_is_ws <= out_r_3_df_is_ws; // @[Reg.scala 39:30]
    out_r_regNext_3_stall <= out_r_3_stall; // @[Reg.scala 39:30]
    out_c_regNext_0_data <= out_c_0_data; // @[Reg.scala 39:30]
    out_c_regNext_0_is_stationary <= out_c_0_is_stationary; // @[Reg.scala 39:30]
    out_c_regNext_1_data <= out_c_1_data; // @[Reg.scala 39:30]
    out_c_regNext_1_is_stationary <= out_c_1_is_stationary; // @[Reg.scala 39:30]
    out_c_regNext_2_data <= out_c_2_data; // @[Reg.scala 39:30]
    out_c_regNext_2_is_stationary <= out_c_2_is_stationary; // @[Reg.scala 39:30]
    out_c_regNext_3_data <= out_c_3_data; // @[Reg.scala 39:30]
    out_c_regNext_3_is_stationary <= out_c_3_is_stationary; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_0_data <= io_in_r_bypass_0_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_0_load_store <= io_in_r_bypass_0_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_0_df_is_ws <= io_in_r_bypass_0_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_0_stall <= io_in_r_bypass_0_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_1_data <= io_in_r_bypass_0_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_1_load_store <= io_in_r_bypass_0_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_1_df_is_ws <= io_in_r_bypass_0_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_1_stall <= io_in_r_bypass_0_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_2_data <= io_in_r_bypass_0_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_2_load_store <= io_in_r_bypass_0_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_2_df_is_ws <= io_in_r_bypass_0_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_2_stall <= io_in_r_bypass_0_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_3_data <= io_in_r_bypass_0_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_3_load_store <= io_in_r_bypass_0_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_3_df_is_ws <= io_in_r_bypass_0_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_3_stall <= io_in_r_bypass_0_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_0_data <= io_in_r_bypass_1_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_0_load_store <= io_in_r_bypass_1_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_0_df_is_ws <= io_in_r_bypass_1_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_0_stall <= io_in_r_bypass_1_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_1_data <= io_in_r_bypass_1_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_1_load_store <= io_in_r_bypass_1_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_1_df_is_ws <= io_in_r_bypass_1_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_1_stall <= io_in_r_bypass_1_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_2_data <= io_in_r_bypass_1_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_2_load_store <= io_in_r_bypass_1_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_2_df_is_ws <= io_in_r_bypass_1_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_2_stall <= io_in_r_bypass_1_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_3_data <= io_in_r_bypass_1_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_3_load_store <= io_in_r_bypass_1_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_3_df_is_ws <= io_in_r_bypass_1_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_3_stall <= io_in_r_bypass_1_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_0_data <= io_in_r_bypass_2_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_0_load_store <= io_in_r_bypass_2_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_0_df_is_ws <= io_in_r_bypass_2_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_0_stall <= io_in_r_bypass_2_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_1_data <= io_in_r_bypass_2_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_1_load_store <= io_in_r_bypass_2_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_1_df_is_ws <= io_in_r_bypass_2_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_1_stall <= io_in_r_bypass_2_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_2_data <= io_in_r_bypass_2_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_2_load_store <= io_in_r_bypass_2_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_2_df_is_ws <= io_in_r_bypass_2_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_2_stall <= io_in_r_bypass_2_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_3_data <= io_in_r_bypass_2_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_3_load_store <= io_in_r_bypass_2_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_3_df_is_ws <= io_in_r_bypass_2_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_3_stall <= io_in_r_bypass_2_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_0_data <= io_in_r_bypass_3_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_0_load_store <= io_in_r_bypass_3_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_0_df_is_ws <= io_in_r_bypass_3_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_0_stall <= io_in_r_bypass_3_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_1_data <= io_in_r_bypass_3_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_1_load_store <= io_in_r_bypass_3_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_1_df_is_ws <= io_in_r_bypass_3_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_1_stall <= io_in_r_bypass_3_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_2_data <= io_in_r_bypass_3_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_2_load_store <= io_in_r_bypass_3_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_2_df_is_ws <= io_in_r_bypass_3_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_2_stall <= io_in_r_bypass_3_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_3_data <= io_in_r_bypass_3_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_3_load_store <= io_in_r_bypass_3_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_3_df_is_ws <= io_in_r_bypass_3_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_3_stall <= io_in_r_bypass_3_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_0_data <= io_in_r_bypass_4_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_0_load_store <= io_in_r_bypass_4_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_0_df_is_ws <= io_in_r_bypass_4_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_0_stall <= io_in_r_bypass_4_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_1_data <= io_in_r_bypass_4_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_1_load_store <= io_in_r_bypass_4_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_1_df_is_ws <= io_in_r_bypass_4_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_1_stall <= io_in_r_bypass_4_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_2_data <= io_in_r_bypass_4_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_2_load_store <= io_in_r_bypass_4_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_2_df_is_ws <= io_in_r_bypass_4_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_2_stall <= io_in_r_bypass_4_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_3_data <= io_in_r_bypass_4_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_3_load_store <= io_in_r_bypass_4_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_3_df_is_ws <= io_in_r_bypass_4_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_3_stall <= io_in_r_bypass_4_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_0_data <= io_in_r_bypass_5_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_0_load_store <= io_in_r_bypass_5_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_0_df_is_ws <= io_in_r_bypass_5_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_0_stall <= io_in_r_bypass_5_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_1_data <= io_in_r_bypass_5_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_1_load_store <= io_in_r_bypass_5_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_1_df_is_ws <= io_in_r_bypass_5_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_1_stall <= io_in_r_bypass_5_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_2_data <= io_in_r_bypass_5_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_2_load_store <= io_in_r_bypass_5_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_2_df_is_ws <= io_in_r_bypass_5_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_2_stall <= io_in_r_bypass_5_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_3_data <= io_in_r_bypass_5_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_3_load_store <= io_in_r_bypass_5_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_3_df_is_ws <= io_in_r_bypass_5_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_3_stall <= io_in_r_bypass_5_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_0_data <= io_in_r_bypass_6_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_0_load_store <= io_in_r_bypass_6_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_0_df_is_ws <= io_in_r_bypass_6_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_0_stall <= io_in_r_bypass_6_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_1_data <= io_in_r_bypass_6_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_1_load_store <= io_in_r_bypass_6_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_1_df_is_ws <= io_in_r_bypass_6_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_1_stall <= io_in_r_bypass_6_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_2_data <= io_in_r_bypass_6_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_2_load_store <= io_in_r_bypass_6_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_2_df_is_ws <= io_in_r_bypass_6_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_2_stall <= io_in_r_bypass_6_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_3_data <= io_in_r_bypass_6_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_3_load_store <= io_in_r_bypass_6_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_3_df_is_ws <= io_in_r_bypass_6_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_3_stall <= io_in_r_bypass_6_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_0_data <= io_in_r_bypass_7_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_0_load_store <= io_in_r_bypass_7_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_0_df_is_ws <= io_in_r_bypass_7_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_0_stall <= io_in_r_bypass_7_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_1_data <= io_in_r_bypass_7_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_1_load_store <= io_in_r_bypass_7_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_1_df_is_ws <= io_in_r_bypass_7_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_1_stall <= io_in_r_bypass_7_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_2_data <= io_in_r_bypass_7_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_2_load_store <= io_in_r_bypass_7_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_2_df_is_ws <= io_in_r_bypass_7_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_2_stall <= io_in_r_bypass_7_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_3_data <= io_in_r_bypass_7_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_3_load_store <= io_in_r_bypass_7_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_3_df_is_ws <= io_in_r_bypass_7_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_3_stall <= io_in_r_bypass_7_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_0_data <= io_in_r_bypass_8_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_0_load_store <= io_in_r_bypass_8_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_0_df_is_ws <= io_in_r_bypass_8_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_0_stall <= io_in_r_bypass_8_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_1_data <= io_in_r_bypass_8_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_1_load_store <= io_in_r_bypass_8_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_1_df_is_ws <= io_in_r_bypass_8_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_1_stall <= io_in_r_bypass_8_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_2_data <= io_in_r_bypass_8_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_2_load_store <= io_in_r_bypass_8_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_2_df_is_ws <= io_in_r_bypass_8_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_2_stall <= io_in_r_bypass_8_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_3_data <= io_in_r_bypass_8_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_3_load_store <= io_in_r_bypass_8_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_3_df_is_ws <= io_in_r_bypass_8_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_3_stall <= io_in_r_bypass_8_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_0_data <= io_in_r_bypass_9_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_0_load_store <= io_in_r_bypass_9_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_0_df_is_ws <= io_in_r_bypass_9_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_0_stall <= io_in_r_bypass_9_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_1_data <= io_in_r_bypass_9_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_1_load_store <= io_in_r_bypass_9_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_1_df_is_ws <= io_in_r_bypass_9_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_1_stall <= io_in_r_bypass_9_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_2_data <= io_in_r_bypass_9_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_2_load_store <= io_in_r_bypass_9_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_2_df_is_ws <= io_in_r_bypass_9_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_2_stall <= io_in_r_bypass_9_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_3_data <= io_in_r_bypass_9_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_3_load_store <= io_in_r_bypass_9_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_3_df_is_ws <= io_in_r_bypass_9_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_3_stall <= io_in_r_bypass_9_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_0_data <= io_in_r_bypass_10_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_0_load_store <= io_in_r_bypass_10_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_0_df_is_ws <= io_in_r_bypass_10_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_0_stall <= io_in_r_bypass_10_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_1_data <= io_in_r_bypass_10_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_1_load_store <= io_in_r_bypass_10_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_1_df_is_ws <= io_in_r_bypass_10_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_1_stall <= io_in_r_bypass_10_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_2_data <= io_in_r_bypass_10_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_2_load_store <= io_in_r_bypass_10_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_2_df_is_ws <= io_in_r_bypass_10_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_2_stall <= io_in_r_bypass_10_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_3_data <= io_in_r_bypass_10_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_3_load_store <= io_in_r_bypass_10_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_3_df_is_ws <= io_in_r_bypass_10_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_3_stall <= io_in_r_bypass_10_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_0_data <= io_in_r_bypass_11_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_0_load_store <= io_in_r_bypass_11_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_0_df_is_ws <= io_in_r_bypass_11_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_0_stall <= io_in_r_bypass_11_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_1_data <= io_in_r_bypass_11_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_1_load_store <= io_in_r_bypass_11_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_1_df_is_ws <= io_in_r_bypass_11_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_1_stall <= io_in_r_bypass_11_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_2_data <= io_in_r_bypass_11_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_2_load_store <= io_in_r_bypass_11_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_2_df_is_ws <= io_in_r_bypass_11_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_2_stall <= io_in_r_bypass_11_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_3_data <= io_in_r_bypass_11_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_3_load_store <= io_in_r_bypass_11_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_3_df_is_ws <= io_in_r_bypass_11_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_3_stall <= io_in_r_bypass_11_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_0_data <= io_in_r_bypass_12_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_0_load_store <= io_in_r_bypass_12_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_0_df_is_ws <= io_in_r_bypass_12_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_0_stall <= io_in_r_bypass_12_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_1_data <= io_in_r_bypass_12_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_1_load_store <= io_in_r_bypass_12_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_1_df_is_ws <= io_in_r_bypass_12_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_1_stall <= io_in_r_bypass_12_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_2_data <= io_in_r_bypass_12_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_2_load_store <= io_in_r_bypass_12_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_2_df_is_ws <= io_in_r_bypass_12_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_2_stall <= io_in_r_bypass_12_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_3_data <= io_in_r_bypass_12_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_3_load_store <= io_in_r_bypass_12_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_3_df_is_ws <= io_in_r_bypass_12_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_3_stall <= io_in_r_bypass_12_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_0_data <= io_in_r_bypass_13_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_0_load_store <= io_in_r_bypass_13_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_0_df_is_ws <= io_in_r_bypass_13_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_0_stall <= io_in_r_bypass_13_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_1_data <= io_in_r_bypass_13_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_1_load_store <= io_in_r_bypass_13_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_1_df_is_ws <= io_in_r_bypass_13_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_1_stall <= io_in_r_bypass_13_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_2_data <= io_in_r_bypass_13_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_2_load_store <= io_in_r_bypass_13_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_2_df_is_ws <= io_in_r_bypass_13_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_2_stall <= io_in_r_bypass_13_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_3_data <= io_in_r_bypass_13_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_3_load_store <= io_in_r_bypass_13_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_3_df_is_ws <= io_in_r_bypass_13_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_3_stall <= io_in_r_bypass_13_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_0_data <= io_in_r_bypass_14_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_0_load_store <= io_in_r_bypass_14_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_0_df_is_ws <= io_in_r_bypass_14_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_0_stall <= io_in_r_bypass_14_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_1_data <= io_in_r_bypass_14_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_1_load_store <= io_in_r_bypass_14_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_1_df_is_ws <= io_in_r_bypass_14_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_1_stall <= io_in_r_bypass_14_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_2_data <= io_in_r_bypass_14_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_2_load_store <= io_in_r_bypass_14_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_2_df_is_ws <= io_in_r_bypass_14_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_2_stall <= io_in_r_bypass_14_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_3_data <= io_in_r_bypass_14_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_3_load_store <= io_in_r_bypass_14_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_3_df_is_ws <= io_in_r_bypass_14_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_3_stall <= io_in_r_bypass_14_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_0_data <= io_in_r_bypass_15_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_0_load_store <= io_in_r_bypass_15_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_0_df_is_ws <= io_in_r_bypass_15_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_0_stall <= io_in_r_bypass_15_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_1_data <= io_in_r_bypass_15_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_1_load_store <= io_in_r_bypass_15_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_1_df_is_ws <= io_in_r_bypass_15_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_1_stall <= io_in_r_bypass_15_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_2_data <= io_in_r_bypass_15_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_2_load_store <= io_in_r_bypass_15_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_2_df_is_ws <= io_in_r_bypass_15_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_2_stall <= io_in_r_bypass_15_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_3_data <= io_in_r_bypass_15_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_3_load_store <= io_in_r_bypass_15_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_3_df_is_ws <= io_in_r_bypass_15_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_3_stall <= io_in_r_bypass_15_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_0_data <= io_in_r_bypass_16_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_0_load_store <= io_in_r_bypass_16_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_0_df_is_ws <= io_in_r_bypass_16_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_0_stall <= io_in_r_bypass_16_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_1_data <= io_in_r_bypass_16_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_1_load_store <= io_in_r_bypass_16_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_1_df_is_ws <= io_in_r_bypass_16_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_1_stall <= io_in_r_bypass_16_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_2_data <= io_in_r_bypass_16_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_2_load_store <= io_in_r_bypass_16_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_2_df_is_ws <= io_in_r_bypass_16_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_2_stall <= io_in_r_bypass_16_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_3_data <= io_in_r_bypass_16_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_3_load_store <= io_in_r_bypass_16_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_3_df_is_ws <= io_in_r_bypass_16_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_3_stall <= io_in_r_bypass_16_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_0_data <= io_in_r_bypass_17_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_0_load_store <= io_in_r_bypass_17_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_0_df_is_ws <= io_in_r_bypass_17_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_0_stall <= io_in_r_bypass_17_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_1_data <= io_in_r_bypass_17_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_1_load_store <= io_in_r_bypass_17_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_1_df_is_ws <= io_in_r_bypass_17_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_1_stall <= io_in_r_bypass_17_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_2_data <= io_in_r_bypass_17_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_2_load_store <= io_in_r_bypass_17_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_2_df_is_ws <= io_in_r_bypass_17_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_2_stall <= io_in_r_bypass_17_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_3_data <= io_in_r_bypass_17_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_3_load_store <= io_in_r_bypass_17_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_3_df_is_ws <= io_in_r_bypass_17_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_3_stall <= io_in_r_bypass_17_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_0_data <= io_in_r_bypass_18_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_0_load_store <= io_in_r_bypass_18_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_0_df_is_ws <= io_in_r_bypass_18_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_0_stall <= io_in_r_bypass_18_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_1_data <= io_in_r_bypass_18_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_1_load_store <= io_in_r_bypass_18_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_1_df_is_ws <= io_in_r_bypass_18_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_1_stall <= io_in_r_bypass_18_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_2_data <= io_in_r_bypass_18_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_2_load_store <= io_in_r_bypass_18_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_2_df_is_ws <= io_in_r_bypass_18_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_2_stall <= io_in_r_bypass_18_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_3_data <= io_in_r_bypass_18_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_3_load_store <= io_in_r_bypass_18_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_3_df_is_ws <= io_in_r_bypass_18_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_3_stall <= io_in_r_bypass_18_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_0_data <= io_in_r_bypass_19_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_0_load_store <= io_in_r_bypass_19_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_0_df_is_ws <= io_in_r_bypass_19_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_0_stall <= io_in_r_bypass_19_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_1_data <= io_in_r_bypass_19_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_1_load_store <= io_in_r_bypass_19_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_1_df_is_ws <= io_in_r_bypass_19_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_1_stall <= io_in_r_bypass_19_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_2_data <= io_in_r_bypass_19_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_2_load_store <= io_in_r_bypass_19_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_2_df_is_ws <= io_in_r_bypass_19_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_2_stall <= io_in_r_bypass_19_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_3_data <= io_in_r_bypass_19_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_3_load_store <= io_in_r_bypass_19_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_3_df_is_ws <= io_in_r_bypass_19_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_3_stall <= io_in_r_bypass_19_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_0_data <= io_in_r_bypass_20_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_0_load_store <= io_in_r_bypass_20_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_0_df_is_ws <= io_in_r_bypass_20_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_0_stall <= io_in_r_bypass_20_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_1_data <= io_in_r_bypass_20_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_1_load_store <= io_in_r_bypass_20_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_1_df_is_ws <= io_in_r_bypass_20_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_1_stall <= io_in_r_bypass_20_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_2_data <= io_in_r_bypass_20_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_2_load_store <= io_in_r_bypass_20_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_2_df_is_ws <= io_in_r_bypass_20_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_2_stall <= io_in_r_bypass_20_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_3_data <= io_in_r_bypass_20_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_3_load_store <= io_in_r_bypass_20_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_3_df_is_ws <= io_in_r_bypass_20_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_3_stall <= io_in_r_bypass_20_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_0_data <= io_in_r_bypass_21_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_0_load_store <= io_in_r_bypass_21_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_0_df_is_ws <= io_in_r_bypass_21_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_0_stall <= io_in_r_bypass_21_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_1_data <= io_in_r_bypass_21_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_1_load_store <= io_in_r_bypass_21_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_1_df_is_ws <= io_in_r_bypass_21_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_1_stall <= io_in_r_bypass_21_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_2_data <= io_in_r_bypass_21_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_2_load_store <= io_in_r_bypass_21_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_2_df_is_ws <= io_in_r_bypass_21_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_2_stall <= io_in_r_bypass_21_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_3_data <= io_in_r_bypass_21_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_3_load_store <= io_in_r_bypass_21_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_3_df_is_ws <= io_in_r_bypass_21_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_3_stall <= io_in_r_bypass_21_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_0_data <= io_in_r_bypass_22_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_0_load_store <= io_in_r_bypass_22_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_0_df_is_ws <= io_in_r_bypass_22_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_0_stall <= io_in_r_bypass_22_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_1_data <= io_in_r_bypass_22_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_1_load_store <= io_in_r_bypass_22_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_1_df_is_ws <= io_in_r_bypass_22_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_1_stall <= io_in_r_bypass_22_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_2_data <= io_in_r_bypass_22_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_2_load_store <= io_in_r_bypass_22_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_2_df_is_ws <= io_in_r_bypass_22_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_2_stall <= io_in_r_bypass_22_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_3_data <= io_in_r_bypass_22_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_3_load_store <= io_in_r_bypass_22_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_3_df_is_ws <= io_in_r_bypass_22_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_3_stall <= io_in_r_bypass_22_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_0_data <= io_in_r_bypass_23_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_0_load_store <= io_in_r_bypass_23_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_0_df_is_ws <= io_in_r_bypass_23_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_0_stall <= io_in_r_bypass_23_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_1_data <= io_in_r_bypass_23_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_1_load_store <= io_in_r_bypass_23_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_1_df_is_ws <= io_in_r_bypass_23_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_1_stall <= io_in_r_bypass_23_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_2_data <= io_in_r_bypass_23_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_2_load_store <= io_in_r_bypass_23_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_2_df_is_ws <= io_in_r_bypass_23_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_2_stall <= io_in_r_bypass_23_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_3_data <= io_in_r_bypass_23_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_3_load_store <= io_in_r_bypass_23_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_3_df_is_ws <= io_in_r_bypass_23_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_3_stall <= io_in_r_bypass_23_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_0_data <= io_in_r_bypass_24_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_0_load_store <= io_in_r_bypass_24_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_0_df_is_ws <= io_in_r_bypass_24_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_0_stall <= io_in_r_bypass_24_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_1_data <= io_in_r_bypass_24_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_1_load_store <= io_in_r_bypass_24_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_1_df_is_ws <= io_in_r_bypass_24_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_1_stall <= io_in_r_bypass_24_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_2_data <= io_in_r_bypass_24_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_2_load_store <= io_in_r_bypass_24_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_2_df_is_ws <= io_in_r_bypass_24_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_2_stall <= io_in_r_bypass_24_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_3_data <= io_in_r_bypass_24_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_3_load_store <= io_in_r_bypass_24_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_3_df_is_ws <= io_in_r_bypass_24_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_3_stall <= io_in_r_bypass_24_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_0_data <= io_in_r_bypass_25_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_0_load_store <= io_in_r_bypass_25_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_0_df_is_ws <= io_in_r_bypass_25_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_0_stall <= io_in_r_bypass_25_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_1_data <= io_in_r_bypass_25_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_1_load_store <= io_in_r_bypass_25_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_1_df_is_ws <= io_in_r_bypass_25_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_1_stall <= io_in_r_bypass_25_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_2_data <= io_in_r_bypass_25_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_2_load_store <= io_in_r_bypass_25_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_2_df_is_ws <= io_in_r_bypass_25_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_2_stall <= io_in_r_bypass_25_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_3_data <= io_in_r_bypass_25_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_3_load_store <= io_in_r_bypass_25_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_3_df_is_ws <= io_in_r_bypass_25_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_3_stall <= io_in_r_bypass_25_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_0_data <= io_in_r_bypass_26_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_0_load_store <= io_in_r_bypass_26_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_0_df_is_ws <= io_in_r_bypass_26_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_0_stall <= io_in_r_bypass_26_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_1_data <= io_in_r_bypass_26_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_1_load_store <= io_in_r_bypass_26_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_1_df_is_ws <= io_in_r_bypass_26_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_1_stall <= io_in_r_bypass_26_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_2_data <= io_in_r_bypass_26_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_2_load_store <= io_in_r_bypass_26_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_2_df_is_ws <= io_in_r_bypass_26_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_2_stall <= io_in_r_bypass_26_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_3_data <= io_in_r_bypass_26_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_3_load_store <= io_in_r_bypass_26_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_3_df_is_ws <= io_in_r_bypass_26_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_3_stall <= io_in_r_bypass_26_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_0_data <= io_in_r_bypass_27_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_0_load_store <= io_in_r_bypass_27_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_0_df_is_ws <= io_in_r_bypass_27_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_0_stall <= io_in_r_bypass_27_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_1_data <= io_in_r_bypass_27_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_1_load_store <= io_in_r_bypass_27_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_1_df_is_ws <= io_in_r_bypass_27_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_1_stall <= io_in_r_bypass_27_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_2_data <= io_in_r_bypass_27_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_2_load_store <= io_in_r_bypass_27_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_2_df_is_ws <= io_in_r_bypass_27_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_2_stall <= io_in_r_bypass_27_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_3_data <= io_in_r_bypass_27_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_3_load_store <= io_in_r_bypass_27_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_3_df_is_ws <= io_in_r_bypass_27_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_3_stall <= io_in_r_bypass_27_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_0_data <= io_in_r_bypass_28_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_0_load_store <= io_in_r_bypass_28_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_0_df_is_ws <= io_in_r_bypass_28_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_0_stall <= io_in_r_bypass_28_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_1_data <= io_in_r_bypass_28_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_1_load_store <= io_in_r_bypass_28_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_1_df_is_ws <= io_in_r_bypass_28_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_1_stall <= io_in_r_bypass_28_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_2_data <= io_in_r_bypass_28_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_2_load_store <= io_in_r_bypass_28_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_2_df_is_ws <= io_in_r_bypass_28_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_2_stall <= io_in_r_bypass_28_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_3_data <= io_in_r_bypass_28_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_3_load_store <= io_in_r_bypass_28_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_3_df_is_ws <= io_in_r_bypass_28_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_3_stall <= io_in_r_bypass_28_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_0_data <= io_in_r_bypass_29_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_0_load_store <= io_in_r_bypass_29_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_0_df_is_ws <= io_in_r_bypass_29_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_0_stall <= io_in_r_bypass_29_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_1_data <= io_in_r_bypass_29_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_1_load_store <= io_in_r_bypass_29_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_1_df_is_ws <= io_in_r_bypass_29_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_1_stall <= io_in_r_bypass_29_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_2_data <= io_in_r_bypass_29_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_2_load_store <= io_in_r_bypass_29_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_2_df_is_ws <= io_in_r_bypass_29_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_2_stall <= io_in_r_bypass_29_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_3_data <= io_in_r_bypass_29_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_3_load_store <= io_in_r_bypass_29_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_3_df_is_ws <= io_in_r_bypass_29_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_3_stall <= io_in_r_bypass_29_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_0_data <= io_in_r_bypass_30_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_0_load_store <= io_in_r_bypass_30_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_0_df_is_ws <= io_in_r_bypass_30_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_0_stall <= io_in_r_bypass_30_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_1_data <= io_in_r_bypass_30_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_1_load_store <= io_in_r_bypass_30_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_1_df_is_ws <= io_in_r_bypass_30_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_1_stall <= io_in_r_bypass_30_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_2_data <= io_in_r_bypass_30_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_2_load_store <= io_in_r_bypass_30_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_2_df_is_ws <= io_in_r_bypass_30_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_2_stall <= io_in_r_bypass_30_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_3_data <= io_in_r_bypass_30_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_3_load_store <= io_in_r_bypass_30_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_3_df_is_ws <= io_in_r_bypass_30_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_3_stall <= io_in_r_bypass_30_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_0_data <= io_in_r_bypass_31_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_0_load_store <= io_in_r_bypass_31_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_0_df_is_ws <= io_in_r_bypass_31_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_0_stall <= io_in_r_bypass_31_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_1_data <= io_in_r_bypass_31_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_1_load_store <= io_in_r_bypass_31_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_1_df_is_ws <= io_in_r_bypass_31_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_1_stall <= io_in_r_bypass_31_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_2_data <= io_in_r_bypass_31_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_2_load_store <= io_in_r_bypass_31_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_2_df_is_ws <= io_in_r_bypass_31_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_2_stall <= io_in_r_bypass_31_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_3_data <= io_in_r_bypass_31_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_3_load_store <= io_in_r_bypass_31_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_3_df_is_ws <= io_in_r_bypass_31_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_3_stall <= io_in_r_bypass_31_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_0_data_1 <= io_in_r_bypass_0_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_0_load_store_1 <= io_in_r_bypass_0_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_0_df_is_ws_1 <= io_in_r_bypass_0_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_0_stall_1 <= io_in_r_bypass_0_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_1_data_1 <= io_in_r_bypass_0_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_1_load_store_1 <= io_in_r_bypass_0_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_1_df_is_ws_1 <= io_in_r_bypass_0_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_1_stall_1 <= io_in_r_bypass_0_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_2_data_1 <= io_in_r_bypass_0_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_2_load_store_1 <= io_in_r_bypass_0_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_2_df_is_ws_1 <= io_in_r_bypass_0_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_2_stall_1 <= io_in_r_bypass_0_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_3_data_1 <= io_in_r_bypass_0_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_3_load_store_1 <= io_in_r_bypass_0_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_3_df_is_ws_1 <= io_in_r_bypass_0_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_3_stall_1 <= io_in_r_bypass_0_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_0_data_1 <= io_in_r_bypass_1_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_0_load_store_1 <= io_in_r_bypass_1_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_0_df_is_ws_1 <= io_in_r_bypass_1_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_0_stall_1 <= io_in_r_bypass_1_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_1_data_1 <= io_in_r_bypass_1_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_1_load_store_1 <= io_in_r_bypass_1_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_1_df_is_ws_1 <= io_in_r_bypass_1_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_1_stall_1 <= io_in_r_bypass_1_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_2_data_1 <= io_in_r_bypass_1_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_2_load_store_1 <= io_in_r_bypass_1_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_2_df_is_ws_1 <= io_in_r_bypass_1_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_2_stall_1 <= io_in_r_bypass_1_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_3_data_1 <= io_in_r_bypass_1_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_3_load_store_1 <= io_in_r_bypass_1_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_3_df_is_ws_1 <= io_in_r_bypass_1_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_3_stall_1 <= io_in_r_bypass_1_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_0_data_1 <= io_in_r_bypass_2_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_0_load_store_1 <= io_in_r_bypass_2_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_0_df_is_ws_1 <= io_in_r_bypass_2_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_0_stall_1 <= io_in_r_bypass_2_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_1_data_1 <= io_in_r_bypass_2_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_1_load_store_1 <= io_in_r_bypass_2_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_1_df_is_ws_1 <= io_in_r_bypass_2_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_1_stall_1 <= io_in_r_bypass_2_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_2_data_1 <= io_in_r_bypass_2_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_2_load_store_1 <= io_in_r_bypass_2_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_2_df_is_ws_1 <= io_in_r_bypass_2_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_2_stall_1 <= io_in_r_bypass_2_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_3_data_1 <= io_in_r_bypass_2_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_3_load_store_1 <= io_in_r_bypass_2_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_3_df_is_ws_1 <= io_in_r_bypass_2_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_3_stall_1 <= io_in_r_bypass_2_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_0_data_1 <= io_in_r_bypass_3_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_0_load_store_1 <= io_in_r_bypass_3_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_0_df_is_ws_1 <= io_in_r_bypass_3_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_0_stall_1 <= io_in_r_bypass_3_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_1_data_1 <= io_in_r_bypass_3_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_1_load_store_1 <= io_in_r_bypass_3_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_1_df_is_ws_1 <= io_in_r_bypass_3_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_1_stall_1 <= io_in_r_bypass_3_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_2_data_1 <= io_in_r_bypass_3_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_2_load_store_1 <= io_in_r_bypass_3_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_2_df_is_ws_1 <= io_in_r_bypass_3_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_2_stall_1 <= io_in_r_bypass_3_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_3_data_1 <= io_in_r_bypass_3_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_3_load_store_1 <= io_in_r_bypass_3_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_3_df_is_ws_1 <= io_in_r_bypass_3_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_3_stall_1 <= io_in_r_bypass_3_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_0_data_1 <= io_in_r_bypass_4_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_0_load_store_1 <= io_in_r_bypass_4_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_0_df_is_ws_1 <= io_in_r_bypass_4_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_0_stall_1 <= io_in_r_bypass_4_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_1_data_1 <= io_in_r_bypass_4_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_1_load_store_1 <= io_in_r_bypass_4_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_1_df_is_ws_1 <= io_in_r_bypass_4_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_1_stall_1 <= io_in_r_bypass_4_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_2_data_1 <= io_in_r_bypass_4_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_2_load_store_1 <= io_in_r_bypass_4_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_2_df_is_ws_1 <= io_in_r_bypass_4_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_2_stall_1 <= io_in_r_bypass_4_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_3_data_1 <= io_in_r_bypass_4_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_3_load_store_1 <= io_in_r_bypass_4_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_3_df_is_ws_1 <= io_in_r_bypass_4_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_3_stall_1 <= io_in_r_bypass_4_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_0_data_1 <= io_in_r_bypass_5_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_0_load_store_1 <= io_in_r_bypass_5_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_0_df_is_ws_1 <= io_in_r_bypass_5_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_0_stall_1 <= io_in_r_bypass_5_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_1_data_1 <= io_in_r_bypass_5_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_1_load_store_1 <= io_in_r_bypass_5_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_1_df_is_ws_1 <= io_in_r_bypass_5_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_1_stall_1 <= io_in_r_bypass_5_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_2_data_1 <= io_in_r_bypass_5_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_2_load_store_1 <= io_in_r_bypass_5_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_2_df_is_ws_1 <= io_in_r_bypass_5_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_2_stall_1 <= io_in_r_bypass_5_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_3_data_1 <= io_in_r_bypass_5_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_3_load_store_1 <= io_in_r_bypass_5_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_3_df_is_ws_1 <= io_in_r_bypass_5_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_3_stall_1 <= io_in_r_bypass_5_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_0_data_1 <= io_in_r_bypass_6_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_0_load_store_1 <= io_in_r_bypass_6_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_0_df_is_ws_1 <= io_in_r_bypass_6_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_0_stall_1 <= io_in_r_bypass_6_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_1_data_1 <= io_in_r_bypass_6_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_1_load_store_1 <= io_in_r_bypass_6_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_1_df_is_ws_1 <= io_in_r_bypass_6_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_1_stall_1 <= io_in_r_bypass_6_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_2_data_1 <= io_in_r_bypass_6_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_2_load_store_1 <= io_in_r_bypass_6_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_2_df_is_ws_1 <= io_in_r_bypass_6_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_2_stall_1 <= io_in_r_bypass_6_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_3_data_1 <= io_in_r_bypass_6_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_3_load_store_1 <= io_in_r_bypass_6_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_3_df_is_ws_1 <= io_in_r_bypass_6_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_3_stall_1 <= io_in_r_bypass_6_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_0_data_1 <= io_in_r_bypass_7_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_0_load_store_1 <= io_in_r_bypass_7_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_0_df_is_ws_1 <= io_in_r_bypass_7_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_0_stall_1 <= io_in_r_bypass_7_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_1_data_1 <= io_in_r_bypass_7_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_1_load_store_1 <= io_in_r_bypass_7_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_1_df_is_ws_1 <= io_in_r_bypass_7_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_1_stall_1 <= io_in_r_bypass_7_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_2_data_1 <= io_in_r_bypass_7_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_2_load_store_1 <= io_in_r_bypass_7_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_2_df_is_ws_1 <= io_in_r_bypass_7_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_2_stall_1 <= io_in_r_bypass_7_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_3_data_1 <= io_in_r_bypass_7_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_3_load_store_1 <= io_in_r_bypass_7_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_3_df_is_ws_1 <= io_in_r_bypass_7_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_3_stall_1 <= io_in_r_bypass_7_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_0_data_1 <= io_in_r_bypass_8_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_0_load_store_1 <= io_in_r_bypass_8_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_0_df_is_ws_1 <= io_in_r_bypass_8_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_0_stall_1 <= io_in_r_bypass_8_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_1_data_1 <= io_in_r_bypass_8_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_1_load_store_1 <= io_in_r_bypass_8_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_1_df_is_ws_1 <= io_in_r_bypass_8_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_1_stall_1 <= io_in_r_bypass_8_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_2_data_1 <= io_in_r_bypass_8_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_2_load_store_1 <= io_in_r_bypass_8_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_2_df_is_ws_1 <= io_in_r_bypass_8_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_2_stall_1 <= io_in_r_bypass_8_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_3_data_1 <= io_in_r_bypass_8_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_3_load_store_1 <= io_in_r_bypass_8_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_3_df_is_ws_1 <= io_in_r_bypass_8_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_3_stall_1 <= io_in_r_bypass_8_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_0_data_1 <= io_in_r_bypass_9_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_0_load_store_1 <= io_in_r_bypass_9_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_0_df_is_ws_1 <= io_in_r_bypass_9_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_0_stall_1 <= io_in_r_bypass_9_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_1_data_1 <= io_in_r_bypass_9_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_1_load_store_1 <= io_in_r_bypass_9_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_1_df_is_ws_1 <= io_in_r_bypass_9_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_1_stall_1 <= io_in_r_bypass_9_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_2_data_1 <= io_in_r_bypass_9_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_2_load_store_1 <= io_in_r_bypass_9_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_2_df_is_ws_1 <= io_in_r_bypass_9_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_2_stall_1 <= io_in_r_bypass_9_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_3_data_1 <= io_in_r_bypass_9_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_3_load_store_1 <= io_in_r_bypass_9_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_3_df_is_ws_1 <= io_in_r_bypass_9_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_3_stall_1 <= io_in_r_bypass_9_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_0_data_1 <= io_in_r_bypass_10_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_0_load_store_1 <= io_in_r_bypass_10_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_0_df_is_ws_1 <= io_in_r_bypass_10_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_0_stall_1 <= io_in_r_bypass_10_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_1_data_1 <= io_in_r_bypass_10_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_1_load_store_1 <= io_in_r_bypass_10_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_1_df_is_ws_1 <= io_in_r_bypass_10_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_1_stall_1 <= io_in_r_bypass_10_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_2_data_1 <= io_in_r_bypass_10_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_2_load_store_1 <= io_in_r_bypass_10_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_2_df_is_ws_1 <= io_in_r_bypass_10_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_2_stall_1 <= io_in_r_bypass_10_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_3_data_1 <= io_in_r_bypass_10_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_3_load_store_1 <= io_in_r_bypass_10_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_3_df_is_ws_1 <= io_in_r_bypass_10_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_3_stall_1 <= io_in_r_bypass_10_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_0_data_1 <= io_in_r_bypass_11_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_0_load_store_1 <= io_in_r_bypass_11_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_0_df_is_ws_1 <= io_in_r_bypass_11_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_0_stall_1 <= io_in_r_bypass_11_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_1_data_1 <= io_in_r_bypass_11_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_1_load_store_1 <= io_in_r_bypass_11_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_1_df_is_ws_1 <= io_in_r_bypass_11_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_1_stall_1 <= io_in_r_bypass_11_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_2_data_1 <= io_in_r_bypass_11_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_2_load_store_1 <= io_in_r_bypass_11_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_2_df_is_ws_1 <= io_in_r_bypass_11_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_2_stall_1 <= io_in_r_bypass_11_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_3_data_1 <= io_in_r_bypass_11_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_3_load_store_1 <= io_in_r_bypass_11_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_3_df_is_ws_1 <= io_in_r_bypass_11_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_3_stall_1 <= io_in_r_bypass_11_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_0_data_1 <= io_in_r_bypass_12_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_0_load_store_1 <= io_in_r_bypass_12_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_0_df_is_ws_1 <= io_in_r_bypass_12_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_0_stall_1 <= io_in_r_bypass_12_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_1_data_1 <= io_in_r_bypass_12_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_1_load_store_1 <= io_in_r_bypass_12_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_1_df_is_ws_1 <= io_in_r_bypass_12_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_1_stall_1 <= io_in_r_bypass_12_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_2_data_1 <= io_in_r_bypass_12_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_2_load_store_1 <= io_in_r_bypass_12_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_2_df_is_ws_1 <= io_in_r_bypass_12_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_2_stall_1 <= io_in_r_bypass_12_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_3_data_1 <= io_in_r_bypass_12_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_3_load_store_1 <= io_in_r_bypass_12_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_3_df_is_ws_1 <= io_in_r_bypass_12_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_3_stall_1 <= io_in_r_bypass_12_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_0_data_1 <= io_in_r_bypass_13_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_0_load_store_1 <= io_in_r_bypass_13_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_0_df_is_ws_1 <= io_in_r_bypass_13_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_0_stall_1 <= io_in_r_bypass_13_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_1_data_1 <= io_in_r_bypass_13_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_1_load_store_1 <= io_in_r_bypass_13_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_1_df_is_ws_1 <= io_in_r_bypass_13_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_1_stall_1 <= io_in_r_bypass_13_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_2_data_1 <= io_in_r_bypass_13_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_2_load_store_1 <= io_in_r_bypass_13_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_2_df_is_ws_1 <= io_in_r_bypass_13_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_2_stall_1 <= io_in_r_bypass_13_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_3_data_1 <= io_in_r_bypass_13_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_3_load_store_1 <= io_in_r_bypass_13_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_3_df_is_ws_1 <= io_in_r_bypass_13_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_3_stall_1 <= io_in_r_bypass_13_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_0_data_1 <= io_in_r_bypass_14_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_0_load_store_1 <= io_in_r_bypass_14_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_0_df_is_ws_1 <= io_in_r_bypass_14_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_0_stall_1 <= io_in_r_bypass_14_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_1_data_1 <= io_in_r_bypass_14_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_1_load_store_1 <= io_in_r_bypass_14_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_1_df_is_ws_1 <= io_in_r_bypass_14_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_1_stall_1 <= io_in_r_bypass_14_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_2_data_1 <= io_in_r_bypass_14_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_2_load_store_1 <= io_in_r_bypass_14_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_2_df_is_ws_1 <= io_in_r_bypass_14_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_2_stall_1 <= io_in_r_bypass_14_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_3_data_1 <= io_in_r_bypass_14_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_3_load_store_1 <= io_in_r_bypass_14_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_3_df_is_ws_1 <= io_in_r_bypass_14_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_3_stall_1 <= io_in_r_bypass_14_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_0_data_1 <= io_in_r_bypass_15_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_0_load_store_1 <= io_in_r_bypass_15_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_0_df_is_ws_1 <= io_in_r_bypass_15_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_0_stall_1 <= io_in_r_bypass_15_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_1_data_1 <= io_in_r_bypass_15_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_1_load_store_1 <= io_in_r_bypass_15_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_1_df_is_ws_1 <= io_in_r_bypass_15_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_1_stall_1 <= io_in_r_bypass_15_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_2_data_1 <= io_in_r_bypass_15_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_2_load_store_1 <= io_in_r_bypass_15_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_2_df_is_ws_1 <= io_in_r_bypass_15_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_2_stall_1 <= io_in_r_bypass_15_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_3_data_1 <= io_in_r_bypass_15_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_3_load_store_1 <= io_in_r_bypass_15_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_3_df_is_ws_1 <= io_in_r_bypass_15_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_3_stall_1 <= io_in_r_bypass_15_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_0_data_1 <= io_in_r_bypass_16_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_0_load_store_1 <= io_in_r_bypass_16_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_0_df_is_ws_1 <= io_in_r_bypass_16_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_0_stall_1 <= io_in_r_bypass_16_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_1_data_1 <= io_in_r_bypass_16_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_1_load_store_1 <= io_in_r_bypass_16_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_1_df_is_ws_1 <= io_in_r_bypass_16_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_1_stall_1 <= io_in_r_bypass_16_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_2_data_1 <= io_in_r_bypass_16_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_2_load_store_1 <= io_in_r_bypass_16_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_2_df_is_ws_1 <= io_in_r_bypass_16_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_2_stall_1 <= io_in_r_bypass_16_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_3_data_1 <= io_in_r_bypass_16_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_3_load_store_1 <= io_in_r_bypass_16_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_3_df_is_ws_1 <= io_in_r_bypass_16_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_3_stall_1 <= io_in_r_bypass_16_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_0_data_1 <= io_in_r_bypass_17_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_0_load_store_1 <= io_in_r_bypass_17_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_0_df_is_ws_1 <= io_in_r_bypass_17_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_0_stall_1 <= io_in_r_bypass_17_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_1_data_1 <= io_in_r_bypass_17_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_1_load_store_1 <= io_in_r_bypass_17_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_1_df_is_ws_1 <= io_in_r_bypass_17_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_1_stall_1 <= io_in_r_bypass_17_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_2_data_1 <= io_in_r_bypass_17_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_2_load_store_1 <= io_in_r_bypass_17_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_2_df_is_ws_1 <= io_in_r_bypass_17_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_2_stall_1 <= io_in_r_bypass_17_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_3_data_1 <= io_in_r_bypass_17_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_3_load_store_1 <= io_in_r_bypass_17_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_3_df_is_ws_1 <= io_in_r_bypass_17_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_3_stall_1 <= io_in_r_bypass_17_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_0_data_1 <= io_in_r_bypass_18_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_0_load_store_1 <= io_in_r_bypass_18_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_0_df_is_ws_1 <= io_in_r_bypass_18_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_0_stall_1 <= io_in_r_bypass_18_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_1_data_1 <= io_in_r_bypass_18_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_1_load_store_1 <= io_in_r_bypass_18_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_1_df_is_ws_1 <= io_in_r_bypass_18_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_1_stall_1 <= io_in_r_bypass_18_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_2_data_1 <= io_in_r_bypass_18_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_2_load_store_1 <= io_in_r_bypass_18_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_2_df_is_ws_1 <= io_in_r_bypass_18_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_2_stall_1 <= io_in_r_bypass_18_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_3_data_1 <= io_in_r_bypass_18_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_3_load_store_1 <= io_in_r_bypass_18_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_3_df_is_ws_1 <= io_in_r_bypass_18_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_3_stall_1 <= io_in_r_bypass_18_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_0_data_1 <= io_in_r_bypass_19_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_0_load_store_1 <= io_in_r_bypass_19_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_0_df_is_ws_1 <= io_in_r_bypass_19_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_0_stall_1 <= io_in_r_bypass_19_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_1_data_1 <= io_in_r_bypass_19_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_1_load_store_1 <= io_in_r_bypass_19_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_1_df_is_ws_1 <= io_in_r_bypass_19_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_1_stall_1 <= io_in_r_bypass_19_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_2_data_1 <= io_in_r_bypass_19_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_2_load_store_1 <= io_in_r_bypass_19_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_2_df_is_ws_1 <= io_in_r_bypass_19_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_2_stall_1 <= io_in_r_bypass_19_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_3_data_1 <= io_in_r_bypass_19_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_3_load_store_1 <= io_in_r_bypass_19_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_3_df_is_ws_1 <= io_in_r_bypass_19_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_3_stall_1 <= io_in_r_bypass_19_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_0_data_1 <= io_in_r_bypass_20_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_0_load_store_1 <= io_in_r_bypass_20_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_0_df_is_ws_1 <= io_in_r_bypass_20_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_0_stall_1 <= io_in_r_bypass_20_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_1_data_1 <= io_in_r_bypass_20_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_1_load_store_1 <= io_in_r_bypass_20_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_1_df_is_ws_1 <= io_in_r_bypass_20_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_1_stall_1 <= io_in_r_bypass_20_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_2_data_1 <= io_in_r_bypass_20_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_2_load_store_1 <= io_in_r_bypass_20_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_2_df_is_ws_1 <= io_in_r_bypass_20_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_2_stall_1 <= io_in_r_bypass_20_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_3_data_1 <= io_in_r_bypass_20_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_3_load_store_1 <= io_in_r_bypass_20_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_3_df_is_ws_1 <= io_in_r_bypass_20_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_3_stall_1 <= io_in_r_bypass_20_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_0_data_1 <= io_in_r_bypass_21_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_0_load_store_1 <= io_in_r_bypass_21_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_0_df_is_ws_1 <= io_in_r_bypass_21_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_0_stall_1 <= io_in_r_bypass_21_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_1_data_1 <= io_in_r_bypass_21_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_1_load_store_1 <= io_in_r_bypass_21_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_1_df_is_ws_1 <= io_in_r_bypass_21_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_1_stall_1 <= io_in_r_bypass_21_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_2_data_1 <= io_in_r_bypass_21_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_2_load_store_1 <= io_in_r_bypass_21_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_2_df_is_ws_1 <= io_in_r_bypass_21_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_2_stall_1 <= io_in_r_bypass_21_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_3_data_1 <= io_in_r_bypass_21_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_3_load_store_1 <= io_in_r_bypass_21_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_3_df_is_ws_1 <= io_in_r_bypass_21_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_3_stall_1 <= io_in_r_bypass_21_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_0_data_1 <= io_in_r_bypass_22_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_0_load_store_1 <= io_in_r_bypass_22_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_0_df_is_ws_1 <= io_in_r_bypass_22_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_0_stall_1 <= io_in_r_bypass_22_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_1_data_1 <= io_in_r_bypass_22_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_1_load_store_1 <= io_in_r_bypass_22_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_1_df_is_ws_1 <= io_in_r_bypass_22_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_1_stall_1 <= io_in_r_bypass_22_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_2_data_1 <= io_in_r_bypass_22_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_2_load_store_1 <= io_in_r_bypass_22_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_2_df_is_ws_1 <= io_in_r_bypass_22_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_2_stall_1 <= io_in_r_bypass_22_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_3_data_1 <= io_in_r_bypass_22_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_3_load_store_1 <= io_in_r_bypass_22_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_3_df_is_ws_1 <= io_in_r_bypass_22_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_3_stall_1 <= io_in_r_bypass_22_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_0_data_1 <= io_in_r_bypass_23_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_0_load_store_1 <= io_in_r_bypass_23_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_0_df_is_ws_1 <= io_in_r_bypass_23_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_0_stall_1 <= io_in_r_bypass_23_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_1_data_1 <= io_in_r_bypass_23_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_1_load_store_1 <= io_in_r_bypass_23_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_1_df_is_ws_1 <= io_in_r_bypass_23_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_1_stall_1 <= io_in_r_bypass_23_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_2_data_1 <= io_in_r_bypass_23_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_2_load_store_1 <= io_in_r_bypass_23_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_2_df_is_ws_1 <= io_in_r_bypass_23_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_2_stall_1 <= io_in_r_bypass_23_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_3_data_1 <= io_in_r_bypass_23_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_3_load_store_1 <= io_in_r_bypass_23_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_3_df_is_ws_1 <= io_in_r_bypass_23_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_3_stall_1 <= io_in_r_bypass_23_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_0_data_1 <= io_in_r_bypass_24_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_0_load_store_1 <= io_in_r_bypass_24_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_0_df_is_ws_1 <= io_in_r_bypass_24_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_0_stall_1 <= io_in_r_bypass_24_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_1_data_1 <= io_in_r_bypass_24_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_1_load_store_1 <= io_in_r_bypass_24_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_1_df_is_ws_1 <= io_in_r_bypass_24_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_1_stall_1 <= io_in_r_bypass_24_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_2_data_1 <= io_in_r_bypass_24_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_2_load_store_1 <= io_in_r_bypass_24_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_2_df_is_ws_1 <= io_in_r_bypass_24_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_2_stall_1 <= io_in_r_bypass_24_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_3_data_1 <= io_in_r_bypass_24_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_3_load_store_1 <= io_in_r_bypass_24_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_3_df_is_ws_1 <= io_in_r_bypass_24_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_3_stall_1 <= io_in_r_bypass_24_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_0_data_1 <= io_in_r_bypass_25_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_0_load_store_1 <= io_in_r_bypass_25_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_0_df_is_ws_1 <= io_in_r_bypass_25_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_0_stall_1 <= io_in_r_bypass_25_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_1_data_1 <= io_in_r_bypass_25_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_1_load_store_1 <= io_in_r_bypass_25_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_1_df_is_ws_1 <= io_in_r_bypass_25_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_1_stall_1 <= io_in_r_bypass_25_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_2_data_1 <= io_in_r_bypass_25_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_2_load_store_1 <= io_in_r_bypass_25_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_2_df_is_ws_1 <= io_in_r_bypass_25_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_2_stall_1 <= io_in_r_bypass_25_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_3_data_1 <= io_in_r_bypass_25_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_3_load_store_1 <= io_in_r_bypass_25_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_3_df_is_ws_1 <= io_in_r_bypass_25_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_3_stall_1 <= io_in_r_bypass_25_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_0_data_1 <= io_in_r_bypass_26_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_0_load_store_1 <= io_in_r_bypass_26_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_0_df_is_ws_1 <= io_in_r_bypass_26_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_0_stall_1 <= io_in_r_bypass_26_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_1_data_1 <= io_in_r_bypass_26_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_1_load_store_1 <= io_in_r_bypass_26_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_1_df_is_ws_1 <= io_in_r_bypass_26_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_1_stall_1 <= io_in_r_bypass_26_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_2_data_1 <= io_in_r_bypass_26_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_2_load_store_1 <= io_in_r_bypass_26_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_2_df_is_ws_1 <= io_in_r_bypass_26_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_2_stall_1 <= io_in_r_bypass_26_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_3_data_1 <= io_in_r_bypass_26_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_3_load_store_1 <= io_in_r_bypass_26_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_3_df_is_ws_1 <= io_in_r_bypass_26_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_3_stall_1 <= io_in_r_bypass_26_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_0_data_1 <= io_in_r_bypass_27_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_0_load_store_1 <= io_in_r_bypass_27_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_0_df_is_ws_1 <= io_in_r_bypass_27_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_0_stall_1 <= io_in_r_bypass_27_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_1_data_1 <= io_in_r_bypass_27_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_1_load_store_1 <= io_in_r_bypass_27_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_1_df_is_ws_1 <= io_in_r_bypass_27_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_1_stall_1 <= io_in_r_bypass_27_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_2_data_1 <= io_in_r_bypass_27_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_2_load_store_1 <= io_in_r_bypass_27_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_2_df_is_ws_1 <= io_in_r_bypass_27_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_2_stall_1 <= io_in_r_bypass_27_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_3_data_1 <= io_in_r_bypass_27_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_3_load_store_1 <= io_in_r_bypass_27_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_3_df_is_ws_1 <= io_in_r_bypass_27_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_3_stall_1 <= io_in_r_bypass_27_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_0_data_1 <= io_in_r_bypass_28_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_0_load_store_1 <= io_in_r_bypass_28_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_0_df_is_ws_1 <= io_in_r_bypass_28_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_0_stall_1 <= io_in_r_bypass_28_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_1_data_1 <= io_in_r_bypass_28_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_1_load_store_1 <= io_in_r_bypass_28_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_1_df_is_ws_1 <= io_in_r_bypass_28_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_1_stall_1 <= io_in_r_bypass_28_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_2_data_1 <= io_in_r_bypass_28_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_2_load_store_1 <= io_in_r_bypass_28_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_2_df_is_ws_1 <= io_in_r_bypass_28_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_2_stall_1 <= io_in_r_bypass_28_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_3_data_1 <= io_in_r_bypass_28_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_3_load_store_1 <= io_in_r_bypass_28_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_3_df_is_ws_1 <= io_in_r_bypass_28_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_3_stall_1 <= io_in_r_bypass_28_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_0_data_1 <= io_in_r_bypass_29_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_0_load_store_1 <= io_in_r_bypass_29_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_0_df_is_ws_1 <= io_in_r_bypass_29_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_0_stall_1 <= io_in_r_bypass_29_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_1_data_1 <= io_in_r_bypass_29_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_1_load_store_1 <= io_in_r_bypass_29_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_1_df_is_ws_1 <= io_in_r_bypass_29_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_1_stall_1 <= io_in_r_bypass_29_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_2_data_1 <= io_in_r_bypass_29_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_2_load_store_1 <= io_in_r_bypass_29_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_2_df_is_ws_1 <= io_in_r_bypass_29_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_2_stall_1 <= io_in_r_bypass_29_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_3_data_1 <= io_in_r_bypass_29_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_3_load_store_1 <= io_in_r_bypass_29_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_3_df_is_ws_1 <= io_in_r_bypass_29_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_3_stall_1 <= io_in_r_bypass_29_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_0_data_1 <= io_in_r_bypass_30_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_0_load_store_1 <= io_in_r_bypass_30_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_0_df_is_ws_1 <= io_in_r_bypass_30_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_0_stall_1 <= io_in_r_bypass_30_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_1_data_1 <= io_in_r_bypass_30_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_1_load_store_1 <= io_in_r_bypass_30_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_1_df_is_ws_1 <= io_in_r_bypass_30_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_1_stall_1 <= io_in_r_bypass_30_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_2_data_1 <= io_in_r_bypass_30_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_2_load_store_1 <= io_in_r_bypass_30_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_2_df_is_ws_1 <= io_in_r_bypass_30_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_2_stall_1 <= io_in_r_bypass_30_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_3_data_1 <= io_in_r_bypass_30_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_3_load_store_1 <= io_in_r_bypass_30_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_3_df_is_ws_1 <= io_in_r_bypass_30_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_3_stall_1 <= io_in_r_bypass_30_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_0_data_1 <= io_in_r_bypass_31_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_0_load_store_1 <= io_in_r_bypass_31_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_0_df_is_ws_1 <= io_in_r_bypass_31_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_0_stall_1 <= io_in_r_bypass_31_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_1_data_1 <= io_in_r_bypass_31_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_1_load_store_1 <= io_in_r_bypass_31_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_1_df_is_ws_1 <= io_in_r_bypass_31_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_1_stall_1 <= io_in_r_bypass_31_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_2_data_1 <= io_in_r_bypass_31_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_2_load_store_1 <= io_in_r_bypass_31_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_2_df_is_ws_1 <= io_in_r_bypass_31_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_2_stall_1 <= io_in_r_bypass_31_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_3_data_1 <= io_in_r_bypass_31_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_3_load_store_1 <= io_in_r_bypass_31_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_3_df_is_ws_1 <= io_in_r_bypass_31_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_3_stall_1 <= io_in_r_bypass_31_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_0_data_2 <= io_in_r_bypass_0_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_0_load_store_2 <= io_in_r_bypass_0_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_0_df_is_ws_2 <= io_in_r_bypass_0_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_0_stall_2 <= io_in_r_bypass_0_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_1_data_2 <= io_in_r_bypass_0_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_1_load_store_2 <= io_in_r_bypass_0_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_1_df_is_ws_2 <= io_in_r_bypass_0_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_1_stall_2 <= io_in_r_bypass_0_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_2_data_2 <= io_in_r_bypass_0_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_2_load_store_2 <= io_in_r_bypass_0_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_2_df_is_ws_2 <= io_in_r_bypass_0_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_2_stall_2 <= io_in_r_bypass_0_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_3_data_2 <= io_in_r_bypass_0_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_3_load_store_2 <= io_in_r_bypass_0_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_3_df_is_ws_2 <= io_in_r_bypass_0_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_3_stall_2 <= io_in_r_bypass_0_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_0_data_2 <= io_in_r_bypass_1_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_0_load_store_2 <= io_in_r_bypass_1_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_0_df_is_ws_2 <= io_in_r_bypass_1_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_0_stall_2 <= io_in_r_bypass_1_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_1_data_2 <= io_in_r_bypass_1_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_1_load_store_2 <= io_in_r_bypass_1_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_1_df_is_ws_2 <= io_in_r_bypass_1_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_1_stall_2 <= io_in_r_bypass_1_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_2_data_2 <= io_in_r_bypass_1_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_2_load_store_2 <= io_in_r_bypass_1_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_2_df_is_ws_2 <= io_in_r_bypass_1_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_2_stall_2 <= io_in_r_bypass_1_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_3_data_2 <= io_in_r_bypass_1_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_3_load_store_2 <= io_in_r_bypass_1_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_3_df_is_ws_2 <= io_in_r_bypass_1_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_3_stall_2 <= io_in_r_bypass_1_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_0_data_2 <= io_in_r_bypass_2_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_0_load_store_2 <= io_in_r_bypass_2_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_0_df_is_ws_2 <= io_in_r_bypass_2_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_0_stall_2 <= io_in_r_bypass_2_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_1_data_2 <= io_in_r_bypass_2_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_1_load_store_2 <= io_in_r_bypass_2_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_1_df_is_ws_2 <= io_in_r_bypass_2_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_1_stall_2 <= io_in_r_bypass_2_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_2_data_2 <= io_in_r_bypass_2_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_2_load_store_2 <= io_in_r_bypass_2_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_2_df_is_ws_2 <= io_in_r_bypass_2_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_2_stall_2 <= io_in_r_bypass_2_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_3_data_2 <= io_in_r_bypass_2_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_3_load_store_2 <= io_in_r_bypass_2_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_3_df_is_ws_2 <= io_in_r_bypass_2_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_3_stall_2 <= io_in_r_bypass_2_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_0_data_2 <= io_in_r_bypass_3_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_0_load_store_2 <= io_in_r_bypass_3_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_0_df_is_ws_2 <= io_in_r_bypass_3_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_0_stall_2 <= io_in_r_bypass_3_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_1_data_2 <= io_in_r_bypass_3_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_1_load_store_2 <= io_in_r_bypass_3_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_1_df_is_ws_2 <= io_in_r_bypass_3_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_1_stall_2 <= io_in_r_bypass_3_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_2_data_2 <= io_in_r_bypass_3_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_2_load_store_2 <= io_in_r_bypass_3_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_2_df_is_ws_2 <= io_in_r_bypass_3_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_2_stall_2 <= io_in_r_bypass_3_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_3_data_2 <= io_in_r_bypass_3_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_3_load_store_2 <= io_in_r_bypass_3_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_3_df_is_ws_2 <= io_in_r_bypass_3_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_3_stall_2 <= io_in_r_bypass_3_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_0_data_2 <= io_in_r_bypass_4_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_0_load_store_2 <= io_in_r_bypass_4_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_0_df_is_ws_2 <= io_in_r_bypass_4_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_0_stall_2 <= io_in_r_bypass_4_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_1_data_2 <= io_in_r_bypass_4_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_1_load_store_2 <= io_in_r_bypass_4_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_1_df_is_ws_2 <= io_in_r_bypass_4_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_1_stall_2 <= io_in_r_bypass_4_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_2_data_2 <= io_in_r_bypass_4_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_2_load_store_2 <= io_in_r_bypass_4_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_2_df_is_ws_2 <= io_in_r_bypass_4_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_2_stall_2 <= io_in_r_bypass_4_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_3_data_2 <= io_in_r_bypass_4_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_3_load_store_2 <= io_in_r_bypass_4_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_3_df_is_ws_2 <= io_in_r_bypass_4_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_3_stall_2 <= io_in_r_bypass_4_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_0_data_2 <= io_in_r_bypass_5_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_0_load_store_2 <= io_in_r_bypass_5_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_0_df_is_ws_2 <= io_in_r_bypass_5_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_0_stall_2 <= io_in_r_bypass_5_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_1_data_2 <= io_in_r_bypass_5_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_1_load_store_2 <= io_in_r_bypass_5_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_1_df_is_ws_2 <= io_in_r_bypass_5_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_1_stall_2 <= io_in_r_bypass_5_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_2_data_2 <= io_in_r_bypass_5_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_2_load_store_2 <= io_in_r_bypass_5_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_2_df_is_ws_2 <= io_in_r_bypass_5_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_2_stall_2 <= io_in_r_bypass_5_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_3_data_2 <= io_in_r_bypass_5_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_3_load_store_2 <= io_in_r_bypass_5_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_3_df_is_ws_2 <= io_in_r_bypass_5_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_3_stall_2 <= io_in_r_bypass_5_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_0_data_2 <= io_in_r_bypass_6_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_0_load_store_2 <= io_in_r_bypass_6_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_0_df_is_ws_2 <= io_in_r_bypass_6_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_0_stall_2 <= io_in_r_bypass_6_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_1_data_2 <= io_in_r_bypass_6_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_1_load_store_2 <= io_in_r_bypass_6_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_1_df_is_ws_2 <= io_in_r_bypass_6_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_1_stall_2 <= io_in_r_bypass_6_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_2_data_2 <= io_in_r_bypass_6_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_2_load_store_2 <= io_in_r_bypass_6_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_2_df_is_ws_2 <= io_in_r_bypass_6_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_2_stall_2 <= io_in_r_bypass_6_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_3_data_2 <= io_in_r_bypass_6_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_3_load_store_2 <= io_in_r_bypass_6_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_3_df_is_ws_2 <= io_in_r_bypass_6_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_3_stall_2 <= io_in_r_bypass_6_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_0_data_2 <= io_in_r_bypass_7_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_0_load_store_2 <= io_in_r_bypass_7_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_0_df_is_ws_2 <= io_in_r_bypass_7_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_0_stall_2 <= io_in_r_bypass_7_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_1_data_2 <= io_in_r_bypass_7_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_1_load_store_2 <= io_in_r_bypass_7_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_1_df_is_ws_2 <= io_in_r_bypass_7_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_1_stall_2 <= io_in_r_bypass_7_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_2_data_2 <= io_in_r_bypass_7_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_2_load_store_2 <= io_in_r_bypass_7_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_2_df_is_ws_2 <= io_in_r_bypass_7_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_2_stall_2 <= io_in_r_bypass_7_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_3_data_2 <= io_in_r_bypass_7_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_3_load_store_2 <= io_in_r_bypass_7_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_3_df_is_ws_2 <= io_in_r_bypass_7_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_3_stall_2 <= io_in_r_bypass_7_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_0_data_2 <= io_in_r_bypass_8_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_0_load_store_2 <= io_in_r_bypass_8_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_0_df_is_ws_2 <= io_in_r_bypass_8_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_0_stall_2 <= io_in_r_bypass_8_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_1_data_2 <= io_in_r_bypass_8_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_1_load_store_2 <= io_in_r_bypass_8_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_1_df_is_ws_2 <= io_in_r_bypass_8_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_1_stall_2 <= io_in_r_bypass_8_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_2_data_2 <= io_in_r_bypass_8_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_2_load_store_2 <= io_in_r_bypass_8_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_2_df_is_ws_2 <= io_in_r_bypass_8_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_2_stall_2 <= io_in_r_bypass_8_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_3_data_2 <= io_in_r_bypass_8_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_3_load_store_2 <= io_in_r_bypass_8_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_3_df_is_ws_2 <= io_in_r_bypass_8_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_3_stall_2 <= io_in_r_bypass_8_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_0_data_2 <= io_in_r_bypass_9_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_0_load_store_2 <= io_in_r_bypass_9_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_0_df_is_ws_2 <= io_in_r_bypass_9_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_0_stall_2 <= io_in_r_bypass_9_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_1_data_2 <= io_in_r_bypass_9_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_1_load_store_2 <= io_in_r_bypass_9_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_1_df_is_ws_2 <= io_in_r_bypass_9_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_1_stall_2 <= io_in_r_bypass_9_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_2_data_2 <= io_in_r_bypass_9_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_2_load_store_2 <= io_in_r_bypass_9_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_2_df_is_ws_2 <= io_in_r_bypass_9_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_2_stall_2 <= io_in_r_bypass_9_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_3_data_2 <= io_in_r_bypass_9_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_3_load_store_2 <= io_in_r_bypass_9_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_3_df_is_ws_2 <= io_in_r_bypass_9_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_3_stall_2 <= io_in_r_bypass_9_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_0_data_2 <= io_in_r_bypass_10_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_0_load_store_2 <= io_in_r_bypass_10_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_0_df_is_ws_2 <= io_in_r_bypass_10_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_0_stall_2 <= io_in_r_bypass_10_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_1_data_2 <= io_in_r_bypass_10_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_1_load_store_2 <= io_in_r_bypass_10_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_1_df_is_ws_2 <= io_in_r_bypass_10_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_1_stall_2 <= io_in_r_bypass_10_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_2_data_2 <= io_in_r_bypass_10_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_2_load_store_2 <= io_in_r_bypass_10_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_2_df_is_ws_2 <= io_in_r_bypass_10_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_2_stall_2 <= io_in_r_bypass_10_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_3_data_2 <= io_in_r_bypass_10_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_3_load_store_2 <= io_in_r_bypass_10_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_3_df_is_ws_2 <= io_in_r_bypass_10_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_3_stall_2 <= io_in_r_bypass_10_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_0_data_2 <= io_in_r_bypass_11_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_0_load_store_2 <= io_in_r_bypass_11_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_0_df_is_ws_2 <= io_in_r_bypass_11_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_0_stall_2 <= io_in_r_bypass_11_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_1_data_2 <= io_in_r_bypass_11_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_1_load_store_2 <= io_in_r_bypass_11_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_1_df_is_ws_2 <= io_in_r_bypass_11_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_1_stall_2 <= io_in_r_bypass_11_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_2_data_2 <= io_in_r_bypass_11_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_2_load_store_2 <= io_in_r_bypass_11_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_2_df_is_ws_2 <= io_in_r_bypass_11_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_2_stall_2 <= io_in_r_bypass_11_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_3_data_2 <= io_in_r_bypass_11_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_3_load_store_2 <= io_in_r_bypass_11_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_3_df_is_ws_2 <= io_in_r_bypass_11_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_3_stall_2 <= io_in_r_bypass_11_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_0_data_2 <= io_in_r_bypass_12_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_0_load_store_2 <= io_in_r_bypass_12_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_0_df_is_ws_2 <= io_in_r_bypass_12_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_0_stall_2 <= io_in_r_bypass_12_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_1_data_2 <= io_in_r_bypass_12_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_1_load_store_2 <= io_in_r_bypass_12_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_1_df_is_ws_2 <= io_in_r_bypass_12_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_1_stall_2 <= io_in_r_bypass_12_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_2_data_2 <= io_in_r_bypass_12_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_2_load_store_2 <= io_in_r_bypass_12_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_2_df_is_ws_2 <= io_in_r_bypass_12_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_2_stall_2 <= io_in_r_bypass_12_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_3_data_2 <= io_in_r_bypass_12_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_3_load_store_2 <= io_in_r_bypass_12_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_3_df_is_ws_2 <= io_in_r_bypass_12_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_3_stall_2 <= io_in_r_bypass_12_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_0_data_2 <= io_in_r_bypass_13_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_0_load_store_2 <= io_in_r_bypass_13_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_0_df_is_ws_2 <= io_in_r_bypass_13_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_0_stall_2 <= io_in_r_bypass_13_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_1_data_2 <= io_in_r_bypass_13_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_1_load_store_2 <= io_in_r_bypass_13_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_1_df_is_ws_2 <= io_in_r_bypass_13_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_1_stall_2 <= io_in_r_bypass_13_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_2_data_2 <= io_in_r_bypass_13_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_2_load_store_2 <= io_in_r_bypass_13_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_2_df_is_ws_2 <= io_in_r_bypass_13_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_2_stall_2 <= io_in_r_bypass_13_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_3_data_2 <= io_in_r_bypass_13_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_3_load_store_2 <= io_in_r_bypass_13_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_3_df_is_ws_2 <= io_in_r_bypass_13_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_3_stall_2 <= io_in_r_bypass_13_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_0_data_2 <= io_in_r_bypass_14_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_0_load_store_2 <= io_in_r_bypass_14_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_0_df_is_ws_2 <= io_in_r_bypass_14_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_0_stall_2 <= io_in_r_bypass_14_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_1_data_2 <= io_in_r_bypass_14_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_1_load_store_2 <= io_in_r_bypass_14_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_1_df_is_ws_2 <= io_in_r_bypass_14_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_1_stall_2 <= io_in_r_bypass_14_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_2_data_2 <= io_in_r_bypass_14_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_2_load_store_2 <= io_in_r_bypass_14_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_2_df_is_ws_2 <= io_in_r_bypass_14_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_2_stall_2 <= io_in_r_bypass_14_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_3_data_2 <= io_in_r_bypass_14_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_3_load_store_2 <= io_in_r_bypass_14_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_3_df_is_ws_2 <= io_in_r_bypass_14_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_3_stall_2 <= io_in_r_bypass_14_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_0_data_2 <= io_in_r_bypass_15_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_0_load_store_2 <= io_in_r_bypass_15_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_0_df_is_ws_2 <= io_in_r_bypass_15_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_0_stall_2 <= io_in_r_bypass_15_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_1_data_2 <= io_in_r_bypass_15_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_1_load_store_2 <= io_in_r_bypass_15_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_1_df_is_ws_2 <= io_in_r_bypass_15_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_1_stall_2 <= io_in_r_bypass_15_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_2_data_2 <= io_in_r_bypass_15_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_2_load_store_2 <= io_in_r_bypass_15_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_2_df_is_ws_2 <= io_in_r_bypass_15_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_2_stall_2 <= io_in_r_bypass_15_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_3_data_2 <= io_in_r_bypass_15_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_3_load_store_2 <= io_in_r_bypass_15_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_3_df_is_ws_2 <= io_in_r_bypass_15_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_3_stall_2 <= io_in_r_bypass_15_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_0_data_2 <= io_in_r_bypass_16_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_0_load_store_2 <= io_in_r_bypass_16_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_0_df_is_ws_2 <= io_in_r_bypass_16_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_0_stall_2 <= io_in_r_bypass_16_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_1_data_2 <= io_in_r_bypass_16_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_1_load_store_2 <= io_in_r_bypass_16_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_1_df_is_ws_2 <= io_in_r_bypass_16_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_1_stall_2 <= io_in_r_bypass_16_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_2_data_2 <= io_in_r_bypass_16_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_2_load_store_2 <= io_in_r_bypass_16_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_2_df_is_ws_2 <= io_in_r_bypass_16_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_2_stall_2 <= io_in_r_bypass_16_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_3_data_2 <= io_in_r_bypass_16_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_3_load_store_2 <= io_in_r_bypass_16_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_3_df_is_ws_2 <= io_in_r_bypass_16_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_3_stall_2 <= io_in_r_bypass_16_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_0_data_2 <= io_in_r_bypass_17_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_0_load_store_2 <= io_in_r_bypass_17_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_0_df_is_ws_2 <= io_in_r_bypass_17_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_0_stall_2 <= io_in_r_bypass_17_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_1_data_2 <= io_in_r_bypass_17_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_1_load_store_2 <= io_in_r_bypass_17_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_1_df_is_ws_2 <= io_in_r_bypass_17_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_1_stall_2 <= io_in_r_bypass_17_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_2_data_2 <= io_in_r_bypass_17_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_2_load_store_2 <= io_in_r_bypass_17_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_2_df_is_ws_2 <= io_in_r_bypass_17_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_2_stall_2 <= io_in_r_bypass_17_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_3_data_2 <= io_in_r_bypass_17_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_3_load_store_2 <= io_in_r_bypass_17_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_3_df_is_ws_2 <= io_in_r_bypass_17_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_3_stall_2 <= io_in_r_bypass_17_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_0_data_2 <= io_in_r_bypass_18_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_0_load_store_2 <= io_in_r_bypass_18_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_0_df_is_ws_2 <= io_in_r_bypass_18_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_0_stall_2 <= io_in_r_bypass_18_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_1_data_2 <= io_in_r_bypass_18_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_1_load_store_2 <= io_in_r_bypass_18_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_1_df_is_ws_2 <= io_in_r_bypass_18_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_1_stall_2 <= io_in_r_bypass_18_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_2_data_2 <= io_in_r_bypass_18_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_2_load_store_2 <= io_in_r_bypass_18_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_2_df_is_ws_2 <= io_in_r_bypass_18_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_2_stall_2 <= io_in_r_bypass_18_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_3_data_2 <= io_in_r_bypass_18_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_3_load_store_2 <= io_in_r_bypass_18_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_3_df_is_ws_2 <= io_in_r_bypass_18_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_3_stall_2 <= io_in_r_bypass_18_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_0_data_2 <= io_in_r_bypass_19_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_0_load_store_2 <= io_in_r_bypass_19_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_0_df_is_ws_2 <= io_in_r_bypass_19_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_0_stall_2 <= io_in_r_bypass_19_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_1_data_2 <= io_in_r_bypass_19_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_1_load_store_2 <= io_in_r_bypass_19_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_1_df_is_ws_2 <= io_in_r_bypass_19_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_1_stall_2 <= io_in_r_bypass_19_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_2_data_2 <= io_in_r_bypass_19_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_2_load_store_2 <= io_in_r_bypass_19_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_2_df_is_ws_2 <= io_in_r_bypass_19_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_2_stall_2 <= io_in_r_bypass_19_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_3_data_2 <= io_in_r_bypass_19_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_3_load_store_2 <= io_in_r_bypass_19_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_3_df_is_ws_2 <= io_in_r_bypass_19_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_3_stall_2 <= io_in_r_bypass_19_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_0_data_2 <= io_in_r_bypass_20_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_0_load_store_2 <= io_in_r_bypass_20_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_0_df_is_ws_2 <= io_in_r_bypass_20_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_0_stall_2 <= io_in_r_bypass_20_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_1_data_2 <= io_in_r_bypass_20_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_1_load_store_2 <= io_in_r_bypass_20_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_1_df_is_ws_2 <= io_in_r_bypass_20_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_1_stall_2 <= io_in_r_bypass_20_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_2_data_2 <= io_in_r_bypass_20_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_2_load_store_2 <= io_in_r_bypass_20_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_2_df_is_ws_2 <= io_in_r_bypass_20_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_2_stall_2 <= io_in_r_bypass_20_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_3_data_2 <= io_in_r_bypass_20_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_3_load_store_2 <= io_in_r_bypass_20_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_3_df_is_ws_2 <= io_in_r_bypass_20_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_3_stall_2 <= io_in_r_bypass_20_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_0_data_2 <= io_in_r_bypass_21_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_0_load_store_2 <= io_in_r_bypass_21_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_0_df_is_ws_2 <= io_in_r_bypass_21_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_0_stall_2 <= io_in_r_bypass_21_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_1_data_2 <= io_in_r_bypass_21_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_1_load_store_2 <= io_in_r_bypass_21_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_1_df_is_ws_2 <= io_in_r_bypass_21_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_1_stall_2 <= io_in_r_bypass_21_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_2_data_2 <= io_in_r_bypass_21_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_2_load_store_2 <= io_in_r_bypass_21_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_2_df_is_ws_2 <= io_in_r_bypass_21_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_2_stall_2 <= io_in_r_bypass_21_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_3_data_2 <= io_in_r_bypass_21_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_3_load_store_2 <= io_in_r_bypass_21_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_3_df_is_ws_2 <= io_in_r_bypass_21_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_3_stall_2 <= io_in_r_bypass_21_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_0_data_2 <= io_in_r_bypass_22_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_0_load_store_2 <= io_in_r_bypass_22_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_0_df_is_ws_2 <= io_in_r_bypass_22_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_0_stall_2 <= io_in_r_bypass_22_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_1_data_2 <= io_in_r_bypass_22_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_1_load_store_2 <= io_in_r_bypass_22_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_1_df_is_ws_2 <= io_in_r_bypass_22_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_1_stall_2 <= io_in_r_bypass_22_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_2_data_2 <= io_in_r_bypass_22_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_2_load_store_2 <= io_in_r_bypass_22_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_2_df_is_ws_2 <= io_in_r_bypass_22_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_2_stall_2 <= io_in_r_bypass_22_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_3_data_2 <= io_in_r_bypass_22_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_3_load_store_2 <= io_in_r_bypass_22_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_3_df_is_ws_2 <= io_in_r_bypass_22_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_3_stall_2 <= io_in_r_bypass_22_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_0_data_2 <= io_in_r_bypass_23_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_0_load_store_2 <= io_in_r_bypass_23_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_0_df_is_ws_2 <= io_in_r_bypass_23_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_0_stall_2 <= io_in_r_bypass_23_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_1_data_2 <= io_in_r_bypass_23_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_1_load_store_2 <= io_in_r_bypass_23_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_1_df_is_ws_2 <= io_in_r_bypass_23_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_1_stall_2 <= io_in_r_bypass_23_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_2_data_2 <= io_in_r_bypass_23_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_2_load_store_2 <= io_in_r_bypass_23_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_2_df_is_ws_2 <= io_in_r_bypass_23_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_2_stall_2 <= io_in_r_bypass_23_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_3_data_2 <= io_in_r_bypass_23_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_3_load_store_2 <= io_in_r_bypass_23_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_3_df_is_ws_2 <= io_in_r_bypass_23_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_3_stall_2 <= io_in_r_bypass_23_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_0_data_2 <= io_in_r_bypass_24_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_0_load_store_2 <= io_in_r_bypass_24_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_0_df_is_ws_2 <= io_in_r_bypass_24_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_0_stall_2 <= io_in_r_bypass_24_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_1_data_2 <= io_in_r_bypass_24_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_1_load_store_2 <= io_in_r_bypass_24_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_1_df_is_ws_2 <= io_in_r_bypass_24_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_1_stall_2 <= io_in_r_bypass_24_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_2_data_2 <= io_in_r_bypass_24_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_2_load_store_2 <= io_in_r_bypass_24_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_2_df_is_ws_2 <= io_in_r_bypass_24_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_2_stall_2 <= io_in_r_bypass_24_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_3_data_2 <= io_in_r_bypass_24_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_3_load_store_2 <= io_in_r_bypass_24_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_3_df_is_ws_2 <= io_in_r_bypass_24_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_3_stall_2 <= io_in_r_bypass_24_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_0_data_2 <= io_in_r_bypass_25_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_0_load_store_2 <= io_in_r_bypass_25_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_0_df_is_ws_2 <= io_in_r_bypass_25_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_0_stall_2 <= io_in_r_bypass_25_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_1_data_2 <= io_in_r_bypass_25_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_1_load_store_2 <= io_in_r_bypass_25_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_1_df_is_ws_2 <= io_in_r_bypass_25_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_1_stall_2 <= io_in_r_bypass_25_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_2_data_2 <= io_in_r_bypass_25_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_2_load_store_2 <= io_in_r_bypass_25_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_2_df_is_ws_2 <= io_in_r_bypass_25_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_2_stall_2 <= io_in_r_bypass_25_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_3_data_2 <= io_in_r_bypass_25_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_3_load_store_2 <= io_in_r_bypass_25_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_3_df_is_ws_2 <= io_in_r_bypass_25_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_3_stall_2 <= io_in_r_bypass_25_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_0_data_2 <= io_in_r_bypass_26_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_0_load_store_2 <= io_in_r_bypass_26_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_0_df_is_ws_2 <= io_in_r_bypass_26_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_0_stall_2 <= io_in_r_bypass_26_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_1_data_2 <= io_in_r_bypass_26_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_1_load_store_2 <= io_in_r_bypass_26_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_1_df_is_ws_2 <= io_in_r_bypass_26_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_1_stall_2 <= io_in_r_bypass_26_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_2_data_2 <= io_in_r_bypass_26_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_2_load_store_2 <= io_in_r_bypass_26_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_2_df_is_ws_2 <= io_in_r_bypass_26_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_2_stall_2 <= io_in_r_bypass_26_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_3_data_2 <= io_in_r_bypass_26_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_3_load_store_2 <= io_in_r_bypass_26_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_3_df_is_ws_2 <= io_in_r_bypass_26_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_3_stall_2 <= io_in_r_bypass_26_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_0_data_2 <= io_in_r_bypass_27_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_0_load_store_2 <= io_in_r_bypass_27_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_0_df_is_ws_2 <= io_in_r_bypass_27_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_0_stall_2 <= io_in_r_bypass_27_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_1_data_2 <= io_in_r_bypass_27_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_1_load_store_2 <= io_in_r_bypass_27_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_1_df_is_ws_2 <= io_in_r_bypass_27_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_1_stall_2 <= io_in_r_bypass_27_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_2_data_2 <= io_in_r_bypass_27_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_2_load_store_2 <= io_in_r_bypass_27_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_2_df_is_ws_2 <= io_in_r_bypass_27_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_2_stall_2 <= io_in_r_bypass_27_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_3_data_2 <= io_in_r_bypass_27_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_3_load_store_2 <= io_in_r_bypass_27_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_3_df_is_ws_2 <= io_in_r_bypass_27_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_3_stall_2 <= io_in_r_bypass_27_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_0_data_2 <= io_in_r_bypass_28_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_0_load_store_2 <= io_in_r_bypass_28_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_0_df_is_ws_2 <= io_in_r_bypass_28_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_0_stall_2 <= io_in_r_bypass_28_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_1_data_2 <= io_in_r_bypass_28_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_1_load_store_2 <= io_in_r_bypass_28_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_1_df_is_ws_2 <= io_in_r_bypass_28_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_1_stall_2 <= io_in_r_bypass_28_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_2_data_2 <= io_in_r_bypass_28_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_2_load_store_2 <= io_in_r_bypass_28_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_2_df_is_ws_2 <= io_in_r_bypass_28_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_2_stall_2 <= io_in_r_bypass_28_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_3_data_2 <= io_in_r_bypass_28_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_3_load_store_2 <= io_in_r_bypass_28_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_3_df_is_ws_2 <= io_in_r_bypass_28_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_3_stall_2 <= io_in_r_bypass_28_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_0_data_2 <= io_in_r_bypass_29_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_0_load_store_2 <= io_in_r_bypass_29_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_0_df_is_ws_2 <= io_in_r_bypass_29_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_0_stall_2 <= io_in_r_bypass_29_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_1_data_2 <= io_in_r_bypass_29_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_1_load_store_2 <= io_in_r_bypass_29_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_1_df_is_ws_2 <= io_in_r_bypass_29_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_1_stall_2 <= io_in_r_bypass_29_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_2_data_2 <= io_in_r_bypass_29_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_2_load_store_2 <= io_in_r_bypass_29_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_2_df_is_ws_2 <= io_in_r_bypass_29_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_2_stall_2 <= io_in_r_bypass_29_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_3_data_2 <= io_in_r_bypass_29_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_3_load_store_2 <= io_in_r_bypass_29_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_3_df_is_ws_2 <= io_in_r_bypass_29_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_3_stall_2 <= io_in_r_bypass_29_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_0_data_2 <= io_in_r_bypass_30_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_0_load_store_2 <= io_in_r_bypass_30_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_0_df_is_ws_2 <= io_in_r_bypass_30_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_0_stall_2 <= io_in_r_bypass_30_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_1_data_2 <= io_in_r_bypass_30_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_1_load_store_2 <= io_in_r_bypass_30_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_1_df_is_ws_2 <= io_in_r_bypass_30_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_1_stall_2 <= io_in_r_bypass_30_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_2_data_2 <= io_in_r_bypass_30_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_2_load_store_2 <= io_in_r_bypass_30_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_2_df_is_ws_2 <= io_in_r_bypass_30_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_2_stall_2 <= io_in_r_bypass_30_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_3_data_2 <= io_in_r_bypass_30_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_3_load_store_2 <= io_in_r_bypass_30_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_3_df_is_ws_2 <= io_in_r_bypass_30_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_3_stall_2 <= io_in_r_bypass_30_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_0_data_2 <= io_in_r_bypass_31_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_0_load_store_2 <= io_in_r_bypass_31_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_0_df_is_ws_2 <= io_in_r_bypass_31_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_0_stall_2 <= io_in_r_bypass_31_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_1_data_2 <= io_in_r_bypass_31_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_1_load_store_2 <= io_in_r_bypass_31_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_1_df_is_ws_2 <= io_in_r_bypass_31_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_1_stall_2 <= io_in_r_bypass_31_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_2_data_2 <= io_in_r_bypass_31_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_2_load_store_2 <= io_in_r_bypass_31_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_2_df_is_ws_2 <= io_in_r_bypass_31_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_2_stall_2 <= io_in_r_bypass_31_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_3_data_2 <= io_in_r_bypass_31_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_3_load_store_2 <= io_in_r_bypass_31_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_3_df_is_ws_2 <= io_in_r_bypass_31_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_3_stall_2 <= io_in_r_bypass_31_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_0_data_3 <= io_in_r_bypass_0_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_0_load_store_3 <= io_in_r_bypass_0_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_0_df_is_ws_3 <= io_in_r_bypass_0_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_0_stall_3 <= io_in_r_bypass_0_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_1_data_3 <= io_in_r_bypass_0_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_1_load_store_3 <= io_in_r_bypass_0_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_1_df_is_ws_3 <= io_in_r_bypass_0_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_1_stall_3 <= io_in_r_bypass_0_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_2_data_3 <= io_in_r_bypass_0_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_2_load_store_3 <= io_in_r_bypass_0_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_2_df_is_ws_3 <= io_in_r_bypass_0_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_2_stall_3 <= io_in_r_bypass_0_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_3_data_3 <= io_in_r_bypass_0_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_3_load_store_3 <= io_in_r_bypass_0_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_3_df_is_ws_3 <= io_in_r_bypass_0_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_3_stall_3 <= io_in_r_bypass_0_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_0_data_3 <= io_in_r_bypass_1_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_0_load_store_3 <= io_in_r_bypass_1_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_0_df_is_ws_3 <= io_in_r_bypass_1_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_0_stall_3 <= io_in_r_bypass_1_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_1_data_3 <= io_in_r_bypass_1_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_1_load_store_3 <= io_in_r_bypass_1_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_1_df_is_ws_3 <= io_in_r_bypass_1_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_1_stall_3 <= io_in_r_bypass_1_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_2_data_3 <= io_in_r_bypass_1_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_2_load_store_3 <= io_in_r_bypass_1_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_2_df_is_ws_3 <= io_in_r_bypass_1_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_2_stall_3 <= io_in_r_bypass_1_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_3_data_3 <= io_in_r_bypass_1_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_3_load_store_3 <= io_in_r_bypass_1_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_3_df_is_ws_3 <= io_in_r_bypass_1_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_3_stall_3 <= io_in_r_bypass_1_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_0_data_3 <= io_in_r_bypass_2_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_0_load_store_3 <= io_in_r_bypass_2_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_0_df_is_ws_3 <= io_in_r_bypass_2_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_0_stall_3 <= io_in_r_bypass_2_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_1_data_3 <= io_in_r_bypass_2_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_1_load_store_3 <= io_in_r_bypass_2_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_1_df_is_ws_3 <= io_in_r_bypass_2_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_1_stall_3 <= io_in_r_bypass_2_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_2_data_3 <= io_in_r_bypass_2_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_2_load_store_3 <= io_in_r_bypass_2_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_2_df_is_ws_3 <= io_in_r_bypass_2_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_2_stall_3 <= io_in_r_bypass_2_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_3_data_3 <= io_in_r_bypass_2_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_3_load_store_3 <= io_in_r_bypass_2_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_3_df_is_ws_3 <= io_in_r_bypass_2_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_3_stall_3 <= io_in_r_bypass_2_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_0_data_3 <= io_in_r_bypass_3_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_0_load_store_3 <= io_in_r_bypass_3_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_0_df_is_ws_3 <= io_in_r_bypass_3_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_0_stall_3 <= io_in_r_bypass_3_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_1_data_3 <= io_in_r_bypass_3_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_1_load_store_3 <= io_in_r_bypass_3_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_1_df_is_ws_3 <= io_in_r_bypass_3_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_1_stall_3 <= io_in_r_bypass_3_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_2_data_3 <= io_in_r_bypass_3_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_2_load_store_3 <= io_in_r_bypass_3_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_2_df_is_ws_3 <= io_in_r_bypass_3_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_2_stall_3 <= io_in_r_bypass_3_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_3_data_3 <= io_in_r_bypass_3_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_3_load_store_3 <= io_in_r_bypass_3_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_3_df_is_ws_3 <= io_in_r_bypass_3_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_3_stall_3 <= io_in_r_bypass_3_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_0_data_3 <= io_in_r_bypass_4_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_0_load_store_3 <= io_in_r_bypass_4_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_0_df_is_ws_3 <= io_in_r_bypass_4_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_0_stall_3 <= io_in_r_bypass_4_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_1_data_3 <= io_in_r_bypass_4_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_1_load_store_3 <= io_in_r_bypass_4_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_1_df_is_ws_3 <= io_in_r_bypass_4_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_1_stall_3 <= io_in_r_bypass_4_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_2_data_3 <= io_in_r_bypass_4_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_2_load_store_3 <= io_in_r_bypass_4_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_2_df_is_ws_3 <= io_in_r_bypass_4_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_2_stall_3 <= io_in_r_bypass_4_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_3_data_3 <= io_in_r_bypass_4_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_3_load_store_3 <= io_in_r_bypass_4_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_3_df_is_ws_3 <= io_in_r_bypass_4_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_3_stall_3 <= io_in_r_bypass_4_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_0_data_3 <= io_in_r_bypass_5_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_0_load_store_3 <= io_in_r_bypass_5_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_0_df_is_ws_3 <= io_in_r_bypass_5_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_0_stall_3 <= io_in_r_bypass_5_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_1_data_3 <= io_in_r_bypass_5_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_1_load_store_3 <= io_in_r_bypass_5_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_1_df_is_ws_3 <= io_in_r_bypass_5_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_1_stall_3 <= io_in_r_bypass_5_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_2_data_3 <= io_in_r_bypass_5_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_2_load_store_3 <= io_in_r_bypass_5_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_2_df_is_ws_3 <= io_in_r_bypass_5_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_2_stall_3 <= io_in_r_bypass_5_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_3_data_3 <= io_in_r_bypass_5_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_3_load_store_3 <= io_in_r_bypass_5_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_3_df_is_ws_3 <= io_in_r_bypass_5_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_3_stall_3 <= io_in_r_bypass_5_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_0_data_3 <= io_in_r_bypass_6_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_0_load_store_3 <= io_in_r_bypass_6_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_0_df_is_ws_3 <= io_in_r_bypass_6_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_0_stall_3 <= io_in_r_bypass_6_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_1_data_3 <= io_in_r_bypass_6_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_1_load_store_3 <= io_in_r_bypass_6_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_1_df_is_ws_3 <= io_in_r_bypass_6_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_1_stall_3 <= io_in_r_bypass_6_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_2_data_3 <= io_in_r_bypass_6_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_2_load_store_3 <= io_in_r_bypass_6_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_2_df_is_ws_3 <= io_in_r_bypass_6_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_2_stall_3 <= io_in_r_bypass_6_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_3_data_3 <= io_in_r_bypass_6_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_3_load_store_3 <= io_in_r_bypass_6_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_3_df_is_ws_3 <= io_in_r_bypass_6_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_3_stall_3 <= io_in_r_bypass_6_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_0_data_3 <= io_in_r_bypass_7_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_0_load_store_3 <= io_in_r_bypass_7_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_0_df_is_ws_3 <= io_in_r_bypass_7_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_0_stall_3 <= io_in_r_bypass_7_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_1_data_3 <= io_in_r_bypass_7_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_1_load_store_3 <= io_in_r_bypass_7_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_1_df_is_ws_3 <= io_in_r_bypass_7_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_1_stall_3 <= io_in_r_bypass_7_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_2_data_3 <= io_in_r_bypass_7_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_2_load_store_3 <= io_in_r_bypass_7_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_2_df_is_ws_3 <= io_in_r_bypass_7_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_2_stall_3 <= io_in_r_bypass_7_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_3_data_3 <= io_in_r_bypass_7_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_3_load_store_3 <= io_in_r_bypass_7_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_3_df_is_ws_3 <= io_in_r_bypass_7_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_3_stall_3 <= io_in_r_bypass_7_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_0_data_3 <= io_in_r_bypass_8_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_0_load_store_3 <= io_in_r_bypass_8_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_0_df_is_ws_3 <= io_in_r_bypass_8_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_0_stall_3 <= io_in_r_bypass_8_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_1_data_3 <= io_in_r_bypass_8_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_1_load_store_3 <= io_in_r_bypass_8_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_1_df_is_ws_3 <= io_in_r_bypass_8_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_1_stall_3 <= io_in_r_bypass_8_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_2_data_3 <= io_in_r_bypass_8_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_2_load_store_3 <= io_in_r_bypass_8_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_2_df_is_ws_3 <= io_in_r_bypass_8_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_2_stall_3 <= io_in_r_bypass_8_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_3_data_3 <= io_in_r_bypass_8_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_3_load_store_3 <= io_in_r_bypass_8_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_3_df_is_ws_3 <= io_in_r_bypass_8_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_3_stall_3 <= io_in_r_bypass_8_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_0_data_3 <= io_in_r_bypass_9_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_0_load_store_3 <= io_in_r_bypass_9_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_0_df_is_ws_3 <= io_in_r_bypass_9_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_0_stall_3 <= io_in_r_bypass_9_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_1_data_3 <= io_in_r_bypass_9_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_1_load_store_3 <= io_in_r_bypass_9_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_1_df_is_ws_3 <= io_in_r_bypass_9_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_1_stall_3 <= io_in_r_bypass_9_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_2_data_3 <= io_in_r_bypass_9_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_2_load_store_3 <= io_in_r_bypass_9_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_2_df_is_ws_3 <= io_in_r_bypass_9_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_2_stall_3 <= io_in_r_bypass_9_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_3_data_3 <= io_in_r_bypass_9_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_3_load_store_3 <= io_in_r_bypass_9_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_3_df_is_ws_3 <= io_in_r_bypass_9_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_3_stall_3 <= io_in_r_bypass_9_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_0_data_3 <= io_in_r_bypass_10_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_0_load_store_3 <= io_in_r_bypass_10_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_0_df_is_ws_3 <= io_in_r_bypass_10_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_0_stall_3 <= io_in_r_bypass_10_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_1_data_3 <= io_in_r_bypass_10_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_1_load_store_3 <= io_in_r_bypass_10_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_1_df_is_ws_3 <= io_in_r_bypass_10_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_1_stall_3 <= io_in_r_bypass_10_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_2_data_3 <= io_in_r_bypass_10_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_2_load_store_3 <= io_in_r_bypass_10_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_2_df_is_ws_3 <= io_in_r_bypass_10_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_2_stall_3 <= io_in_r_bypass_10_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_3_data_3 <= io_in_r_bypass_10_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_3_load_store_3 <= io_in_r_bypass_10_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_3_df_is_ws_3 <= io_in_r_bypass_10_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_3_stall_3 <= io_in_r_bypass_10_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_0_data_3 <= io_in_r_bypass_11_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_0_load_store_3 <= io_in_r_bypass_11_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_0_df_is_ws_3 <= io_in_r_bypass_11_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_0_stall_3 <= io_in_r_bypass_11_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_1_data_3 <= io_in_r_bypass_11_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_1_load_store_3 <= io_in_r_bypass_11_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_1_df_is_ws_3 <= io_in_r_bypass_11_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_1_stall_3 <= io_in_r_bypass_11_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_2_data_3 <= io_in_r_bypass_11_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_2_load_store_3 <= io_in_r_bypass_11_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_2_df_is_ws_3 <= io_in_r_bypass_11_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_2_stall_3 <= io_in_r_bypass_11_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_3_data_3 <= io_in_r_bypass_11_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_3_load_store_3 <= io_in_r_bypass_11_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_3_df_is_ws_3 <= io_in_r_bypass_11_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_3_stall_3 <= io_in_r_bypass_11_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_0_data_3 <= io_in_r_bypass_12_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_0_load_store_3 <= io_in_r_bypass_12_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_0_df_is_ws_3 <= io_in_r_bypass_12_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_0_stall_3 <= io_in_r_bypass_12_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_1_data_3 <= io_in_r_bypass_12_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_1_load_store_3 <= io_in_r_bypass_12_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_1_df_is_ws_3 <= io_in_r_bypass_12_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_1_stall_3 <= io_in_r_bypass_12_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_2_data_3 <= io_in_r_bypass_12_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_2_load_store_3 <= io_in_r_bypass_12_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_2_df_is_ws_3 <= io_in_r_bypass_12_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_2_stall_3 <= io_in_r_bypass_12_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_3_data_3 <= io_in_r_bypass_12_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_3_load_store_3 <= io_in_r_bypass_12_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_3_df_is_ws_3 <= io_in_r_bypass_12_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_3_stall_3 <= io_in_r_bypass_12_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_0_data_3 <= io_in_r_bypass_13_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_0_load_store_3 <= io_in_r_bypass_13_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_0_df_is_ws_3 <= io_in_r_bypass_13_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_0_stall_3 <= io_in_r_bypass_13_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_1_data_3 <= io_in_r_bypass_13_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_1_load_store_3 <= io_in_r_bypass_13_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_1_df_is_ws_3 <= io_in_r_bypass_13_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_1_stall_3 <= io_in_r_bypass_13_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_2_data_3 <= io_in_r_bypass_13_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_2_load_store_3 <= io_in_r_bypass_13_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_2_df_is_ws_3 <= io_in_r_bypass_13_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_2_stall_3 <= io_in_r_bypass_13_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_3_data_3 <= io_in_r_bypass_13_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_3_load_store_3 <= io_in_r_bypass_13_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_3_df_is_ws_3 <= io_in_r_bypass_13_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_3_stall_3 <= io_in_r_bypass_13_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_0_data_3 <= io_in_r_bypass_14_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_0_load_store_3 <= io_in_r_bypass_14_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_0_df_is_ws_3 <= io_in_r_bypass_14_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_0_stall_3 <= io_in_r_bypass_14_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_1_data_3 <= io_in_r_bypass_14_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_1_load_store_3 <= io_in_r_bypass_14_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_1_df_is_ws_3 <= io_in_r_bypass_14_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_1_stall_3 <= io_in_r_bypass_14_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_2_data_3 <= io_in_r_bypass_14_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_2_load_store_3 <= io_in_r_bypass_14_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_2_df_is_ws_3 <= io_in_r_bypass_14_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_2_stall_3 <= io_in_r_bypass_14_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_3_data_3 <= io_in_r_bypass_14_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_3_load_store_3 <= io_in_r_bypass_14_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_3_df_is_ws_3 <= io_in_r_bypass_14_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_3_stall_3 <= io_in_r_bypass_14_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_0_data_3 <= io_in_r_bypass_15_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_0_load_store_3 <= io_in_r_bypass_15_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_0_df_is_ws_3 <= io_in_r_bypass_15_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_0_stall_3 <= io_in_r_bypass_15_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_1_data_3 <= io_in_r_bypass_15_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_1_load_store_3 <= io_in_r_bypass_15_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_1_df_is_ws_3 <= io_in_r_bypass_15_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_1_stall_3 <= io_in_r_bypass_15_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_2_data_3 <= io_in_r_bypass_15_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_2_load_store_3 <= io_in_r_bypass_15_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_2_df_is_ws_3 <= io_in_r_bypass_15_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_2_stall_3 <= io_in_r_bypass_15_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_3_data_3 <= io_in_r_bypass_15_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_3_load_store_3 <= io_in_r_bypass_15_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_3_df_is_ws_3 <= io_in_r_bypass_15_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_3_stall_3 <= io_in_r_bypass_15_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_0_data_3 <= io_in_r_bypass_16_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_0_load_store_3 <= io_in_r_bypass_16_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_0_df_is_ws_3 <= io_in_r_bypass_16_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_0_stall_3 <= io_in_r_bypass_16_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_1_data_3 <= io_in_r_bypass_16_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_1_load_store_3 <= io_in_r_bypass_16_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_1_df_is_ws_3 <= io_in_r_bypass_16_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_1_stall_3 <= io_in_r_bypass_16_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_2_data_3 <= io_in_r_bypass_16_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_2_load_store_3 <= io_in_r_bypass_16_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_2_df_is_ws_3 <= io_in_r_bypass_16_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_2_stall_3 <= io_in_r_bypass_16_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_3_data_3 <= io_in_r_bypass_16_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_3_load_store_3 <= io_in_r_bypass_16_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_3_df_is_ws_3 <= io_in_r_bypass_16_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_3_stall_3 <= io_in_r_bypass_16_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_0_data_3 <= io_in_r_bypass_17_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_0_load_store_3 <= io_in_r_bypass_17_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_0_df_is_ws_3 <= io_in_r_bypass_17_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_0_stall_3 <= io_in_r_bypass_17_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_1_data_3 <= io_in_r_bypass_17_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_1_load_store_3 <= io_in_r_bypass_17_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_1_df_is_ws_3 <= io_in_r_bypass_17_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_1_stall_3 <= io_in_r_bypass_17_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_2_data_3 <= io_in_r_bypass_17_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_2_load_store_3 <= io_in_r_bypass_17_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_2_df_is_ws_3 <= io_in_r_bypass_17_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_2_stall_3 <= io_in_r_bypass_17_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_3_data_3 <= io_in_r_bypass_17_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_3_load_store_3 <= io_in_r_bypass_17_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_3_df_is_ws_3 <= io_in_r_bypass_17_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_3_stall_3 <= io_in_r_bypass_17_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_0_data_3 <= io_in_r_bypass_18_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_0_load_store_3 <= io_in_r_bypass_18_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_0_df_is_ws_3 <= io_in_r_bypass_18_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_0_stall_3 <= io_in_r_bypass_18_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_1_data_3 <= io_in_r_bypass_18_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_1_load_store_3 <= io_in_r_bypass_18_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_1_df_is_ws_3 <= io_in_r_bypass_18_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_1_stall_3 <= io_in_r_bypass_18_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_2_data_3 <= io_in_r_bypass_18_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_2_load_store_3 <= io_in_r_bypass_18_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_2_df_is_ws_3 <= io_in_r_bypass_18_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_2_stall_3 <= io_in_r_bypass_18_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_3_data_3 <= io_in_r_bypass_18_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_3_load_store_3 <= io_in_r_bypass_18_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_3_df_is_ws_3 <= io_in_r_bypass_18_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_3_stall_3 <= io_in_r_bypass_18_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_0_data_3 <= io_in_r_bypass_19_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_0_load_store_3 <= io_in_r_bypass_19_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_0_df_is_ws_3 <= io_in_r_bypass_19_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_0_stall_3 <= io_in_r_bypass_19_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_1_data_3 <= io_in_r_bypass_19_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_1_load_store_3 <= io_in_r_bypass_19_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_1_df_is_ws_3 <= io_in_r_bypass_19_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_1_stall_3 <= io_in_r_bypass_19_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_2_data_3 <= io_in_r_bypass_19_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_2_load_store_3 <= io_in_r_bypass_19_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_2_df_is_ws_3 <= io_in_r_bypass_19_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_2_stall_3 <= io_in_r_bypass_19_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_3_data_3 <= io_in_r_bypass_19_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_3_load_store_3 <= io_in_r_bypass_19_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_3_df_is_ws_3 <= io_in_r_bypass_19_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_3_stall_3 <= io_in_r_bypass_19_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_0_data_3 <= io_in_r_bypass_20_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_0_load_store_3 <= io_in_r_bypass_20_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_0_df_is_ws_3 <= io_in_r_bypass_20_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_0_stall_3 <= io_in_r_bypass_20_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_1_data_3 <= io_in_r_bypass_20_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_1_load_store_3 <= io_in_r_bypass_20_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_1_df_is_ws_3 <= io_in_r_bypass_20_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_1_stall_3 <= io_in_r_bypass_20_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_2_data_3 <= io_in_r_bypass_20_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_2_load_store_3 <= io_in_r_bypass_20_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_2_df_is_ws_3 <= io_in_r_bypass_20_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_2_stall_3 <= io_in_r_bypass_20_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_3_data_3 <= io_in_r_bypass_20_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_3_load_store_3 <= io_in_r_bypass_20_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_3_df_is_ws_3 <= io_in_r_bypass_20_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_3_stall_3 <= io_in_r_bypass_20_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_0_data_3 <= io_in_r_bypass_21_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_0_load_store_3 <= io_in_r_bypass_21_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_0_df_is_ws_3 <= io_in_r_bypass_21_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_0_stall_3 <= io_in_r_bypass_21_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_1_data_3 <= io_in_r_bypass_21_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_1_load_store_3 <= io_in_r_bypass_21_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_1_df_is_ws_3 <= io_in_r_bypass_21_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_1_stall_3 <= io_in_r_bypass_21_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_2_data_3 <= io_in_r_bypass_21_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_2_load_store_3 <= io_in_r_bypass_21_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_2_df_is_ws_3 <= io_in_r_bypass_21_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_2_stall_3 <= io_in_r_bypass_21_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_3_data_3 <= io_in_r_bypass_21_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_3_load_store_3 <= io_in_r_bypass_21_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_3_df_is_ws_3 <= io_in_r_bypass_21_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_3_stall_3 <= io_in_r_bypass_21_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_0_data_3 <= io_in_r_bypass_22_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_0_load_store_3 <= io_in_r_bypass_22_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_0_df_is_ws_3 <= io_in_r_bypass_22_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_0_stall_3 <= io_in_r_bypass_22_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_1_data_3 <= io_in_r_bypass_22_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_1_load_store_3 <= io_in_r_bypass_22_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_1_df_is_ws_3 <= io_in_r_bypass_22_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_1_stall_3 <= io_in_r_bypass_22_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_2_data_3 <= io_in_r_bypass_22_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_2_load_store_3 <= io_in_r_bypass_22_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_2_df_is_ws_3 <= io_in_r_bypass_22_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_2_stall_3 <= io_in_r_bypass_22_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_3_data_3 <= io_in_r_bypass_22_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_3_load_store_3 <= io_in_r_bypass_22_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_3_df_is_ws_3 <= io_in_r_bypass_22_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_3_stall_3 <= io_in_r_bypass_22_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_0_data_3 <= io_in_r_bypass_23_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_0_load_store_3 <= io_in_r_bypass_23_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_0_df_is_ws_3 <= io_in_r_bypass_23_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_0_stall_3 <= io_in_r_bypass_23_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_1_data_3 <= io_in_r_bypass_23_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_1_load_store_3 <= io_in_r_bypass_23_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_1_df_is_ws_3 <= io_in_r_bypass_23_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_1_stall_3 <= io_in_r_bypass_23_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_2_data_3 <= io_in_r_bypass_23_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_2_load_store_3 <= io_in_r_bypass_23_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_2_df_is_ws_3 <= io_in_r_bypass_23_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_2_stall_3 <= io_in_r_bypass_23_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_3_data_3 <= io_in_r_bypass_23_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_3_load_store_3 <= io_in_r_bypass_23_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_3_df_is_ws_3 <= io_in_r_bypass_23_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_3_stall_3 <= io_in_r_bypass_23_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_0_data_3 <= io_in_r_bypass_24_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_0_load_store_3 <= io_in_r_bypass_24_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_0_df_is_ws_3 <= io_in_r_bypass_24_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_0_stall_3 <= io_in_r_bypass_24_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_1_data_3 <= io_in_r_bypass_24_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_1_load_store_3 <= io_in_r_bypass_24_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_1_df_is_ws_3 <= io_in_r_bypass_24_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_1_stall_3 <= io_in_r_bypass_24_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_2_data_3 <= io_in_r_bypass_24_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_2_load_store_3 <= io_in_r_bypass_24_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_2_df_is_ws_3 <= io_in_r_bypass_24_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_2_stall_3 <= io_in_r_bypass_24_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_3_data_3 <= io_in_r_bypass_24_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_3_load_store_3 <= io_in_r_bypass_24_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_3_df_is_ws_3 <= io_in_r_bypass_24_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_3_stall_3 <= io_in_r_bypass_24_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_0_data_3 <= io_in_r_bypass_25_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_0_load_store_3 <= io_in_r_bypass_25_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_0_df_is_ws_3 <= io_in_r_bypass_25_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_0_stall_3 <= io_in_r_bypass_25_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_1_data_3 <= io_in_r_bypass_25_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_1_load_store_3 <= io_in_r_bypass_25_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_1_df_is_ws_3 <= io_in_r_bypass_25_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_1_stall_3 <= io_in_r_bypass_25_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_2_data_3 <= io_in_r_bypass_25_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_2_load_store_3 <= io_in_r_bypass_25_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_2_df_is_ws_3 <= io_in_r_bypass_25_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_2_stall_3 <= io_in_r_bypass_25_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_3_data_3 <= io_in_r_bypass_25_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_3_load_store_3 <= io_in_r_bypass_25_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_3_df_is_ws_3 <= io_in_r_bypass_25_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_3_stall_3 <= io_in_r_bypass_25_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_0_data_3 <= io_in_r_bypass_26_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_0_load_store_3 <= io_in_r_bypass_26_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_0_df_is_ws_3 <= io_in_r_bypass_26_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_0_stall_3 <= io_in_r_bypass_26_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_1_data_3 <= io_in_r_bypass_26_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_1_load_store_3 <= io_in_r_bypass_26_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_1_df_is_ws_3 <= io_in_r_bypass_26_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_1_stall_3 <= io_in_r_bypass_26_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_2_data_3 <= io_in_r_bypass_26_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_2_load_store_3 <= io_in_r_bypass_26_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_2_df_is_ws_3 <= io_in_r_bypass_26_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_2_stall_3 <= io_in_r_bypass_26_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_3_data_3 <= io_in_r_bypass_26_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_3_load_store_3 <= io_in_r_bypass_26_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_3_df_is_ws_3 <= io_in_r_bypass_26_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_3_stall_3 <= io_in_r_bypass_26_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_0_data_3 <= io_in_r_bypass_27_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_0_load_store_3 <= io_in_r_bypass_27_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_0_df_is_ws_3 <= io_in_r_bypass_27_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_0_stall_3 <= io_in_r_bypass_27_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_1_data_3 <= io_in_r_bypass_27_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_1_load_store_3 <= io_in_r_bypass_27_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_1_df_is_ws_3 <= io_in_r_bypass_27_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_1_stall_3 <= io_in_r_bypass_27_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_2_data_3 <= io_in_r_bypass_27_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_2_load_store_3 <= io_in_r_bypass_27_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_2_df_is_ws_3 <= io_in_r_bypass_27_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_2_stall_3 <= io_in_r_bypass_27_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_3_data_3 <= io_in_r_bypass_27_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_3_load_store_3 <= io_in_r_bypass_27_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_3_df_is_ws_3 <= io_in_r_bypass_27_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_3_stall_3 <= io_in_r_bypass_27_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_0_data_3 <= io_in_r_bypass_28_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_0_load_store_3 <= io_in_r_bypass_28_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_0_df_is_ws_3 <= io_in_r_bypass_28_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_0_stall_3 <= io_in_r_bypass_28_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_1_data_3 <= io_in_r_bypass_28_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_1_load_store_3 <= io_in_r_bypass_28_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_1_df_is_ws_3 <= io_in_r_bypass_28_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_1_stall_3 <= io_in_r_bypass_28_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_2_data_3 <= io_in_r_bypass_28_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_2_load_store_3 <= io_in_r_bypass_28_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_2_df_is_ws_3 <= io_in_r_bypass_28_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_2_stall_3 <= io_in_r_bypass_28_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_3_data_3 <= io_in_r_bypass_28_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_3_load_store_3 <= io_in_r_bypass_28_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_3_df_is_ws_3 <= io_in_r_bypass_28_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_3_stall_3 <= io_in_r_bypass_28_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_0_data_3 <= io_in_r_bypass_29_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_0_load_store_3 <= io_in_r_bypass_29_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_0_df_is_ws_3 <= io_in_r_bypass_29_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_0_stall_3 <= io_in_r_bypass_29_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_1_data_3 <= io_in_r_bypass_29_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_1_load_store_3 <= io_in_r_bypass_29_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_1_df_is_ws_3 <= io_in_r_bypass_29_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_1_stall_3 <= io_in_r_bypass_29_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_2_data_3 <= io_in_r_bypass_29_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_2_load_store_3 <= io_in_r_bypass_29_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_2_df_is_ws_3 <= io_in_r_bypass_29_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_2_stall_3 <= io_in_r_bypass_29_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_3_data_3 <= io_in_r_bypass_29_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_3_load_store_3 <= io_in_r_bypass_29_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_3_df_is_ws_3 <= io_in_r_bypass_29_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_3_stall_3 <= io_in_r_bypass_29_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_0_data_3 <= io_in_r_bypass_30_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_0_load_store_3 <= io_in_r_bypass_30_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_0_df_is_ws_3 <= io_in_r_bypass_30_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_0_stall_3 <= io_in_r_bypass_30_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_1_data_3 <= io_in_r_bypass_30_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_1_load_store_3 <= io_in_r_bypass_30_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_1_df_is_ws_3 <= io_in_r_bypass_30_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_1_stall_3 <= io_in_r_bypass_30_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_2_data_3 <= io_in_r_bypass_30_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_2_load_store_3 <= io_in_r_bypass_30_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_2_df_is_ws_3 <= io_in_r_bypass_30_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_2_stall_3 <= io_in_r_bypass_30_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_3_data_3 <= io_in_r_bypass_30_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_3_load_store_3 <= io_in_r_bypass_30_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_3_df_is_ws_3 <= io_in_r_bypass_30_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_3_stall_3 <= io_in_r_bypass_30_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_0_data_3 <= io_in_r_bypass_31_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_0_load_store_3 <= io_in_r_bypass_31_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_0_df_is_ws_3 <= io_in_r_bypass_31_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_0_stall_3 <= io_in_r_bypass_31_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_1_data_3 <= io_in_r_bypass_31_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_1_load_store_3 <= io_in_r_bypass_31_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_1_df_is_ws_3 <= io_in_r_bypass_31_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_1_stall_3 <= io_in_r_bypass_31_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_2_data_3 <= io_in_r_bypass_31_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_2_load_store_3 <= io_in_r_bypass_31_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_2_df_is_ws_3 <= io_in_r_bypass_31_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_2_stall_3 <= io_in_r_bypass_31_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_3_data_3 <= io_in_r_bypass_31_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_3_load_store_3 <= io_in_r_bypass_31_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_3_df_is_ws_3 <= io_in_r_bypass_31_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_3_stall_3 <= io_in_r_bypass_31_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_0_data_4 <= io_in_r_bypass_0_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_0_load_store_4 <= io_in_r_bypass_0_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_0_df_is_ws_4 <= io_in_r_bypass_0_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_0_stall_4 <= io_in_r_bypass_0_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_1_data_4 <= io_in_r_bypass_0_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_1_load_store_4 <= io_in_r_bypass_0_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_1_df_is_ws_4 <= io_in_r_bypass_0_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_1_stall_4 <= io_in_r_bypass_0_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_2_data_4 <= io_in_r_bypass_0_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_2_load_store_4 <= io_in_r_bypass_0_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_2_df_is_ws_4 <= io_in_r_bypass_0_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_2_stall_4 <= io_in_r_bypass_0_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_3_data_4 <= io_in_r_bypass_0_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_3_load_store_4 <= io_in_r_bypass_0_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_3_df_is_ws_4 <= io_in_r_bypass_0_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_3_stall_4 <= io_in_r_bypass_0_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_0_data_4 <= io_in_r_bypass_1_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_0_load_store_4 <= io_in_r_bypass_1_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_0_df_is_ws_4 <= io_in_r_bypass_1_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_0_stall_4 <= io_in_r_bypass_1_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_1_data_4 <= io_in_r_bypass_1_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_1_load_store_4 <= io_in_r_bypass_1_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_1_df_is_ws_4 <= io_in_r_bypass_1_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_1_stall_4 <= io_in_r_bypass_1_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_2_data_4 <= io_in_r_bypass_1_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_2_load_store_4 <= io_in_r_bypass_1_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_2_df_is_ws_4 <= io_in_r_bypass_1_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_2_stall_4 <= io_in_r_bypass_1_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_3_data_4 <= io_in_r_bypass_1_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_3_load_store_4 <= io_in_r_bypass_1_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_3_df_is_ws_4 <= io_in_r_bypass_1_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_3_stall_4 <= io_in_r_bypass_1_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_0_data_4 <= io_in_r_bypass_2_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_0_load_store_4 <= io_in_r_bypass_2_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_0_df_is_ws_4 <= io_in_r_bypass_2_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_0_stall_4 <= io_in_r_bypass_2_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_1_data_4 <= io_in_r_bypass_2_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_1_load_store_4 <= io_in_r_bypass_2_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_1_df_is_ws_4 <= io_in_r_bypass_2_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_1_stall_4 <= io_in_r_bypass_2_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_2_data_4 <= io_in_r_bypass_2_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_2_load_store_4 <= io_in_r_bypass_2_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_2_df_is_ws_4 <= io_in_r_bypass_2_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_2_stall_4 <= io_in_r_bypass_2_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_3_data_4 <= io_in_r_bypass_2_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_3_load_store_4 <= io_in_r_bypass_2_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_3_df_is_ws_4 <= io_in_r_bypass_2_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_3_stall_4 <= io_in_r_bypass_2_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_0_data_4 <= io_in_r_bypass_3_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_0_load_store_4 <= io_in_r_bypass_3_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_0_df_is_ws_4 <= io_in_r_bypass_3_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_0_stall_4 <= io_in_r_bypass_3_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_1_data_4 <= io_in_r_bypass_3_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_1_load_store_4 <= io_in_r_bypass_3_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_1_df_is_ws_4 <= io_in_r_bypass_3_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_1_stall_4 <= io_in_r_bypass_3_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_2_data_4 <= io_in_r_bypass_3_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_2_load_store_4 <= io_in_r_bypass_3_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_2_df_is_ws_4 <= io_in_r_bypass_3_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_2_stall_4 <= io_in_r_bypass_3_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_3_data_4 <= io_in_r_bypass_3_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_3_load_store_4 <= io_in_r_bypass_3_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_3_df_is_ws_4 <= io_in_r_bypass_3_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_3_stall_4 <= io_in_r_bypass_3_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_0_data_4 <= io_in_r_bypass_4_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_0_load_store_4 <= io_in_r_bypass_4_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_0_df_is_ws_4 <= io_in_r_bypass_4_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_0_stall_4 <= io_in_r_bypass_4_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_1_data_4 <= io_in_r_bypass_4_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_1_load_store_4 <= io_in_r_bypass_4_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_1_df_is_ws_4 <= io_in_r_bypass_4_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_1_stall_4 <= io_in_r_bypass_4_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_2_data_4 <= io_in_r_bypass_4_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_2_load_store_4 <= io_in_r_bypass_4_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_2_df_is_ws_4 <= io_in_r_bypass_4_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_2_stall_4 <= io_in_r_bypass_4_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_3_data_4 <= io_in_r_bypass_4_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_3_load_store_4 <= io_in_r_bypass_4_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_3_df_is_ws_4 <= io_in_r_bypass_4_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_3_stall_4 <= io_in_r_bypass_4_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_0_data_4 <= io_in_r_bypass_5_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_0_load_store_4 <= io_in_r_bypass_5_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_0_df_is_ws_4 <= io_in_r_bypass_5_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_0_stall_4 <= io_in_r_bypass_5_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_1_data_4 <= io_in_r_bypass_5_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_1_load_store_4 <= io_in_r_bypass_5_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_1_df_is_ws_4 <= io_in_r_bypass_5_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_1_stall_4 <= io_in_r_bypass_5_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_2_data_4 <= io_in_r_bypass_5_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_2_load_store_4 <= io_in_r_bypass_5_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_2_df_is_ws_4 <= io_in_r_bypass_5_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_2_stall_4 <= io_in_r_bypass_5_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_3_data_4 <= io_in_r_bypass_5_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_3_load_store_4 <= io_in_r_bypass_5_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_3_df_is_ws_4 <= io_in_r_bypass_5_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_3_stall_4 <= io_in_r_bypass_5_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_0_data_4 <= io_in_r_bypass_6_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_0_load_store_4 <= io_in_r_bypass_6_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_0_df_is_ws_4 <= io_in_r_bypass_6_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_0_stall_4 <= io_in_r_bypass_6_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_1_data_4 <= io_in_r_bypass_6_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_1_load_store_4 <= io_in_r_bypass_6_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_1_df_is_ws_4 <= io_in_r_bypass_6_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_1_stall_4 <= io_in_r_bypass_6_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_2_data_4 <= io_in_r_bypass_6_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_2_load_store_4 <= io_in_r_bypass_6_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_2_df_is_ws_4 <= io_in_r_bypass_6_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_2_stall_4 <= io_in_r_bypass_6_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_3_data_4 <= io_in_r_bypass_6_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_3_load_store_4 <= io_in_r_bypass_6_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_3_df_is_ws_4 <= io_in_r_bypass_6_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_3_stall_4 <= io_in_r_bypass_6_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_0_data_4 <= io_in_r_bypass_7_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_0_load_store_4 <= io_in_r_bypass_7_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_0_df_is_ws_4 <= io_in_r_bypass_7_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_0_stall_4 <= io_in_r_bypass_7_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_1_data_4 <= io_in_r_bypass_7_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_1_load_store_4 <= io_in_r_bypass_7_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_1_df_is_ws_4 <= io_in_r_bypass_7_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_1_stall_4 <= io_in_r_bypass_7_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_2_data_4 <= io_in_r_bypass_7_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_2_load_store_4 <= io_in_r_bypass_7_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_2_df_is_ws_4 <= io_in_r_bypass_7_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_2_stall_4 <= io_in_r_bypass_7_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_3_data_4 <= io_in_r_bypass_7_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_3_load_store_4 <= io_in_r_bypass_7_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_3_df_is_ws_4 <= io_in_r_bypass_7_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_3_stall_4 <= io_in_r_bypass_7_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_0_data_4 <= io_in_r_bypass_8_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_0_load_store_4 <= io_in_r_bypass_8_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_0_df_is_ws_4 <= io_in_r_bypass_8_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_0_stall_4 <= io_in_r_bypass_8_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_1_data_4 <= io_in_r_bypass_8_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_1_load_store_4 <= io_in_r_bypass_8_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_1_df_is_ws_4 <= io_in_r_bypass_8_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_1_stall_4 <= io_in_r_bypass_8_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_2_data_4 <= io_in_r_bypass_8_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_2_load_store_4 <= io_in_r_bypass_8_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_2_df_is_ws_4 <= io_in_r_bypass_8_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_2_stall_4 <= io_in_r_bypass_8_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_3_data_4 <= io_in_r_bypass_8_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_3_load_store_4 <= io_in_r_bypass_8_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_3_df_is_ws_4 <= io_in_r_bypass_8_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_3_stall_4 <= io_in_r_bypass_8_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_0_data_4 <= io_in_r_bypass_9_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_0_load_store_4 <= io_in_r_bypass_9_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_0_df_is_ws_4 <= io_in_r_bypass_9_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_0_stall_4 <= io_in_r_bypass_9_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_1_data_4 <= io_in_r_bypass_9_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_1_load_store_4 <= io_in_r_bypass_9_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_1_df_is_ws_4 <= io_in_r_bypass_9_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_1_stall_4 <= io_in_r_bypass_9_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_2_data_4 <= io_in_r_bypass_9_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_2_load_store_4 <= io_in_r_bypass_9_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_2_df_is_ws_4 <= io_in_r_bypass_9_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_2_stall_4 <= io_in_r_bypass_9_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_3_data_4 <= io_in_r_bypass_9_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_3_load_store_4 <= io_in_r_bypass_9_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_3_df_is_ws_4 <= io_in_r_bypass_9_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_3_stall_4 <= io_in_r_bypass_9_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_0_data_4 <= io_in_r_bypass_10_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_0_load_store_4 <= io_in_r_bypass_10_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_0_df_is_ws_4 <= io_in_r_bypass_10_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_0_stall_4 <= io_in_r_bypass_10_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_1_data_4 <= io_in_r_bypass_10_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_1_load_store_4 <= io_in_r_bypass_10_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_1_df_is_ws_4 <= io_in_r_bypass_10_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_1_stall_4 <= io_in_r_bypass_10_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_2_data_4 <= io_in_r_bypass_10_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_2_load_store_4 <= io_in_r_bypass_10_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_2_df_is_ws_4 <= io_in_r_bypass_10_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_2_stall_4 <= io_in_r_bypass_10_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_3_data_4 <= io_in_r_bypass_10_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_3_load_store_4 <= io_in_r_bypass_10_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_3_df_is_ws_4 <= io_in_r_bypass_10_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_3_stall_4 <= io_in_r_bypass_10_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_0_data_4 <= io_in_r_bypass_11_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_0_load_store_4 <= io_in_r_bypass_11_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_0_df_is_ws_4 <= io_in_r_bypass_11_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_0_stall_4 <= io_in_r_bypass_11_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_1_data_4 <= io_in_r_bypass_11_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_1_load_store_4 <= io_in_r_bypass_11_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_1_df_is_ws_4 <= io_in_r_bypass_11_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_1_stall_4 <= io_in_r_bypass_11_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_2_data_4 <= io_in_r_bypass_11_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_2_load_store_4 <= io_in_r_bypass_11_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_2_df_is_ws_4 <= io_in_r_bypass_11_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_2_stall_4 <= io_in_r_bypass_11_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_3_data_4 <= io_in_r_bypass_11_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_3_load_store_4 <= io_in_r_bypass_11_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_3_df_is_ws_4 <= io_in_r_bypass_11_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_3_stall_4 <= io_in_r_bypass_11_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_0_data_4 <= io_in_r_bypass_12_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_0_load_store_4 <= io_in_r_bypass_12_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_0_df_is_ws_4 <= io_in_r_bypass_12_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_0_stall_4 <= io_in_r_bypass_12_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_1_data_4 <= io_in_r_bypass_12_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_1_load_store_4 <= io_in_r_bypass_12_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_1_df_is_ws_4 <= io_in_r_bypass_12_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_1_stall_4 <= io_in_r_bypass_12_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_2_data_4 <= io_in_r_bypass_12_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_2_load_store_4 <= io_in_r_bypass_12_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_2_df_is_ws_4 <= io_in_r_bypass_12_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_2_stall_4 <= io_in_r_bypass_12_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_3_data_4 <= io_in_r_bypass_12_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_3_load_store_4 <= io_in_r_bypass_12_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_3_df_is_ws_4 <= io_in_r_bypass_12_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_3_stall_4 <= io_in_r_bypass_12_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_0_data_4 <= io_in_r_bypass_13_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_0_load_store_4 <= io_in_r_bypass_13_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_0_df_is_ws_4 <= io_in_r_bypass_13_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_0_stall_4 <= io_in_r_bypass_13_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_1_data_4 <= io_in_r_bypass_13_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_1_load_store_4 <= io_in_r_bypass_13_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_1_df_is_ws_4 <= io_in_r_bypass_13_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_1_stall_4 <= io_in_r_bypass_13_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_2_data_4 <= io_in_r_bypass_13_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_2_load_store_4 <= io_in_r_bypass_13_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_2_df_is_ws_4 <= io_in_r_bypass_13_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_2_stall_4 <= io_in_r_bypass_13_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_3_data_4 <= io_in_r_bypass_13_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_3_load_store_4 <= io_in_r_bypass_13_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_3_df_is_ws_4 <= io_in_r_bypass_13_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_3_stall_4 <= io_in_r_bypass_13_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_0_data_4 <= io_in_r_bypass_14_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_0_load_store_4 <= io_in_r_bypass_14_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_0_df_is_ws_4 <= io_in_r_bypass_14_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_0_stall_4 <= io_in_r_bypass_14_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_1_data_4 <= io_in_r_bypass_14_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_1_load_store_4 <= io_in_r_bypass_14_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_1_df_is_ws_4 <= io_in_r_bypass_14_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_1_stall_4 <= io_in_r_bypass_14_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_2_data_4 <= io_in_r_bypass_14_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_2_load_store_4 <= io_in_r_bypass_14_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_2_df_is_ws_4 <= io_in_r_bypass_14_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_2_stall_4 <= io_in_r_bypass_14_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_3_data_4 <= io_in_r_bypass_14_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_3_load_store_4 <= io_in_r_bypass_14_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_3_df_is_ws_4 <= io_in_r_bypass_14_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_3_stall_4 <= io_in_r_bypass_14_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_0_data_4 <= io_in_r_bypass_15_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_0_load_store_4 <= io_in_r_bypass_15_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_0_df_is_ws_4 <= io_in_r_bypass_15_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_0_stall_4 <= io_in_r_bypass_15_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_1_data_4 <= io_in_r_bypass_15_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_1_load_store_4 <= io_in_r_bypass_15_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_1_df_is_ws_4 <= io_in_r_bypass_15_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_1_stall_4 <= io_in_r_bypass_15_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_2_data_4 <= io_in_r_bypass_15_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_2_load_store_4 <= io_in_r_bypass_15_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_2_df_is_ws_4 <= io_in_r_bypass_15_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_2_stall_4 <= io_in_r_bypass_15_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_3_data_4 <= io_in_r_bypass_15_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_3_load_store_4 <= io_in_r_bypass_15_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_3_df_is_ws_4 <= io_in_r_bypass_15_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_3_stall_4 <= io_in_r_bypass_15_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_0_data_4 <= io_in_r_bypass_16_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_0_load_store_4 <= io_in_r_bypass_16_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_0_df_is_ws_4 <= io_in_r_bypass_16_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_0_stall_4 <= io_in_r_bypass_16_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_1_data_4 <= io_in_r_bypass_16_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_1_load_store_4 <= io_in_r_bypass_16_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_1_df_is_ws_4 <= io_in_r_bypass_16_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_1_stall_4 <= io_in_r_bypass_16_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_2_data_4 <= io_in_r_bypass_16_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_2_load_store_4 <= io_in_r_bypass_16_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_2_df_is_ws_4 <= io_in_r_bypass_16_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_2_stall_4 <= io_in_r_bypass_16_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_3_data_4 <= io_in_r_bypass_16_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_3_load_store_4 <= io_in_r_bypass_16_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_3_df_is_ws_4 <= io_in_r_bypass_16_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_3_stall_4 <= io_in_r_bypass_16_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_0_data_4 <= io_in_r_bypass_17_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_0_load_store_4 <= io_in_r_bypass_17_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_0_df_is_ws_4 <= io_in_r_bypass_17_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_0_stall_4 <= io_in_r_bypass_17_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_1_data_4 <= io_in_r_bypass_17_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_1_load_store_4 <= io_in_r_bypass_17_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_1_df_is_ws_4 <= io_in_r_bypass_17_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_1_stall_4 <= io_in_r_bypass_17_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_2_data_4 <= io_in_r_bypass_17_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_2_load_store_4 <= io_in_r_bypass_17_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_2_df_is_ws_4 <= io_in_r_bypass_17_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_2_stall_4 <= io_in_r_bypass_17_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_3_data_4 <= io_in_r_bypass_17_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_3_load_store_4 <= io_in_r_bypass_17_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_3_df_is_ws_4 <= io_in_r_bypass_17_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_3_stall_4 <= io_in_r_bypass_17_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_0_data_4 <= io_in_r_bypass_18_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_0_load_store_4 <= io_in_r_bypass_18_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_0_df_is_ws_4 <= io_in_r_bypass_18_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_0_stall_4 <= io_in_r_bypass_18_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_1_data_4 <= io_in_r_bypass_18_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_1_load_store_4 <= io_in_r_bypass_18_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_1_df_is_ws_4 <= io_in_r_bypass_18_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_1_stall_4 <= io_in_r_bypass_18_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_2_data_4 <= io_in_r_bypass_18_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_2_load_store_4 <= io_in_r_bypass_18_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_2_df_is_ws_4 <= io_in_r_bypass_18_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_2_stall_4 <= io_in_r_bypass_18_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_3_data_4 <= io_in_r_bypass_18_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_3_load_store_4 <= io_in_r_bypass_18_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_3_df_is_ws_4 <= io_in_r_bypass_18_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_3_stall_4 <= io_in_r_bypass_18_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_0_data_4 <= io_in_r_bypass_19_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_0_load_store_4 <= io_in_r_bypass_19_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_0_df_is_ws_4 <= io_in_r_bypass_19_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_0_stall_4 <= io_in_r_bypass_19_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_1_data_4 <= io_in_r_bypass_19_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_1_load_store_4 <= io_in_r_bypass_19_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_1_df_is_ws_4 <= io_in_r_bypass_19_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_1_stall_4 <= io_in_r_bypass_19_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_2_data_4 <= io_in_r_bypass_19_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_2_load_store_4 <= io_in_r_bypass_19_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_2_df_is_ws_4 <= io_in_r_bypass_19_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_2_stall_4 <= io_in_r_bypass_19_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_3_data_4 <= io_in_r_bypass_19_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_3_load_store_4 <= io_in_r_bypass_19_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_3_df_is_ws_4 <= io_in_r_bypass_19_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_3_stall_4 <= io_in_r_bypass_19_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_0_data_4 <= io_in_r_bypass_20_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_0_load_store_4 <= io_in_r_bypass_20_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_0_df_is_ws_4 <= io_in_r_bypass_20_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_0_stall_4 <= io_in_r_bypass_20_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_1_data_4 <= io_in_r_bypass_20_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_1_load_store_4 <= io_in_r_bypass_20_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_1_df_is_ws_4 <= io_in_r_bypass_20_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_1_stall_4 <= io_in_r_bypass_20_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_2_data_4 <= io_in_r_bypass_20_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_2_load_store_4 <= io_in_r_bypass_20_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_2_df_is_ws_4 <= io_in_r_bypass_20_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_2_stall_4 <= io_in_r_bypass_20_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_3_data_4 <= io_in_r_bypass_20_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_3_load_store_4 <= io_in_r_bypass_20_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_3_df_is_ws_4 <= io_in_r_bypass_20_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_3_stall_4 <= io_in_r_bypass_20_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_0_data_4 <= io_in_r_bypass_21_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_0_load_store_4 <= io_in_r_bypass_21_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_0_df_is_ws_4 <= io_in_r_bypass_21_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_0_stall_4 <= io_in_r_bypass_21_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_1_data_4 <= io_in_r_bypass_21_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_1_load_store_4 <= io_in_r_bypass_21_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_1_df_is_ws_4 <= io_in_r_bypass_21_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_1_stall_4 <= io_in_r_bypass_21_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_2_data_4 <= io_in_r_bypass_21_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_2_load_store_4 <= io_in_r_bypass_21_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_2_df_is_ws_4 <= io_in_r_bypass_21_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_2_stall_4 <= io_in_r_bypass_21_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_3_data_4 <= io_in_r_bypass_21_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_3_load_store_4 <= io_in_r_bypass_21_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_3_df_is_ws_4 <= io_in_r_bypass_21_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_3_stall_4 <= io_in_r_bypass_21_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_0_data_4 <= io_in_r_bypass_22_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_0_load_store_4 <= io_in_r_bypass_22_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_0_df_is_ws_4 <= io_in_r_bypass_22_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_0_stall_4 <= io_in_r_bypass_22_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_1_data_4 <= io_in_r_bypass_22_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_1_load_store_4 <= io_in_r_bypass_22_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_1_df_is_ws_4 <= io_in_r_bypass_22_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_1_stall_4 <= io_in_r_bypass_22_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_2_data_4 <= io_in_r_bypass_22_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_2_load_store_4 <= io_in_r_bypass_22_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_2_df_is_ws_4 <= io_in_r_bypass_22_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_2_stall_4 <= io_in_r_bypass_22_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_3_data_4 <= io_in_r_bypass_22_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_3_load_store_4 <= io_in_r_bypass_22_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_3_df_is_ws_4 <= io_in_r_bypass_22_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_3_stall_4 <= io_in_r_bypass_22_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_0_data_4 <= io_in_r_bypass_23_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_0_load_store_4 <= io_in_r_bypass_23_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_0_df_is_ws_4 <= io_in_r_bypass_23_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_0_stall_4 <= io_in_r_bypass_23_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_1_data_4 <= io_in_r_bypass_23_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_1_load_store_4 <= io_in_r_bypass_23_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_1_df_is_ws_4 <= io_in_r_bypass_23_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_1_stall_4 <= io_in_r_bypass_23_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_2_data_4 <= io_in_r_bypass_23_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_2_load_store_4 <= io_in_r_bypass_23_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_2_df_is_ws_4 <= io_in_r_bypass_23_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_2_stall_4 <= io_in_r_bypass_23_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_3_data_4 <= io_in_r_bypass_23_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_3_load_store_4 <= io_in_r_bypass_23_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_3_df_is_ws_4 <= io_in_r_bypass_23_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_3_stall_4 <= io_in_r_bypass_23_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_0_data_4 <= io_in_r_bypass_24_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_0_load_store_4 <= io_in_r_bypass_24_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_0_df_is_ws_4 <= io_in_r_bypass_24_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_0_stall_4 <= io_in_r_bypass_24_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_1_data_4 <= io_in_r_bypass_24_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_1_load_store_4 <= io_in_r_bypass_24_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_1_df_is_ws_4 <= io_in_r_bypass_24_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_1_stall_4 <= io_in_r_bypass_24_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_2_data_4 <= io_in_r_bypass_24_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_2_load_store_4 <= io_in_r_bypass_24_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_2_df_is_ws_4 <= io_in_r_bypass_24_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_2_stall_4 <= io_in_r_bypass_24_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_3_data_4 <= io_in_r_bypass_24_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_3_load_store_4 <= io_in_r_bypass_24_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_3_df_is_ws_4 <= io_in_r_bypass_24_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_3_stall_4 <= io_in_r_bypass_24_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_0_data_4 <= io_in_r_bypass_25_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_0_load_store_4 <= io_in_r_bypass_25_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_0_df_is_ws_4 <= io_in_r_bypass_25_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_0_stall_4 <= io_in_r_bypass_25_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_1_data_4 <= io_in_r_bypass_25_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_1_load_store_4 <= io_in_r_bypass_25_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_1_df_is_ws_4 <= io_in_r_bypass_25_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_1_stall_4 <= io_in_r_bypass_25_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_2_data_4 <= io_in_r_bypass_25_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_2_load_store_4 <= io_in_r_bypass_25_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_2_df_is_ws_4 <= io_in_r_bypass_25_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_2_stall_4 <= io_in_r_bypass_25_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_3_data_4 <= io_in_r_bypass_25_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_3_load_store_4 <= io_in_r_bypass_25_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_3_df_is_ws_4 <= io_in_r_bypass_25_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_3_stall_4 <= io_in_r_bypass_25_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_0_data_4 <= io_in_r_bypass_26_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_0_load_store_4 <= io_in_r_bypass_26_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_0_df_is_ws_4 <= io_in_r_bypass_26_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_0_stall_4 <= io_in_r_bypass_26_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_1_data_4 <= io_in_r_bypass_26_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_1_load_store_4 <= io_in_r_bypass_26_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_1_df_is_ws_4 <= io_in_r_bypass_26_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_1_stall_4 <= io_in_r_bypass_26_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_2_data_4 <= io_in_r_bypass_26_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_2_load_store_4 <= io_in_r_bypass_26_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_2_df_is_ws_4 <= io_in_r_bypass_26_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_2_stall_4 <= io_in_r_bypass_26_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_3_data_4 <= io_in_r_bypass_26_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_3_load_store_4 <= io_in_r_bypass_26_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_3_df_is_ws_4 <= io_in_r_bypass_26_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_3_stall_4 <= io_in_r_bypass_26_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_0_data_4 <= io_in_r_bypass_27_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_0_load_store_4 <= io_in_r_bypass_27_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_0_df_is_ws_4 <= io_in_r_bypass_27_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_0_stall_4 <= io_in_r_bypass_27_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_1_data_4 <= io_in_r_bypass_27_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_1_load_store_4 <= io_in_r_bypass_27_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_1_df_is_ws_4 <= io_in_r_bypass_27_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_1_stall_4 <= io_in_r_bypass_27_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_2_data_4 <= io_in_r_bypass_27_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_2_load_store_4 <= io_in_r_bypass_27_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_2_df_is_ws_4 <= io_in_r_bypass_27_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_2_stall_4 <= io_in_r_bypass_27_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_3_data_4 <= io_in_r_bypass_27_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_3_load_store_4 <= io_in_r_bypass_27_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_3_df_is_ws_4 <= io_in_r_bypass_27_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_3_stall_4 <= io_in_r_bypass_27_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_0_data_4 <= io_in_r_bypass_28_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_0_load_store_4 <= io_in_r_bypass_28_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_0_df_is_ws_4 <= io_in_r_bypass_28_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_0_stall_4 <= io_in_r_bypass_28_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_1_data_4 <= io_in_r_bypass_28_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_1_load_store_4 <= io_in_r_bypass_28_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_1_df_is_ws_4 <= io_in_r_bypass_28_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_1_stall_4 <= io_in_r_bypass_28_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_2_data_4 <= io_in_r_bypass_28_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_2_load_store_4 <= io_in_r_bypass_28_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_2_df_is_ws_4 <= io_in_r_bypass_28_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_2_stall_4 <= io_in_r_bypass_28_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_3_data_4 <= io_in_r_bypass_28_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_3_load_store_4 <= io_in_r_bypass_28_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_3_df_is_ws_4 <= io_in_r_bypass_28_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_3_stall_4 <= io_in_r_bypass_28_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_0_data_4 <= io_in_r_bypass_29_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_0_load_store_4 <= io_in_r_bypass_29_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_0_df_is_ws_4 <= io_in_r_bypass_29_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_0_stall_4 <= io_in_r_bypass_29_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_1_data_4 <= io_in_r_bypass_29_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_1_load_store_4 <= io_in_r_bypass_29_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_1_df_is_ws_4 <= io_in_r_bypass_29_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_1_stall_4 <= io_in_r_bypass_29_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_2_data_4 <= io_in_r_bypass_29_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_2_load_store_4 <= io_in_r_bypass_29_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_2_df_is_ws_4 <= io_in_r_bypass_29_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_2_stall_4 <= io_in_r_bypass_29_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_3_data_4 <= io_in_r_bypass_29_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_3_load_store_4 <= io_in_r_bypass_29_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_3_df_is_ws_4 <= io_in_r_bypass_29_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_3_stall_4 <= io_in_r_bypass_29_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_0_data_4 <= io_in_r_bypass_30_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_0_load_store_4 <= io_in_r_bypass_30_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_0_df_is_ws_4 <= io_in_r_bypass_30_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_0_stall_4 <= io_in_r_bypass_30_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_1_data_4 <= io_in_r_bypass_30_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_1_load_store_4 <= io_in_r_bypass_30_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_1_df_is_ws_4 <= io_in_r_bypass_30_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_1_stall_4 <= io_in_r_bypass_30_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_2_data_4 <= io_in_r_bypass_30_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_2_load_store_4 <= io_in_r_bypass_30_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_2_df_is_ws_4 <= io_in_r_bypass_30_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_2_stall_4 <= io_in_r_bypass_30_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_3_data_4 <= io_in_r_bypass_30_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_3_load_store_4 <= io_in_r_bypass_30_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_3_df_is_ws_4 <= io_in_r_bypass_30_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_3_stall_4 <= io_in_r_bypass_30_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_0_data_4 <= io_in_r_bypass_31_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_0_load_store_4 <= io_in_r_bypass_31_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_0_df_is_ws_4 <= io_in_r_bypass_31_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_0_stall_4 <= io_in_r_bypass_31_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_1_data_4 <= io_in_r_bypass_31_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_1_load_store_4 <= io_in_r_bypass_31_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_1_df_is_ws_4 <= io_in_r_bypass_31_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_1_stall_4 <= io_in_r_bypass_31_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_2_data_4 <= io_in_r_bypass_31_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_2_load_store_4 <= io_in_r_bypass_31_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_2_df_is_ws_4 <= io_in_r_bypass_31_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_2_stall_4 <= io_in_r_bypass_31_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_3_data_4 <= io_in_r_bypass_31_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_3_load_store_4 <= io_in_r_bypass_31_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_3_df_is_ws_4 <= io_in_r_bypass_31_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_3_stall_4 <= io_in_r_bypass_31_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_0_data_5 <= io_in_r_bypass_0_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_0_load_store_5 <= io_in_r_bypass_0_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_0_df_is_ws_5 <= io_in_r_bypass_0_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_0_stall_5 <= io_in_r_bypass_0_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_1_data_5 <= io_in_r_bypass_0_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_1_load_store_5 <= io_in_r_bypass_0_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_1_df_is_ws_5 <= io_in_r_bypass_0_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_1_stall_5 <= io_in_r_bypass_0_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_2_data_5 <= io_in_r_bypass_0_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_2_load_store_5 <= io_in_r_bypass_0_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_2_df_is_ws_5 <= io_in_r_bypass_0_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_2_stall_5 <= io_in_r_bypass_0_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_3_data_5 <= io_in_r_bypass_0_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_3_load_store_5 <= io_in_r_bypass_0_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_3_df_is_ws_5 <= io_in_r_bypass_0_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_3_stall_5 <= io_in_r_bypass_0_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_0_data_5 <= io_in_r_bypass_1_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_0_load_store_5 <= io_in_r_bypass_1_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_0_df_is_ws_5 <= io_in_r_bypass_1_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_0_stall_5 <= io_in_r_bypass_1_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_1_data_5 <= io_in_r_bypass_1_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_1_load_store_5 <= io_in_r_bypass_1_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_1_df_is_ws_5 <= io_in_r_bypass_1_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_1_stall_5 <= io_in_r_bypass_1_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_2_data_5 <= io_in_r_bypass_1_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_2_load_store_5 <= io_in_r_bypass_1_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_2_df_is_ws_5 <= io_in_r_bypass_1_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_2_stall_5 <= io_in_r_bypass_1_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_3_data_5 <= io_in_r_bypass_1_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_3_load_store_5 <= io_in_r_bypass_1_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_3_df_is_ws_5 <= io_in_r_bypass_1_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_3_stall_5 <= io_in_r_bypass_1_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_0_data_5 <= io_in_r_bypass_2_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_0_load_store_5 <= io_in_r_bypass_2_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_0_df_is_ws_5 <= io_in_r_bypass_2_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_0_stall_5 <= io_in_r_bypass_2_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_1_data_5 <= io_in_r_bypass_2_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_1_load_store_5 <= io_in_r_bypass_2_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_1_df_is_ws_5 <= io_in_r_bypass_2_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_1_stall_5 <= io_in_r_bypass_2_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_2_data_5 <= io_in_r_bypass_2_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_2_load_store_5 <= io_in_r_bypass_2_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_2_df_is_ws_5 <= io_in_r_bypass_2_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_2_stall_5 <= io_in_r_bypass_2_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_3_data_5 <= io_in_r_bypass_2_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_3_load_store_5 <= io_in_r_bypass_2_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_3_df_is_ws_5 <= io_in_r_bypass_2_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_3_stall_5 <= io_in_r_bypass_2_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_0_data_5 <= io_in_r_bypass_3_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_0_load_store_5 <= io_in_r_bypass_3_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_0_df_is_ws_5 <= io_in_r_bypass_3_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_0_stall_5 <= io_in_r_bypass_3_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_1_data_5 <= io_in_r_bypass_3_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_1_load_store_5 <= io_in_r_bypass_3_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_1_df_is_ws_5 <= io_in_r_bypass_3_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_1_stall_5 <= io_in_r_bypass_3_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_2_data_5 <= io_in_r_bypass_3_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_2_load_store_5 <= io_in_r_bypass_3_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_2_df_is_ws_5 <= io_in_r_bypass_3_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_2_stall_5 <= io_in_r_bypass_3_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_3_data_5 <= io_in_r_bypass_3_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_3_load_store_5 <= io_in_r_bypass_3_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_3_df_is_ws_5 <= io_in_r_bypass_3_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_3_stall_5 <= io_in_r_bypass_3_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_0_data_5 <= io_in_r_bypass_4_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_0_load_store_5 <= io_in_r_bypass_4_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_0_df_is_ws_5 <= io_in_r_bypass_4_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_0_stall_5 <= io_in_r_bypass_4_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_1_data_5 <= io_in_r_bypass_4_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_1_load_store_5 <= io_in_r_bypass_4_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_1_df_is_ws_5 <= io_in_r_bypass_4_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_1_stall_5 <= io_in_r_bypass_4_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_2_data_5 <= io_in_r_bypass_4_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_2_load_store_5 <= io_in_r_bypass_4_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_2_df_is_ws_5 <= io_in_r_bypass_4_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_2_stall_5 <= io_in_r_bypass_4_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_3_data_5 <= io_in_r_bypass_4_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_3_load_store_5 <= io_in_r_bypass_4_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_3_df_is_ws_5 <= io_in_r_bypass_4_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_3_stall_5 <= io_in_r_bypass_4_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_0_data_5 <= io_in_r_bypass_5_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_0_load_store_5 <= io_in_r_bypass_5_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_0_df_is_ws_5 <= io_in_r_bypass_5_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_0_stall_5 <= io_in_r_bypass_5_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_1_data_5 <= io_in_r_bypass_5_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_1_load_store_5 <= io_in_r_bypass_5_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_1_df_is_ws_5 <= io_in_r_bypass_5_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_1_stall_5 <= io_in_r_bypass_5_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_2_data_5 <= io_in_r_bypass_5_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_2_load_store_5 <= io_in_r_bypass_5_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_2_df_is_ws_5 <= io_in_r_bypass_5_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_2_stall_5 <= io_in_r_bypass_5_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_3_data_5 <= io_in_r_bypass_5_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_3_load_store_5 <= io_in_r_bypass_5_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_3_df_is_ws_5 <= io_in_r_bypass_5_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_3_stall_5 <= io_in_r_bypass_5_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_0_data_5 <= io_in_r_bypass_6_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_0_load_store_5 <= io_in_r_bypass_6_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_0_df_is_ws_5 <= io_in_r_bypass_6_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_0_stall_5 <= io_in_r_bypass_6_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_1_data_5 <= io_in_r_bypass_6_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_1_load_store_5 <= io_in_r_bypass_6_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_1_df_is_ws_5 <= io_in_r_bypass_6_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_1_stall_5 <= io_in_r_bypass_6_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_2_data_5 <= io_in_r_bypass_6_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_2_load_store_5 <= io_in_r_bypass_6_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_2_df_is_ws_5 <= io_in_r_bypass_6_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_2_stall_5 <= io_in_r_bypass_6_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_3_data_5 <= io_in_r_bypass_6_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_3_load_store_5 <= io_in_r_bypass_6_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_3_df_is_ws_5 <= io_in_r_bypass_6_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_3_stall_5 <= io_in_r_bypass_6_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_0_data_5 <= io_in_r_bypass_7_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_0_load_store_5 <= io_in_r_bypass_7_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_0_df_is_ws_5 <= io_in_r_bypass_7_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_0_stall_5 <= io_in_r_bypass_7_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_1_data_5 <= io_in_r_bypass_7_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_1_load_store_5 <= io_in_r_bypass_7_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_1_df_is_ws_5 <= io_in_r_bypass_7_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_1_stall_5 <= io_in_r_bypass_7_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_2_data_5 <= io_in_r_bypass_7_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_2_load_store_5 <= io_in_r_bypass_7_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_2_df_is_ws_5 <= io_in_r_bypass_7_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_2_stall_5 <= io_in_r_bypass_7_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_3_data_5 <= io_in_r_bypass_7_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_3_load_store_5 <= io_in_r_bypass_7_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_3_df_is_ws_5 <= io_in_r_bypass_7_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_3_stall_5 <= io_in_r_bypass_7_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_0_data_5 <= io_in_r_bypass_8_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_0_load_store_5 <= io_in_r_bypass_8_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_0_df_is_ws_5 <= io_in_r_bypass_8_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_0_stall_5 <= io_in_r_bypass_8_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_1_data_5 <= io_in_r_bypass_8_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_1_load_store_5 <= io_in_r_bypass_8_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_1_df_is_ws_5 <= io_in_r_bypass_8_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_1_stall_5 <= io_in_r_bypass_8_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_2_data_5 <= io_in_r_bypass_8_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_2_load_store_5 <= io_in_r_bypass_8_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_2_df_is_ws_5 <= io_in_r_bypass_8_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_2_stall_5 <= io_in_r_bypass_8_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_3_data_5 <= io_in_r_bypass_8_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_3_load_store_5 <= io_in_r_bypass_8_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_3_df_is_ws_5 <= io_in_r_bypass_8_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_3_stall_5 <= io_in_r_bypass_8_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_0_data_5 <= io_in_r_bypass_9_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_0_load_store_5 <= io_in_r_bypass_9_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_0_df_is_ws_5 <= io_in_r_bypass_9_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_0_stall_5 <= io_in_r_bypass_9_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_1_data_5 <= io_in_r_bypass_9_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_1_load_store_5 <= io_in_r_bypass_9_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_1_df_is_ws_5 <= io_in_r_bypass_9_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_1_stall_5 <= io_in_r_bypass_9_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_2_data_5 <= io_in_r_bypass_9_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_2_load_store_5 <= io_in_r_bypass_9_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_2_df_is_ws_5 <= io_in_r_bypass_9_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_2_stall_5 <= io_in_r_bypass_9_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_3_data_5 <= io_in_r_bypass_9_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_3_load_store_5 <= io_in_r_bypass_9_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_3_df_is_ws_5 <= io_in_r_bypass_9_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_3_stall_5 <= io_in_r_bypass_9_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_0_data_5 <= io_in_r_bypass_10_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_0_load_store_5 <= io_in_r_bypass_10_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_0_df_is_ws_5 <= io_in_r_bypass_10_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_0_stall_5 <= io_in_r_bypass_10_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_1_data_5 <= io_in_r_bypass_10_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_1_load_store_5 <= io_in_r_bypass_10_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_1_df_is_ws_5 <= io_in_r_bypass_10_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_1_stall_5 <= io_in_r_bypass_10_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_2_data_5 <= io_in_r_bypass_10_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_2_load_store_5 <= io_in_r_bypass_10_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_2_df_is_ws_5 <= io_in_r_bypass_10_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_2_stall_5 <= io_in_r_bypass_10_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_3_data_5 <= io_in_r_bypass_10_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_3_load_store_5 <= io_in_r_bypass_10_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_3_df_is_ws_5 <= io_in_r_bypass_10_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_3_stall_5 <= io_in_r_bypass_10_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_0_data_5 <= io_in_r_bypass_11_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_0_load_store_5 <= io_in_r_bypass_11_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_0_df_is_ws_5 <= io_in_r_bypass_11_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_0_stall_5 <= io_in_r_bypass_11_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_1_data_5 <= io_in_r_bypass_11_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_1_load_store_5 <= io_in_r_bypass_11_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_1_df_is_ws_5 <= io_in_r_bypass_11_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_1_stall_5 <= io_in_r_bypass_11_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_2_data_5 <= io_in_r_bypass_11_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_2_load_store_5 <= io_in_r_bypass_11_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_2_df_is_ws_5 <= io_in_r_bypass_11_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_2_stall_5 <= io_in_r_bypass_11_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_3_data_5 <= io_in_r_bypass_11_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_3_load_store_5 <= io_in_r_bypass_11_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_3_df_is_ws_5 <= io_in_r_bypass_11_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_3_stall_5 <= io_in_r_bypass_11_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_0_data_5 <= io_in_r_bypass_12_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_0_load_store_5 <= io_in_r_bypass_12_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_0_df_is_ws_5 <= io_in_r_bypass_12_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_0_stall_5 <= io_in_r_bypass_12_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_1_data_5 <= io_in_r_bypass_12_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_1_load_store_5 <= io_in_r_bypass_12_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_1_df_is_ws_5 <= io_in_r_bypass_12_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_1_stall_5 <= io_in_r_bypass_12_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_2_data_5 <= io_in_r_bypass_12_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_2_load_store_5 <= io_in_r_bypass_12_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_2_df_is_ws_5 <= io_in_r_bypass_12_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_2_stall_5 <= io_in_r_bypass_12_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_3_data_5 <= io_in_r_bypass_12_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_3_load_store_5 <= io_in_r_bypass_12_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_3_df_is_ws_5 <= io_in_r_bypass_12_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_3_stall_5 <= io_in_r_bypass_12_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_0_data_5 <= io_in_r_bypass_13_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_0_load_store_5 <= io_in_r_bypass_13_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_0_df_is_ws_5 <= io_in_r_bypass_13_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_0_stall_5 <= io_in_r_bypass_13_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_1_data_5 <= io_in_r_bypass_13_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_1_load_store_5 <= io_in_r_bypass_13_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_1_df_is_ws_5 <= io_in_r_bypass_13_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_1_stall_5 <= io_in_r_bypass_13_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_2_data_5 <= io_in_r_bypass_13_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_2_load_store_5 <= io_in_r_bypass_13_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_2_df_is_ws_5 <= io_in_r_bypass_13_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_2_stall_5 <= io_in_r_bypass_13_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_3_data_5 <= io_in_r_bypass_13_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_3_load_store_5 <= io_in_r_bypass_13_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_3_df_is_ws_5 <= io_in_r_bypass_13_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_3_stall_5 <= io_in_r_bypass_13_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_0_data_5 <= io_in_r_bypass_14_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_0_load_store_5 <= io_in_r_bypass_14_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_0_df_is_ws_5 <= io_in_r_bypass_14_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_0_stall_5 <= io_in_r_bypass_14_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_1_data_5 <= io_in_r_bypass_14_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_1_load_store_5 <= io_in_r_bypass_14_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_1_df_is_ws_5 <= io_in_r_bypass_14_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_1_stall_5 <= io_in_r_bypass_14_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_2_data_5 <= io_in_r_bypass_14_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_2_load_store_5 <= io_in_r_bypass_14_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_2_df_is_ws_5 <= io_in_r_bypass_14_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_2_stall_5 <= io_in_r_bypass_14_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_3_data_5 <= io_in_r_bypass_14_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_3_load_store_5 <= io_in_r_bypass_14_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_3_df_is_ws_5 <= io_in_r_bypass_14_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_3_stall_5 <= io_in_r_bypass_14_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_0_data_5 <= io_in_r_bypass_15_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_0_load_store_5 <= io_in_r_bypass_15_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_0_df_is_ws_5 <= io_in_r_bypass_15_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_0_stall_5 <= io_in_r_bypass_15_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_1_data_5 <= io_in_r_bypass_15_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_1_load_store_5 <= io_in_r_bypass_15_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_1_df_is_ws_5 <= io_in_r_bypass_15_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_1_stall_5 <= io_in_r_bypass_15_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_2_data_5 <= io_in_r_bypass_15_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_2_load_store_5 <= io_in_r_bypass_15_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_2_df_is_ws_5 <= io_in_r_bypass_15_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_2_stall_5 <= io_in_r_bypass_15_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_3_data_5 <= io_in_r_bypass_15_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_3_load_store_5 <= io_in_r_bypass_15_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_3_df_is_ws_5 <= io_in_r_bypass_15_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_3_stall_5 <= io_in_r_bypass_15_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_0_data_5 <= io_in_r_bypass_16_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_0_load_store_5 <= io_in_r_bypass_16_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_0_df_is_ws_5 <= io_in_r_bypass_16_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_0_stall_5 <= io_in_r_bypass_16_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_1_data_5 <= io_in_r_bypass_16_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_1_load_store_5 <= io_in_r_bypass_16_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_1_df_is_ws_5 <= io_in_r_bypass_16_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_1_stall_5 <= io_in_r_bypass_16_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_2_data_5 <= io_in_r_bypass_16_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_2_load_store_5 <= io_in_r_bypass_16_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_2_df_is_ws_5 <= io_in_r_bypass_16_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_2_stall_5 <= io_in_r_bypass_16_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_3_data_5 <= io_in_r_bypass_16_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_3_load_store_5 <= io_in_r_bypass_16_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_3_df_is_ws_5 <= io_in_r_bypass_16_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_3_stall_5 <= io_in_r_bypass_16_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_0_data_5 <= io_in_r_bypass_17_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_0_load_store_5 <= io_in_r_bypass_17_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_0_df_is_ws_5 <= io_in_r_bypass_17_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_0_stall_5 <= io_in_r_bypass_17_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_1_data_5 <= io_in_r_bypass_17_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_1_load_store_5 <= io_in_r_bypass_17_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_1_df_is_ws_5 <= io_in_r_bypass_17_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_1_stall_5 <= io_in_r_bypass_17_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_2_data_5 <= io_in_r_bypass_17_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_2_load_store_5 <= io_in_r_bypass_17_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_2_df_is_ws_5 <= io_in_r_bypass_17_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_2_stall_5 <= io_in_r_bypass_17_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_3_data_5 <= io_in_r_bypass_17_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_3_load_store_5 <= io_in_r_bypass_17_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_3_df_is_ws_5 <= io_in_r_bypass_17_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_3_stall_5 <= io_in_r_bypass_17_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_0_data_5 <= io_in_r_bypass_18_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_0_load_store_5 <= io_in_r_bypass_18_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_0_df_is_ws_5 <= io_in_r_bypass_18_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_0_stall_5 <= io_in_r_bypass_18_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_1_data_5 <= io_in_r_bypass_18_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_1_load_store_5 <= io_in_r_bypass_18_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_1_df_is_ws_5 <= io_in_r_bypass_18_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_1_stall_5 <= io_in_r_bypass_18_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_2_data_5 <= io_in_r_bypass_18_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_2_load_store_5 <= io_in_r_bypass_18_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_2_df_is_ws_5 <= io_in_r_bypass_18_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_2_stall_5 <= io_in_r_bypass_18_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_3_data_5 <= io_in_r_bypass_18_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_3_load_store_5 <= io_in_r_bypass_18_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_3_df_is_ws_5 <= io_in_r_bypass_18_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_3_stall_5 <= io_in_r_bypass_18_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_0_data_5 <= io_in_r_bypass_19_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_0_load_store_5 <= io_in_r_bypass_19_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_0_df_is_ws_5 <= io_in_r_bypass_19_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_0_stall_5 <= io_in_r_bypass_19_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_1_data_5 <= io_in_r_bypass_19_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_1_load_store_5 <= io_in_r_bypass_19_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_1_df_is_ws_5 <= io_in_r_bypass_19_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_1_stall_5 <= io_in_r_bypass_19_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_2_data_5 <= io_in_r_bypass_19_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_2_load_store_5 <= io_in_r_bypass_19_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_2_df_is_ws_5 <= io_in_r_bypass_19_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_2_stall_5 <= io_in_r_bypass_19_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_3_data_5 <= io_in_r_bypass_19_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_3_load_store_5 <= io_in_r_bypass_19_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_3_df_is_ws_5 <= io_in_r_bypass_19_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_3_stall_5 <= io_in_r_bypass_19_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_0_data_5 <= io_in_r_bypass_20_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_0_load_store_5 <= io_in_r_bypass_20_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_0_df_is_ws_5 <= io_in_r_bypass_20_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_0_stall_5 <= io_in_r_bypass_20_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_1_data_5 <= io_in_r_bypass_20_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_1_load_store_5 <= io_in_r_bypass_20_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_1_df_is_ws_5 <= io_in_r_bypass_20_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_1_stall_5 <= io_in_r_bypass_20_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_2_data_5 <= io_in_r_bypass_20_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_2_load_store_5 <= io_in_r_bypass_20_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_2_df_is_ws_5 <= io_in_r_bypass_20_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_2_stall_5 <= io_in_r_bypass_20_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_3_data_5 <= io_in_r_bypass_20_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_3_load_store_5 <= io_in_r_bypass_20_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_3_df_is_ws_5 <= io_in_r_bypass_20_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_3_stall_5 <= io_in_r_bypass_20_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_0_data_5 <= io_in_r_bypass_21_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_0_load_store_5 <= io_in_r_bypass_21_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_0_df_is_ws_5 <= io_in_r_bypass_21_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_0_stall_5 <= io_in_r_bypass_21_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_1_data_5 <= io_in_r_bypass_21_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_1_load_store_5 <= io_in_r_bypass_21_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_1_df_is_ws_5 <= io_in_r_bypass_21_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_1_stall_5 <= io_in_r_bypass_21_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_2_data_5 <= io_in_r_bypass_21_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_2_load_store_5 <= io_in_r_bypass_21_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_2_df_is_ws_5 <= io_in_r_bypass_21_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_2_stall_5 <= io_in_r_bypass_21_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_3_data_5 <= io_in_r_bypass_21_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_3_load_store_5 <= io_in_r_bypass_21_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_3_df_is_ws_5 <= io_in_r_bypass_21_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_3_stall_5 <= io_in_r_bypass_21_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_0_data_5 <= io_in_r_bypass_22_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_0_load_store_5 <= io_in_r_bypass_22_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_0_df_is_ws_5 <= io_in_r_bypass_22_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_0_stall_5 <= io_in_r_bypass_22_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_1_data_5 <= io_in_r_bypass_22_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_1_load_store_5 <= io_in_r_bypass_22_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_1_df_is_ws_5 <= io_in_r_bypass_22_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_1_stall_5 <= io_in_r_bypass_22_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_2_data_5 <= io_in_r_bypass_22_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_2_load_store_5 <= io_in_r_bypass_22_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_2_df_is_ws_5 <= io_in_r_bypass_22_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_2_stall_5 <= io_in_r_bypass_22_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_3_data_5 <= io_in_r_bypass_22_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_3_load_store_5 <= io_in_r_bypass_22_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_3_df_is_ws_5 <= io_in_r_bypass_22_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_3_stall_5 <= io_in_r_bypass_22_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_0_data_5 <= io_in_r_bypass_23_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_0_load_store_5 <= io_in_r_bypass_23_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_0_df_is_ws_5 <= io_in_r_bypass_23_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_0_stall_5 <= io_in_r_bypass_23_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_1_data_5 <= io_in_r_bypass_23_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_1_load_store_5 <= io_in_r_bypass_23_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_1_df_is_ws_5 <= io_in_r_bypass_23_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_1_stall_5 <= io_in_r_bypass_23_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_2_data_5 <= io_in_r_bypass_23_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_2_load_store_5 <= io_in_r_bypass_23_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_2_df_is_ws_5 <= io_in_r_bypass_23_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_2_stall_5 <= io_in_r_bypass_23_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_3_data_5 <= io_in_r_bypass_23_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_3_load_store_5 <= io_in_r_bypass_23_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_3_df_is_ws_5 <= io_in_r_bypass_23_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_3_stall_5 <= io_in_r_bypass_23_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_0_data_5 <= io_in_r_bypass_24_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_0_load_store_5 <= io_in_r_bypass_24_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_0_df_is_ws_5 <= io_in_r_bypass_24_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_0_stall_5 <= io_in_r_bypass_24_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_1_data_5 <= io_in_r_bypass_24_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_1_load_store_5 <= io_in_r_bypass_24_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_1_df_is_ws_5 <= io_in_r_bypass_24_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_1_stall_5 <= io_in_r_bypass_24_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_2_data_5 <= io_in_r_bypass_24_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_2_load_store_5 <= io_in_r_bypass_24_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_2_df_is_ws_5 <= io_in_r_bypass_24_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_2_stall_5 <= io_in_r_bypass_24_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_3_data_5 <= io_in_r_bypass_24_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_3_load_store_5 <= io_in_r_bypass_24_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_3_df_is_ws_5 <= io_in_r_bypass_24_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_3_stall_5 <= io_in_r_bypass_24_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_0_data_5 <= io_in_r_bypass_25_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_0_load_store_5 <= io_in_r_bypass_25_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_0_df_is_ws_5 <= io_in_r_bypass_25_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_0_stall_5 <= io_in_r_bypass_25_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_1_data_5 <= io_in_r_bypass_25_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_1_load_store_5 <= io_in_r_bypass_25_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_1_df_is_ws_5 <= io_in_r_bypass_25_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_1_stall_5 <= io_in_r_bypass_25_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_2_data_5 <= io_in_r_bypass_25_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_2_load_store_5 <= io_in_r_bypass_25_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_2_df_is_ws_5 <= io_in_r_bypass_25_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_2_stall_5 <= io_in_r_bypass_25_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_3_data_5 <= io_in_r_bypass_25_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_3_load_store_5 <= io_in_r_bypass_25_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_3_df_is_ws_5 <= io_in_r_bypass_25_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_3_stall_5 <= io_in_r_bypass_25_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_0_data_5 <= io_in_r_bypass_26_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_0_load_store_5 <= io_in_r_bypass_26_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_0_df_is_ws_5 <= io_in_r_bypass_26_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_0_stall_5 <= io_in_r_bypass_26_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_1_data_5 <= io_in_r_bypass_26_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_1_load_store_5 <= io_in_r_bypass_26_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_1_df_is_ws_5 <= io_in_r_bypass_26_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_1_stall_5 <= io_in_r_bypass_26_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_2_data_5 <= io_in_r_bypass_26_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_2_load_store_5 <= io_in_r_bypass_26_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_2_df_is_ws_5 <= io_in_r_bypass_26_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_2_stall_5 <= io_in_r_bypass_26_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_3_data_5 <= io_in_r_bypass_26_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_3_load_store_5 <= io_in_r_bypass_26_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_3_df_is_ws_5 <= io_in_r_bypass_26_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_3_stall_5 <= io_in_r_bypass_26_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_0_data_5 <= io_in_r_bypass_27_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_0_load_store_5 <= io_in_r_bypass_27_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_0_df_is_ws_5 <= io_in_r_bypass_27_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_0_stall_5 <= io_in_r_bypass_27_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_1_data_5 <= io_in_r_bypass_27_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_1_load_store_5 <= io_in_r_bypass_27_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_1_df_is_ws_5 <= io_in_r_bypass_27_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_1_stall_5 <= io_in_r_bypass_27_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_2_data_5 <= io_in_r_bypass_27_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_2_load_store_5 <= io_in_r_bypass_27_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_2_df_is_ws_5 <= io_in_r_bypass_27_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_2_stall_5 <= io_in_r_bypass_27_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_3_data_5 <= io_in_r_bypass_27_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_3_load_store_5 <= io_in_r_bypass_27_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_3_df_is_ws_5 <= io_in_r_bypass_27_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_3_stall_5 <= io_in_r_bypass_27_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_0_data_5 <= io_in_r_bypass_28_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_0_load_store_5 <= io_in_r_bypass_28_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_0_df_is_ws_5 <= io_in_r_bypass_28_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_0_stall_5 <= io_in_r_bypass_28_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_1_data_5 <= io_in_r_bypass_28_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_1_load_store_5 <= io_in_r_bypass_28_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_1_df_is_ws_5 <= io_in_r_bypass_28_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_1_stall_5 <= io_in_r_bypass_28_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_2_data_5 <= io_in_r_bypass_28_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_2_load_store_5 <= io_in_r_bypass_28_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_2_df_is_ws_5 <= io_in_r_bypass_28_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_2_stall_5 <= io_in_r_bypass_28_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_3_data_5 <= io_in_r_bypass_28_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_3_load_store_5 <= io_in_r_bypass_28_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_3_df_is_ws_5 <= io_in_r_bypass_28_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_3_stall_5 <= io_in_r_bypass_28_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_0_data_5 <= io_in_r_bypass_29_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_0_load_store_5 <= io_in_r_bypass_29_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_0_df_is_ws_5 <= io_in_r_bypass_29_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_0_stall_5 <= io_in_r_bypass_29_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_1_data_5 <= io_in_r_bypass_29_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_1_load_store_5 <= io_in_r_bypass_29_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_1_df_is_ws_5 <= io_in_r_bypass_29_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_1_stall_5 <= io_in_r_bypass_29_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_2_data_5 <= io_in_r_bypass_29_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_2_load_store_5 <= io_in_r_bypass_29_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_2_df_is_ws_5 <= io_in_r_bypass_29_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_2_stall_5 <= io_in_r_bypass_29_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_3_data_5 <= io_in_r_bypass_29_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_3_load_store_5 <= io_in_r_bypass_29_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_3_df_is_ws_5 <= io_in_r_bypass_29_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_3_stall_5 <= io_in_r_bypass_29_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_0_data_5 <= io_in_r_bypass_30_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_0_load_store_5 <= io_in_r_bypass_30_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_0_df_is_ws_5 <= io_in_r_bypass_30_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_0_stall_5 <= io_in_r_bypass_30_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_1_data_5 <= io_in_r_bypass_30_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_1_load_store_5 <= io_in_r_bypass_30_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_1_df_is_ws_5 <= io_in_r_bypass_30_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_1_stall_5 <= io_in_r_bypass_30_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_2_data_5 <= io_in_r_bypass_30_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_2_load_store_5 <= io_in_r_bypass_30_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_2_df_is_ws_5 <= io_in_r_bypass_30_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_2_stall_5 <= io_in_r_bypass_30_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_3_data_5 <= io_in_r_bypass_30_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_3_load_store_5 <= io_in_r_bypass_30_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_3_df_is_ws_5 <= io_in_r_bypass_30_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_3_stall_5 <= io_in_r_bypass_30_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_0_data_5 <= io_in_r_bypass_31_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_0_load_store_5 <= io_in_r_bypass_31_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_0_df_is_ws_5 <= io_in_r_bypass_31_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_0_stall_5 <= io_in_r_bypass_31_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_1_data_5 <= io_in_r_bypass_31_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_1_load_store_5 <= io_in_r_bypass_31_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_1_df_is_ws_5 <= io_in_r_bypass_31_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_1_stall_5 <= io_in_r_bypass_31_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_2_data_5 <= io_in_r_bypass_31_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_2_load_store_5 <= io_in_r_bypass_31_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_2_df_is_ws_5 <= io_in_r_bypass_31_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_2_stall_5 <= io_in_r_bypass_31_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_3_data_5 <= io_in_r_bypass_31_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_3_load_store_5 <= io_in_r_bypass_31_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_3_df_is_ws_5 <= io_in_r_bypass_31_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_3_stall_5 <= io_in_r_bypass_31_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_0_data_6 <= io_in_r_bypass_0_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_0_load_store_6 <= io_in_r_bypass_0_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_0_df_is_ws_6 <= io_in_r_bypass_0_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_0_stall_6 <= io_in_r_bypass_0_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_1_data_6 <= io_in_r_bypass_0_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_1_load_store_6 <= io_in_r_bypass_0_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_1_df_is_ws_6 <= io_in_r_bypass_0_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_1_stall_6 <= io_in_r_bypass_0_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_2_data_6 <= io_in_r_bypass_0_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_2_load_store_6 <= io_in_r_bypass_0_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_2_df_is_ws_6 <= io_in_r_bypass_0_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_2_stall_6 <= io_in_r_bypass_0_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_3_data_6 <= io_in_r_bypass_0_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_3_load_store_6 <= io_in_r_bypass_0_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_3_df_is_ws_6 <= io_in_r_bypass_0_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_3_stall_6 <= io_in_r_bypass_0_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_0_data_6 <= io_in_r_bypass_1_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_0_load_store_6 <= io_in_r_bypass_1_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_0_df_is_ws_6 <= io_in_r_bypass_1_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_0_stall_6 <= io_in_r_bypass_1_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_1_data_6 <= io_in_r_bypass_1_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_1_load_store_6 <= io_in_r_bypass_1_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_1_df_is_ws_6 <= io_in_r_bypass_1_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_1_stall_6 <= io_in_r_bypass_1_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_2_data_6 <= io_in_r_bypass_1_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_2_load_store_6 <= io_in_r_bypass_1_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_2_df_is_ws_6 <= io_in_r_bypass_1_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_2_stall_6 <= io_in_r_bypass_1_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_3_data_6 <= io_in_r_bypass_1_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_3_load_store_6 <= io_in_r_bypass_1_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_3_df_is_ws_6 <= io_in_r_bypass_1_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_3_stall_6 <= io_in_r_bypass_1_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_0_data_6 <= io_in_r_bypass_2_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_0_load_store_6 <= io_in_r_bypass_2_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_0_df_is_ws_6 <= io_in_r_bypass_2_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_0_stall_6 <= io_in_r_bypass_2_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_1_data_6 <= io_in_r_bypass_2_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_1_load_store_6 <= io_in_r_bypass_2_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_1_df_is_ws_6 <= io_in_r_bypass_2_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_1_stall_6 <= io_in_r_bypass_2_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_2_data_6 <= io_in_r_bypass_2_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_2_load_store_6 <= io_in_r_bypass_2_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_2_df_is_ws_6 <= io_in_r_bypass_2_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_2_stall_6 <= io_in_r_bypass_2_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_3_data_6 <= io_in_r_bypass_2_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_3_load_store_6 <= io_in_r_bypass_2_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_3_df_is_ws_6 <= io_in_r_bypass_2_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_3_stall_6 <= io_in_r_bypass_2_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_0_data_6 <= io_in_r_bypass_3_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_0_load_store_6 <= io_in_r_bypass_3_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_0_df_is_ws_6 <= io_in_r_bypass_3_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_0_stall_6 <= io_in_r_bypass_3_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_1_data_6 <= io_in_r_bypass_3_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_1_load_store_6 <= io_in_r_bypass_3_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_1_df_is_ws_6 <= io_in_r_bypass_3_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_1_stall_6 <= io_in_r_bypass_3_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_2_data_6 <= io_in_r_bypass_3_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_2_load_store_6 <= io_in_r_bypass_3_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_2_df_is_ws_6 <= io_in_r_bypass_3_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_2_stall_6 <= io_in_r_bypass_3_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_3_data_6 <= io_in_r_bypass_3_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_3_load_store_6 <= io_in_r_bypass_3_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_3_df_is_ws_6 <= io_in_r_bypass_3_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_3_stall_6 <= io_in_r_bypass_3_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_0_data_6 <= io_in_r_bypass_4_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_0_load_store_6 <= io_in_r_bypass_4_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_0_df_is_ws_6 <= io_in_r_bypass_4_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_0_stall_6 <= io_in_r_bypass_4_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_1_data_6 <= io_in_r_bypass_4_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_1_load_store_6 <= io_in_r_bypass_4_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_1_df_is_ws_6 <= io_in_r_bypass_4_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_1_stall_6 <= io_in_r_bypass_4_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_2_data_6 <= io_in_r_bypass_4_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_2_load_store_6 <= io_in_r_bypass_4_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_2_df_is_ws_6 <= io_in_r_bypass_4_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_2_stall_6 <= io_in_r_bypass_4_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_3_data_6 <= io_in_r_bypass_4_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_3_load_store_6 <= io_in_r_bypass_4_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_3_df_is_ws_6 <= io_in_r_bypass_4_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_3_stall_6 <= io_in_r_bypass_4_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_0_data_6 <= io_in_r_bypass_5_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_0_load_store_6 <= io_in_r_bypass_5_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_0_df_is_ws_6 <= io_in_r_bypass_5_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_0_stall_6 <= io_in_r_bypass_5_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_1_data_6 <= io_in_r_bypass_5_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_1_load_store_6 <= io_in_r_bypass_5_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_1_df_is_ws_6 <= io_in_r_bypass_5_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_1_stall_6 <= io_in_r_bypass_5_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_2_data_6 <= io_in_r_bypass_5_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_2_load_store_6 <= io_in_r_bypass_5_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_2_df_is_ws_6 <= io_in_r_bypass_5_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_2_stall_6 <= io_in_r_bypass_5_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_3_data_6 <= io_in_r_bypass_5_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_3_load_store_6 <= io_in_r_bypass_5_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_3_df_is_ws_6 <= io_in_r_bypass_5_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_3_stall_6 <= io_in_r_bypass_5_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_0_data_6 <= io_in_r_bypass_6_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_0_load_store_6 <= io_in_r_bypass_6_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_0_df_is_ws_6 <= io_in_r_bypass_6_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_0_stall_6 <= io_in_r_bypass_6_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_1_data_6 <= io_in_r_bypass_6_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_1_load_store_6 <= io_in_r_bypass_6_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_1_df_is_ws_6 <= io_in_r_bypass_6_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_1_stall_6 <= io_in_r_bypass_6_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_2_data_6 <= io_in_r_bypass_6_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_2_load_store_6 <= io_in_r_bypass_6_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_2_df_is_ws_6 <= io_in_r_bypass_6_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_2_stall_6 <= io_in_r_bypass_6_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_3_data_6 <= io_in_r_bypass_6_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_3_load_store_6 <= io_in_r_bypass_6_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_3_df_is_ws_6 <= io_in_r_bypass_6_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_3_stall_6 <= io_in_r_bypass_6_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_0_data_6 <= io_in_r_bypass_7_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_0_load_store_6 <= io_in_r_bypass_7_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_0_df_is_ws_6 <= io_in_r_bypass_7_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_0_stall_6 <= io_in_r_bypass_7_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_1_data_6 <= io_in_r_bypass_7_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_1_load_store_6 <= io_in_r_bypass_7_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_1_df_is_ws_6 <= io_in_r_bypass_7_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_1_stall_6 <= io_in_r_bypass_7_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_2_data_6 <= io_in_r_bypass_7_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_2_load_store_6 <= io_in_r_bypass_7_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_2_df_is_ws_6 <= io_in_r_bypass_7_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_2_stall_6 <= io_in_r_bypass_7_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_3_data_6 <= io_in_r_bypass_7_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_3_load_store_6 <= io_in_r_bypass_7_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_3_df_is_ws_6 <= io_in_r_bypass_7_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_3_stall_6 <= io_in_r_bypass_7_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_0_data_6 <= io_in_r_bypass_8_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_0_load_store_6 <= io_in_r_bypass_8_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_0_df_is_ws_6 <= io_in_r_bypass_8_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_0_stall_6 <= io_in_r_bypass_8_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_1_data_6 <= io_in_r_bypass_8_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_1_load_store_6 <= io_in_r_bypass_8_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_1_df_is_ws_6 <= io_in_r_bypass_8_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_1_stall_6 <= io_in_r_bypass_8_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_2_data_6 <= io_in_r_bypass_8_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_2_load_store_6 <= io_in_r_bypass_8_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_2_df_is_ws_6 <= io_in_r_bypass_8_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_2_stall_6 <= io_in_r_bypass_8_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_3_data_6 <= io_in_r_bypass_8_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_3_load_store_6 <= io_in_r_bypass_8_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_3_df_is_ws_6 <= io_in_r_bypass_8_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_3_stall_6 <= io_in_r_bypass_8_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_0_data_6 <= io_in_r_bypass_9_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_0_load_store_6 <= io_in_r_bypass_9_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_0_df_is_ws_6 <= io_in_r_bypass_9_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_0_stall_6 <= io_in_r_bypass_9_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_1_data_6 <= io_in_r_bypass_9_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_1_load_store_6 <= io_in_r_bypass_9_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_1_df_is_ws_6 <= io_in_r_bypass_9_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_1_stall_6 <= io_in_r_bypass_9_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_2_data_6 <= io_in_r_bypass_9_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_2_load_store_6 <= io_in_r_bypass_9_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_2_df_is_ws_6 <= io_in_r_bypass_9_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_2_stall_6 <= io_in_r_bypass_9_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_3_data_6 <= io_in_r_bypass_9_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_3_load_store_6 <= io_in_r_bypass_9_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_3_df_is_ws_6 <= io_in_r_bypass_9_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_3_stall_6 <= io_in_r_bypass_9_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_0_data_6 <= io_in_r_bypass_10_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_0_load_store_6 <= io_in_r_bypass_10_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_0_df_is_ws_6 <= io_in_r_bypass_10_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_0_stall_6 <= io_in_r_bypass_10_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_1_data_6 <= io_in_r_bypass_10_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_1_load_store_6 <= io_in_r_bypass_10_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_1_df_is_ws_6 <= io_in_r_bypass_10_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_1_stall_6 <= io_in_r_bypass_10_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_2_data_6 <= io_in_r_bypass_10_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_2_load_store_6 <= io_in_r_bypass_10_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_2_df_is_ws_6 <= io_in_r_bypass_10_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_2_stall_6 <= io_in_r_bypass_10_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_3_data_6 <= io_in_r_bypass_10_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_3_load_store_6 <= io_in_r_bypass_10_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_3_df_is_ws_6 <= io_in_r_bypass_10_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_3_stall_6 <= io_in_r_bypass_10_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_0_data_6 <= io_in_r_bypass_11_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_0_load_store_6 <= io_in_r_bypass_11_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_0_df_is_ws_6 <= io_in_r_bypass_11_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_0_stall_6 <= io_in_r_bypass_11_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_1_data_6 <= io_in_r_bypass_11_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_1_load_store_6 <= io_in_r_bypass_11_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_1_df_is_ws_6 <= io_in_r_bypass_11_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_1_stall_6 <= io_in_r_bypass_11_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_2_data_6 <= io_in_r_bypass_11_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_2_load_store_6 <= io_in_r_bypass_11_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_2_df_is_ws_6 <= io_in_r_bypass_11_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_2_stall_6 <= io_in_r_bypass_11_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_3_data_6 <= io_in_r_bypass_11_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_3_load_store_6 <= io_in_r_bypass_11_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_3_df_is_ws_6 <= io_in_r_bypass_11_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_3_stall_6 <= io_in_r_bypass_11_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_0_data_6 <= io_in_r_bypass_12_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_0_load_store_6 <= io_in_r_bypass_12_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_0_df_is_ws_6 <= io_in_r_bypass_12_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_0_stall_6 <= io_in_r_bypass_12_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_1_data_6 <= io_in_r_bypass_12_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_1_load_store_6 <= io_in_r_bypass_12_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_1_df_is_ws_6 <= io_in_r_bypass_12_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_1_stall_6 <= io_in_r_bypass_12_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_2_data_6 <= io_in_r_bypass_12_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_2_load_store_6 <= io_in_r_bypass_12_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_2_df_is_ws_6 <= io_in_r_bypass_12_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_2_stall_6 <= io_in_r_bypass_12_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_3_data_6 <= io_in_r_bypass_12_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_3_load_store_6 <= io_in_r_bypass_12_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_3_df_is_ws_6 <= io_in_r_bypass_12_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_3_stall_6 <= io_in_r_bypass_12_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_0_data_6 <= io_in_r_bypass_13_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_0_load_store_6 <= io_in_r_bypass_13_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_0_df_is_ws_6 <= io_in_r_bypass_13_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_0_stall_6 <= io_in_r_bypass_13_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_1_data_6 <= io_in_r_bypass_13_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_1_load_store_6 <= io_in_r_bypass_13_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_1_df_is_ws_6 <= io_in_r_bypass_13_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_1_stall_6 <= io_in_r_bypass_13_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_2_data_6 <= io_in_r_bypass_13_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_2_load_store_6 <= io_in_r_bypass_13_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_2_df_is_ws_6 <= io_in_r_bypass_13_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_2_stall_6 <= io_in_r_bypass_13_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_3_data_6 <= io_in_r_bypass_13_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_3_load_store_6 <= io_in_r_bypass_13_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_3_df_is_ws_6 <= io_in_r_bypass_13_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_3_stall_6 <= io_in_r_bypass_13_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_0_data_6 <= io_in_r_bypass_14_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_0_load_store_6 <= io_in_r_bypass_14_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_0_df_is_ws_6 <= io_in_r_bypass_14_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_0_stall_6 <= io_in_r_bypass_14_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_1_data_6 <= io_in_r_bypass_14_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_1_load_store_6 <= io_in_r_bypass_14_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_1_df_is_ws_6 <= io_in_r_bypass_14_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_1_stall_6 <= io_in_r_bypass_14_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_2_data_6 <= io_in_r_bypass_14_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_2_load_store_6 <= io_in_r_bypass_14_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_2_df_is_ws_6 <= io_in_r_bypass_14_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_2_stall_6 <= io_in_r_bypass_14_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_3_data_6 <= io_in_r_bypass_14_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_3_load_store_6 <= io_in_r_bypass_14_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_3_df_is_ws_6 <= io_in_r_bypass_14_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_3_stall_6 <= io_in_r_bypass_14_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_0_data_6 <= io_in_r_bypass_15_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_0_load_store_6 <= io_in_r_bypass_15_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_0_df_is_ws_6 <= io_in_r_bypass_15_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_0_stall_6 <= io_in_r_bypass_15_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_1_data_6 <= io_in_r_bypass_15_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_1_load_store_6 <= io_in_r_bypass_15_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_1_df_is_ws_6 <= io_in_r_bypass_15_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_1_stall_6 <= io_in_r_bypass_15_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_2_data_6 <= io_in_r_bypass_15_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_2_load_store_6 <= io_in_r_bypass_15_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_2_df_is_ws_6 <= io_in_r_bypass_15_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_2_stall_6 <= io_in_r_bypass_15_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_3_data_6 <= io_in_r_bypass_15_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_3_load_store_6 <= io_in_r_bypass_15_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_3_df_is_ws_6 <= io_in_r_bypass_15_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_3_stall_6 <= io_in_r_bypass_15_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_0_data_6 <= io_in_r_bypass_16_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_0_load_store_6 <= io_in_r_bypass_16_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_0_df_is_ws_6 <= io_in_r_bypass_16_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_0_stall_6 <= io_in_r_bypass_16_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_1_data_6 <= io_in_r_bypass_16_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_1_load_store_6 <= io_in_r_bypass_16_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_1_df_is_ws_6 <= io_in_r_bypass_16_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_1_stall_6 <= io_in_r_bypass_16_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_2_data_6 <= io_in_r_bypass_16_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_2_load_store_6 <= io_in_r_bypass_16_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_2_df_is_ws_6 <= io_in_r_bypass_16_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_2_stall_6 <= io_in_r_bypass_16_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_3_data_6 <= io_in_r_bypass_16_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_3_load_store_6 <= io_in_r_bypass_16_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_3_df_is_ws_6 <= io_in_r_bypass_16_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_3_stall_6 <= io_in_r_bypass_16_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_0_data_6 <= io_in_r_bypass_17_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_0_load_store_6 <= io_in_r_bypass_17_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_0_df_is_ws_6 <= io_in_r_bypass_17_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_0_stall_6 <= io_in_r_bypass_17_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_1_data_6 <= io_in_r_bypass_17_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_1_load_store_6 <= io_in_r_bypass_17_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_1_df_is_ws_6 <= io_in_r_bypass_17_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_1_stall_6 <= io_in_r_bypass_17_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_2_data_6 <= io_in_r_bypass_17_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_2_load_store_6 <= io_in_r_bypass_17_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_2_df_is_ws_6 <= io_in_r_bypass_17_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_2_stall_6 <= io_in_r_bypass_17_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_3_data_6 <= io_in_r_bypass_17_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_3_load_store_6 <= io_in_r_bypass_17_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_3_df_is_ws_6 <= io_in_r_bypass_17_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_3_stall_6 <= io_in_r_bypass_17_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_0_data_6 <= io_in_r_bypass_18_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_0_load_store_6 <= io_in_r_bypass_18_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_0_df_is_ws_6 <= io_in_r_bypass_18_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_0_stall_6 <= io_in_r_bypass_18_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_1_data_6 <= io_in_r_bypass_18_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_1_load_store_6 <= io_in_r_bypass_18_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_1_df_is_ws_6 <= io_in_r_bypass_18_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_1_stall_6 <= io_in_r_bypass_18_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_2_data_6 <= io_in_r_bypass_18_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_2_load_store_6 <= io_in_r_bypass_18_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_2_df_is_ws_6 <= io_in_r_bypass_18_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_2_stall_6 <= io_in_r_bypass_18_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_3_data_6 <= io_in_r_bypass_18_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_3_load_store_6 <= io_in_r_bypass_18_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_3_df_is_ws_6 <= io_in_r_bypass_18_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_3_stall_6 <= io_in_r_bypass_18_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_0_data_6 <= io_in_r_bypass_19_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_0_load_store_6 <= io_in_r_bypass_19_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_0_df_is_ws_6 <= io_in_r_bypass_19_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_0_stall_6 <= io_in_r_bypass_19_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_1_data_6 <= io_in_r_bypass_19_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_1_load_store_6 <= io_in_r_bypass_19_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_1_df_is_ws_6 <= io_in_r_bypass_19_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_1_stall_6 <= io_in_r_bypass_19_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_2_data_6 <= io_in_r_bypass_19_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_2_load_store_6 <= io_in_r_bypass_19_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_2_df_is_ws_6 <= io_in_r_bypass_19_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_2_stall_6 <= io_in_r_bypass_19_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_3_data_6 <= io_in_r_bypass_19_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_3_load_store_6 <= io_in_r_bypass_19_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_3_df_is_ws_6 <= io_in_r_bypass_19_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_3_stall_6 <= io_in_r_bypass_19_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_0_data_6 <= io_in_r_bypass_20_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_0_load_store_6 <= io_in_r_bypass_20_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_0_df_is_ws_6 <= io_in_r_bypass_20_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_0_stall_6 <= io_in_r_bypass_20_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_1_data_6 <= io_in_r_bypass_20_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_1_load_store_6 <= io_in_r_bypass_20_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_1_df_is_ws_6 <= io_in_r_bypass_20_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_1_stall_6 <= io_in_r_bypass_20_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_2_data_6 <= io_in_r_bypass_20_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_2_load_store_6 <= io_in_r_bypass_20_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_2_df_is_ws_6 <= io_in_r_bypass_20_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_2_stall_6 <= io_in_r_bypass_20_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_3_data_6 <= io_in_r_bypass_20_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_3_load_store_6 <= io_in_r_bypass_20_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_3_df_is_ws_6 <= io_in_r_bypass_20_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_3_stall_6 <= io_in_r_bypass_20_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_0_data_6 <= io_in_r_bypass_21_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_0_load_store_6 <= io_in_r_bypass_21_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_0_df_is_ws_6 <= io_in_r_bypass_21_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_0_stall_6 <= io_in_r_bypass_21_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_1_data_6 <= io_in_r_bypass_21_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_1_load_store_6 <= io_in_r_bypass_21_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_1_df_is_ws_6 <= io_in_r_bypass_21_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_1_stall_6 <= io_in_r_bypass_21_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_2_data_6 <= io_in_r_bypass_21_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_2_load_store_6 <= io_in_r_bypass_21_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_2_df_is_ws_6 <= io_in_r_bypass_21_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_2_stall_6 <= io_in_r_bypass_21_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_3_data_6 <= io_in_r_bypass_21_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_3_load_store_6 <= io_in_r_bypass_21_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_3_df_is_ws_6 <= io_in_r_bypass_21_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_3_stall_6 <= io_in_r_bypass_21_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_0_data_6 <= io_in_r_bypass_22_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_0_load_store_6 <= io_in_r_bypass_22_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_0_df_is_ws_6 <= io_in_r_bypass_22_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_0_stall_6 <= io_in_r_bypass_22_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_1_data_6 <= io_in_r_bypass_22_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_1_load_store_6 <= io_in_r_bypass_22_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_1_df_is_ws_6 <= io_in_r_bypass_22_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_1_stall_6 <= io_in_r_bypass_22_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_2_data_6 <= io_in_r_bypass_22_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_2_load_store_6 <= io_in_r_bypass_22_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_2_df_is_ws_6 <= io_in_r_bypass_22_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_2_stall_6 <= io_in_r_bypass_22_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_3_data_6 <= io_in_r_bypass_22_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_3_load_store_6 <= io_in_r_bypass_22_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_3_df_is_ws_6 <= io_in_r_bypass_22_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_3_stall_6 <= io_in_r_bypass_22_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_0_data_6 <= io_in_r_bypass_23_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_0_load_store_6 <= io_in_r_bypass_23_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_0_df_is_ws_6 <= io_in_r_bypass_23_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_0_stall_6 <= io_in_r_bypass_23_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_1_data_6 <= io_in_r_bypass_23_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_1_load_store_6 <= io_in_r_bypass_23_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_1_df_is_ws_6 <= io_in_r_bypass_23_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_1_stall_6 <= io_in_r_bypass_23_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_2_data_6 <= io_in_r_bypass_23_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_2_load_store_6 <= io_in_r_bypass_23_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_2_df_is_ws_6 <= io_in_r_bypass_23_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_2_stall_6 <= io_in_r_bypass_23_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_3_data_6 <= io_in_r_bypass_23_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_3_load_store_6 <= io_in_r_bypass_23_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_3_df_is_ws_6 <= io_in_r_bypass_23_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_3_stall_6 <= io_in_r_bypass_23_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_0_data_6 <= io_in_r_bypass_24_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_0_load_store_6 <= io_in_r_bypass_24_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_0_df_is_ws_6 <= io_in_r_bypass_24_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_0_stall_6 <= io_in_r_bypass_24_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_1_data_6 <= io_in_r_bypass_24_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_1_load_store_6 <= io_in_r_bypass_24_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_1_df_is_ws_6 <= io_in_r_bypass_24_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_1_stall_6 <= io_in_r_bypass_24_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_2_data_6 <= io_in_r_bypass_24_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_2_load_store_6 <= io_in_r_bypass_24_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_2_df_is_ws_6 <= io_in_r_bypass_24_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_2_stall_6 <= io_in_r_bypass_24_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_3_data_6 <= io_in_r_bypass_24_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_3_load_store_6 <= io_in_r_bypass_24_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_3_df_is_ws_6 <= io_in_r_bypass_24_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_3_stall_6 <= io_in_r_bypass_24_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_0_data_6 <= io_in_r_bypass_25_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_0_load_store_6 <= io_in_r_bypass_25_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_0_df_is_ws_6 <= io_in_r_bypass_25_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_0_stall_6 <= io_in_r_bypass_25_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_1_data_6 <= io_in_r_bypass_25_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_1_load_store_6 <= io_in_r_bypass_25_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_1_df_is_ws_6 <= io_in_r_bypass_25_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_1_stall_6 <= io_in_r_bypass_25_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_2_data_6 <= io_in_r_bypass_25_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_2_load_store_6 <= io_in_r_bypass_25_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_2_df_is_ws_6 <= io_in_r_bypass_25_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_2_stall_6 <= io_in_r_bypass_25_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_3_data_6 <= io_in_r_bypass_25_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_3_load_store_6 <= io_in_r_bypass_25_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_3_df_is_ws_6 <= io_in_r_bypass_25_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_3_stall_6 <= io_in_r_bypass_25_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_0_data_6 <= io_in_r_bypass_26_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_0_load_store_6 <= io_in_r_bypass_26_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_0_df_is_ws_6 <= io_in_r_bypass_26_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_0_stall_6 <= io_in_r_bypass_26_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_1_data_6 <= io_in_r_bypass_26_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_1_load_store_6 <= io_in_r_bypass_26_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_1_df_is_ws_6 <= io_in_r_bypass_26_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_1_stall_6 <= io_in_r_bypass_26_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_2_data_6 <= io_in_r_bypass_26_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_2_load_store_6 <= io_in_r_bypass_26_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_2_df_is_ws_6 <= io_in_r_bypass_26_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_2_stall_6 <= io_in_r_bypass_26_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_3_data_6 <= io_in_r_bypass_26_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_3_load_store_6 <= io_in_r_bypass_26_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_3_df_is_ws_6 <= io_in_r_bypass_26_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_3_stall_6 <= io_in_r_bypass_26_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_0_data_6 <= io_in_r_bypass_27_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_0_load_store_6 <= io_in_r_bypass_27_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_0_df_is_ws_6 <= io_in_r_bypass_27_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_0_stall_6 <= io_in_r_bypass_27_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_1_data_6 <= io_in_r_bypass_27_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_1_load_store_6 <= io_in_r_bypass_27_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_1_df_is_ws_6 <= io_in_r_bypass_27_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_1_stall_6 <= io_in_r_bypass_27_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_2_data_6 <= io_in_r_bypass_27_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_2_load_store_6 <= io_in_r_bypass_27_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_2_df_is_ws_6 <= io_in_r_bypass_27_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_2_stall_6 <= io_in_r_bypass_27_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_3_data_6 <= io_in_r_bypass_27_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_3_load_store_6 <= io_in_r_bypass_27_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_3_df_is_ws_6 <= io_in_r_bypass_27_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_3_stall_6 <= io_in_r_bypass_27_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_0_data_6 <= io_in_r_bypass_28_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_0_load_store_6 <= io_in_r_bypass_28_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_0_df_is_ws_6 <= io_in_r_bypass_28_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_0_stall_6 <= io_in_r_bypass_28_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_1_data_6 <= io_in_r_bypass_28_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_1_load_store_6 <= io_in_r_bypass_28_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_1_df_is_ws_6 <= io_in_r_bypass_28_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_1_stall_6 <= io_in_r_bypass_28_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_2_data_6 <= io_in_r_bypass_28_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_2_load_store_6 <= io_in_r_bypass_28_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_2_df_is_ws_6 <= io_in_r_bypass_28_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_2_stall_6 <= io_in_r_bypass_28_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_3_data_6 <= io_in_r_bypass_28_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_3_load_store_6 <= io_in_r_bypass_28_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_3_df_is_ws_6 <= io_in_r_bypass_28_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_3_stall_6 <= io_in_r_bypass_28_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_0_data_6 <= io_in_r_bypass_29_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_0_load_store_6 <= io_in_r_bypass_29_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_0_df_is_ws_6 <= io_in_r_bypass_29_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_0_stall_6 <= io_in_r_bypass_29_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_1_data_6 <= io_in_r_bypass_29_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_1_load_store_6 <= io_in_r_bypass_29_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_1_df_is_ws_6 <= io_in_r_bypass_29_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_1_stall_6 <= io_in_r_bypass_29_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_2_data_6 <= io_in_r_bypass_29_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_2_load_store_6 <= io_in_r_bypass_29_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_2_df_is_ws_6 <= io_in_r_bypass_29_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_2_stall_6 <= io_in_r_bypass_29_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_3_data_6 <= io_in_r_bypass_29_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_3_load_store_6 <= io_in_r_bypass_29_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_3_df_is_ws_6 <= io_in_r_bypass_29_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_3_stall_6 <= io_in_r_bypass_29_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_0_data_6 <= io_in_r_bypass_30_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_0_load_store_6 <= io_in_r_bypass_30_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_0_df_is_ws_6 <= io_in_r_bypass_30_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_0_stall_6 <= io_in_r_bypass_30_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_1_data_6 <= io_in_r_bypass_30_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_1_load_store_6 <= io_in_r_bypass_30_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_1_df_is_ws_6 <= io_in_r_bypass_30_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_1_stall_6 <= io_in_r_bypass_30_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_2_data_6 <= io_in_r_bypass_30_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_2_load_store_6 <= io_in_r_bypass_30_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_2_df_is_ws_6 <= io_in_r_bypass_30_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_2_stall_6 <= io_in_r_bypass_30_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_3_data_6 <= io_in_r_bypass_30_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_3_load_store_6 <= io_in_r_bypass_30_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_3_df_is_ws_6 <= io_in_r_bypass_30_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_3_stall_6 <= io_in_r_bypass_30_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_0_data_6 <= io_in_r_bypass_31_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_0_load_store_6 <= io_in_r_bypass_31_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_0_df_is_ws_6 <= io_in_r_bypass_31_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_0_stall_6 <= io_in_r_bypass_31_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_1_data_6 <= io_in_r_bypass_31_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_1_load_store_6 <= io_in_r_bypass_31_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_1_df_is_ws_6 <= io_in_r_bypass_31_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_1_stall_6 <= io_in_r_bypass_31_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_2_data_6 <= io_in_r_bypass_31_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_2_load_store_6 <= io_in_r_bypass_31_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_2_df_is_ws_6 <= io_in_r_bypass_31_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_2_stall_6 <= io_in_r_bypass_31_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_3_data_6 <= io_in_r_bypass_31_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_3_load_store_6 <= io_in_r_bypass_31_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_3_df_is_ws_6 <= io_in_r_bypass_31_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_3_stall_6 <= io_in_r_bypass_31_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_0_data_7 <= io_in_r_bypass_0_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_0_load_store_7 <= io_in_r_bypass_0_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_0_df_is_ws_7 <= io_in_r_bypass_0_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_0_stall_7 <= io_in_r_bypass_0_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_1_data_7 <= io_in_r_bypass_0_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_1_load_store_7 <= io_in_r_bypass_0_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_1_df_is_ws_7 <= io_in_r_bypass_0_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_1_stall_7 <= io_in_r_bypass_0_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_2_data_7 <= io_in_r_bypass_0_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_2_load_store_7 <= io_in_r_bypass_0_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_2_df_is_ws_7 <= io_in_r_bypass_0_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_2_stall_7 <= io_in_r_bypass_0_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_3_data_7 <= io_in_r_bypass_0_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_3_load_store_7 <= io_in_r_bypass_0_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_3_df_is_ws_7 <= io_in_r_bypass_0_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_3_stall_7 <= io_in_r_bypass_0_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_0_data_7 <= io_in_r_bypass_1_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_0_load_store_7 <= io_in_r_bypass_1_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_0_df_is_ws_7 <= io_in_r_bypass_1_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_0_stall_7 <= io_in_r_bypass_1_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_1_data_7 <= io_in_r_bypass_1_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_1_load_store_7 <= io_in_r_bypass_1_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_1_df_is_ws_7 <= io_in_r_bypass_1_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_1_stall_7 <= io_in_r_bypass_1_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_2_data_7 <= io_in_r_bypass_1_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_2_load_store_7 <= io_in_r_bypass_1_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_2_df_is_ws_7 <= io_in_r_bypass_1_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_2_stall_7 <= io_in_r_bypass_1_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_3_data_7 <= io_in_r_bypass_1_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_3_load_store_7 <= io_in_r_bypass_1_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_3_df_is_ws_7 <= io_in_r_bypass_1_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_3_stall_7 <= io_in_r_bypass_1_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_0_data_7 <= io_in_r_bypass_2_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_0_load_store_7 <= io_in_r_bypass_2_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_0_df_is_ws_7 <= io_in_r_bypass_2_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_0_stall_7 <= io_in_r_bypass_2_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_1_data_7 <= io_in_r_bypass_2_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_1_load_store_7 <= io_in_r_bypass_2_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_1_df_is_ws_7 <= io_in_r_bypass_2_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_1_stall_7 <= io_in_r_bypass_2_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_2_data_7 <= io_in_r_bypass_2_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_2_load_store_7 <= io_in_r_bypass_2_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_2_df_is_ws_7 <= io_in_r_bypass_2_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_2_stall_7 <= io_in_r_bypass_2_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_3_data_7 <= io_in_r_bypass_2_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_3_load_store_7 <= io_in_r_bypass_2_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_3_df_is_ws_7 <= io_in_r_bypass_2_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_3_stall_7 <= io_in_r_bypass_2_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_0_data_7 <= io_in_r_bypass_3_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_0_load_store_7 <= io_in_r_bypass_3_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_0_df_is_ws_7 <= io_in_r_bypass_3_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_0_stall_7 <= io_in_r_bypass_3_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_1_data_7 <= io_in_r_bypass_3_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_1_load_store_7 <= io_in_r_bypass_3_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_1_df_is_ws_7 <= io_in_r_bypass_3_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_1_stall_7 <= io_in_r_bypass_3_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_2_data_7 <= io_in_r_bypass_3_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_2_load_store_7 <= io_in_r_bypass_3_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_2_df_is_ws_7 <= io_in_r_bypass_3_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_2_stall_7 <= io_in_r_bypass_3_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_3_data_7 <= io_in_r_bypass_3_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_3_load_store_7 <= io_in_r_bypass_3_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_3_df_is_ws_7 <= io_in_r_bypass_3_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_3_stall_7 <= io_in_r_bypass_3_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_0_data_7 <= io_in_r_bypass_4_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_0_load_store_7 <= io_in_r_bypass_4_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_0_df_is_ws_7 <= io_in_r_bypass_4_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_0_stall_7 <= io_in_r_bypass_4_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_1_data_7 <= io_in_r_bypass_4_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_1_load_store_7 <= io_in_r_bypass_4_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_1_df_is_ws_7 <= io_in_r_bypass_4_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_1_stall_7 <= io_in_r_bypass_4_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_2_data_7 <= io_in_r_bypass_4_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_2_load_store_7 <= io_in_r_bypass_4_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_2_df_is_ws_7 <= io_in_r_bypass_4_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_2_stall_7 <= io_in_r_bypass_4_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_3_data_7 <= io_in_r_bypass_4_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_3_load_store_7 <= io_in_r_bypass_4_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_3_df_is_ws_7 <= io_in_r_bypass_4_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_3_stall_7 <= io_in_r_bypass_4_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_0_data_7 <= io_in_r_bypass_5_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_0_load_store_7 <= io_in_r_bypass_5_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_0_df_is_ws_7 <= io_in_r_bypass_5_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_0_stall_7 <= io_in_r_bypass_5_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_1_data_7 <= io_in_r_bypass_5_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_1_load_store_7 <= io_in_r_bypass_5_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_1_df_is_ws_7 <= io_in_r_bypass_5_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_1_stall_7 <= io_in_r_bypass_5_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_2_data_7 <= io_in_r_bypass_5_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_2_load_store_7 <= io_in_r_bypass_5_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_2_df_is_ws_7 <= io_in_r_bypass_5_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_2_stall_7 <= io_in_r_bypass_5_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_3_data_7 <= io_in_r_bypass_5_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_3_load_store_7 <= io_in_r_bypass_5_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_3_df_is_ws_7 <= io_in_r_bypass_5_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_3_stall_7 <= io_in_r_bypass_5_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_0_data_7 <= io_in_r_bypass_6_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_0_load_store_7 <= io_in_r_bypass_6_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_0_df_is_ws_7 <= io_in_r_bypass_6_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_0_stall_7 <= io_in_r_bypass_6_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_1_data_7 <= io_in_r_bypass_6_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_1_load_store_7 <= io_in_r_bypass_6_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_1_df_is_ws_7 <= io_in_r_bypass_6_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_1_stall_7 <= io_in_r_bypass_6_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_2_data_7 <= io_in_r_bypass_6_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_2_load_store_7 <= io_in_r_bypass_6_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_2_df_is_ws_7 <= io_in_r_bypass_6_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_2_stall_7 <= io_in_r_bypass_6_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_3_data_7 <= io_in_r_bypass_6_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_3_load_store_7 <= io_in_r_bypass_6_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_3_df_is_ws_7 <= io_in_r_bypass_6_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_3_stall_7 <= io_in_r_bypass_6_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_0_data_7 <= io_in_r_bypass_7_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_0_load_store_7 <= io_in_r_bypass_7_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_0_df_is_ws_7 <= io_in_r_bypass_7_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_0_stall_7 <= io_in_r_bypass_7_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_1_data_7 <= io_in_r_bypass_7_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_1_load_store_7 <= io_in_r_bypass_7_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_1_df_is_ws_7 <= io_in_r_bypass_7_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_1_stall_7 <= io_in_r_bypass_7_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_2_data_7 <= io_in_r_bypass_7_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_2_load_store_7 <= io_in_r_bypass_7_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_2_df_is_ws_7 <= io_in_r_bypass_7_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_2_stall_7 <= io_in_r_bypass_7_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_3_data_7 <= io_in_r_bypass_7_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_3_load_store_7 <= io_in_r_bypass_7_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_3_df_is_ws_7 <= io_in_r_bypass_7_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_3_stall_7 <= io_in_r_bypass_7_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_0_data_7 <= io_in_r_bypass_8_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_0_load_store_7 <= io_in_r_bypass_8_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_0_df_is_ws_7 <= io_in_r_bypass_8_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_0_stall_7 <= io_in_r_bypass_8_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_1_data_7 <= io_in_r_bypass_8_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_1_load_store_7 <= io_in_r_bypass_8_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_1_df_is_ws_7 <= io_in_r_bypass_8_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_1_stall_7 <= io_in_r_bypass_8_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_2_data_7 <= io_in_r_bypass_8_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_2_load_store_7 <= io_in_r_bypass_8_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_2_df_is_ws_7 <= io_in_r_bypass_8_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_2_stall_7 <= io_in_r_bypass_8_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_3_data_7 <= io_in_r_bypass_8_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_3_load_store_7 <= io_in_r_bypass_8_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_3_df_is_ws_7 <= io_in_r_bypass_8_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_3_stall_7 <= io_in_r_bypass_8_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_0_data_7 <= io_in_r_bypass_9_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_0_load_store_7 <= io_in_r_bypass_9_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_0_df_is_ws_7 <= io_in_r_bypass_9_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_0_stall_7 <= io_in_r_bypass_9_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_1_data_7 <= io_in_r_bypass_9_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_1_load_store_7 <= io_in_r_bypass_9_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_1_df_is_ws_7 <= io_in_r_bypass_9_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_1_stall_7 <= io_in_r_bypass_9_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_2_data_7 <= io_in_r_bypass_9_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_2_load_store_7 <= io_in_r_bypass_9_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_2_df_is_ws_7 <= io_in_r_bypass_9_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_2_stall_7 <= io_in_r_bypass_9_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_3_data_7 <= io_in_r_bypass_9_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_3_load_store_7 <= io_in_r_bypass_9_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_3_df_is_ws_7 <= io_in_r_bypass_9_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_3_stall_7 <= io_in_r_bypass_9_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_0_data_7 <= io_in_r_bypass_10_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_0_load_store_7 <= io_in_r_bypass_10_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_0_df_is_ws_7 <= io_in_r_bypass_10_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_0_stall_7 <= io_in_r_bypass_10_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_1_data_7 <= io_in_r_bypass_10_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_1_load_store_7 <= io_in_r_bypass_10_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_1_df_is_ws_7 <= io_in_r_bypass_10_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_1_stall_7 <= io_in_r_bypass_10_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_2_data_7 <= io_in_r_bypass_10_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_2_load_store_7 <= io_in_r_bypass_10_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_2_df_is_ws_7 <= io_in_r_bypass_10_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_2_stall_7 <= io_in_r_bypass_10_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_3_data_7 <= io_in_r_bypass_10_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_3_load_store_7 <= io_in_r_bypass_10_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_3_df_is_ws_7 <= io_in_r_bypass_10_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_3_stall_7 <= io_in_r_bypass_10_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_0_data_7 <= io_in_r_bypass_11_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_0_load_store_7 <= io_in_r_bypass_11_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_0_df_is_ws_7 <= io_in_r_bypass_11_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_0_stall_7 <= io_in_r_bypass_11_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_1_data_7 <= io_in_r_bypass_11_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_1_load_store_7 <= io_in_r_bypass_11_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_1_df_is_ws_7 <= io_in_r_bypass_11_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_1_stall_7 <= io_in_r_bypass_11_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_2_data_7 <= io_in_r_bypass_11_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_2_load_store_7 <= io_in_r_bypass_11_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_2_df_is_ws_7 <= io_in_r_bypass_11_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_2_stall_7 <= io_in_r_bypass_11_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_3_data_7 <= io_in_r_bypass_11_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_3_load_store_7 <= io_in_r_bypass_11_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_3_df_is_ws_7 <= io_in_r_bypass_11_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_3_stall_7 <= io_in_r_bypass_11_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_0_data_7 <= io_in_r_bypass_12_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_0_load_store_7 <= io_in_r_bypass_12_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_0_df_is_ws_7 <= io_in_r_bypass_12_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_0_stall_7 <= io_in_r_bypass_12_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_1_data_7 <= io_in_r_bypass_12_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_1_load_store_7 <= io_in_r_bypass_12_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_1_df_is_ws_7 <= io_in_r_bypass_12_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_1_stall_7 <= io_in_r_bypass_12_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_2_data_7 <= io_in_r_bypass_12_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_2_load_store_7 <= io_in_r_bypass_12_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_2_df_is_ws_7 <= io_in_r_bypass_12_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_2_stall_7 <= io_in_r_bypass_12_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_3_data_7 <= io_in_r_bypass_12_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_3_load_store_7 <= io_in_r_bypass_12_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_3_df_is_ws_7 <= io_in_r_bypass_12_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_3_stall_7 <= io_in_r_bypass_12_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_0_data_7 <= io_in_r_bypass_13_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_0_load_store_7 <= io_in_r_bypass_13_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_0_df_is_ws_7 <= io_in_r_bypass_13_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_0_stall_7 <= io_in_r_bypass_13_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_1_data_7 <= io_in_r_bypass_13_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_1_load_store_7 <= io_in_r_bypass_13_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_1_df_is_ws_7 <= io_in_r_bypass_13_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_1_stall_7 <= io_in_r_bypass_13_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_2_data_7 <= io_in_r_bypass_13_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_2_load_store_7 <= io_in_r_bypass_13_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_2_df_is_ws_7 <= io_in_r_bypass_13_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_2_stall_7 <= io_in_r_bypass_13_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_3_data_7 <= io_in_r_bypass_13_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_3_load_store_7 <= io_in_r_bypass_13_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_3_df_is_ws_7 <= io_in_r_bypass_13_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_3_stall_7 <= io_in_r_bypass_13_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_0_data_7 <= io_in_r_bypass_14_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_0_load_store_7 <= io_in_r_bypass_14_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_0_df_is_ws_7 <= io_in_r_bypass_14_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_0_stall_7 <= io_in_r_bypass_14_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_1_data_7 <= io_in_r_bypass_14_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_1_load_store_7 <= io_in_r_bypass_14_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_1_df_is_ws_7 <= io_in_r_bypass_14_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_1_stall_7 <= io_in_r_bypass_14_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_2_data_7 <= io_in_r_bypass_14_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_2_load_store_7 <= io_in_r_bypass_14_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_2_df_is_ws_7 <= io_in_r_bypass_14_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_2_stall_7 <= io_in_r_bypass_14_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_3_data_7 <= io_in_r_bypass_14_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_3_load_store_7 <= io_in_r_bypass_14_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_3_df_is_ws_7 <= io_in_r_bypass_14_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_3_stall_7 <= io_in_r_bypass_14_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_0_data_7 <= io_in_r_bypass_15_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_0_load_store_7 <= io_in_r_bypass_15_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_0_df_is_ws_7 <= io_in_r_bypass_15_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_0_stall_7 <= io_in_r_bypass_15_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_1_data_7 <= io_in_r_bypass_15_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_1_load_store_7 <= io_in_r_bypass_15_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_1_df_is_ws_7 <= io_in_r_bypass_15_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_1_stall_7 <= io_in_r_bypass_15_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_2_data_7 <= io_in_r_bypass_15_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_2_load_store_7 <= io_in_r_bypass_15_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_2_df_is_ws_7 <= io_in_r_bypass_15_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_2_stall_7 <= io_in_r_bypass_15_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_3_data_7 <= io_in_r_bypass_15_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_3_load_store_7 <= io_in_r_bypass_15_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_3_df_is_ws_7 <= io_in_r_bypass_15_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_3_stall_7 <= io_in_r_bypass_15_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_0_data_7 <= io_in_r_bypass_16_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_0_load_store_7 <= io_in_r_bypass_16_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_0_df_is_ws_7 <= io_in_r_bypass_16_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_0_stall_7 <= io_in_r_bypass_16_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_1_data_7 <= io_in_r_bypass_16_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_1_load_store_7 <= io_in_r_bypass_16_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_1_df_is_ws_7 <= io_in_r_bypass_16_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_1_stall_7 <= io_in_r_bypass_16_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_2_data_7 <= io_in_r_bypass_16_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_2_load_store_7 <= io_in_r_bypass_16_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_2_df_is_ws_7 <= io_in_r_bypass_16_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_2_stall_7 <= io_in_r_bypass_16_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_3_data_7 <= io_in_r_bypass_16_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_3_load_store_7 <= io_in_r_bypass_16_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_3_df_is_ws_7 <= io_in_r_bypass_16_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_3_stall_7 <= io_in_r_bypass_16_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_0_data_7 <= io_in_r_bypass_17_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_0_load_store_7 <= io_in_r_bypass_17_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_0_df_is_ws_7 <= io_in_r_bypass_17_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_0_stall_7 <= io_in_r_bypass_17_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_1_data_7 <= io_in_r_bypass_17_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_1_load_store_7 <= io_in_r_bypass_17_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_1_df_is_ws_7 <= io_in_r_bypass_17_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_1_stall_7 <= io_in_r_bypass_17_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_2_data_7 <= io_in_r_bypass_17_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_2_load_store_7 <= io_in_r_bypass_17_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_2_df_is_ws_7 <= io_in_r_bypass_17_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_2_stall_7 <= io_in_r_bypass_17_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_3_data_7 <= io_in_r_bypass_17_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_3_load_store_7 <= io_in_r_bypass_17_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_3_df_is_ws_7 <= io_in_r_bypass_17_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_3_stall_7 <= io_in_r_bypass_17_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_0_data_7 <= io_in_r_bypass_18_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_0_load_store_7 <= io_in_r_bypass_18_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_0_df_is_ws_7 <= io_in_r_bypass_18_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_0_stall_7 <= io_in_r_bypass_18_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_1_data_7 <= io_in_r_bypass_18_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_1_load_store_7 <= io_in_r_bypass_18_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_1_df_is_ws_7 <= io_in_r_bypass_18_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_1_stall_7 <= io_in_r_bypass_18_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_2_data_7 <= io_in_r_bypass_18_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_2_load_store_7 <= io_in_r_bypass_18_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_2_df_is_ws_7 <= io_in_r_bypass_18_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_2_stall_7 <= io_in_r_bypass_18_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_3_data_7 <= io_in_r_bypass_18_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_3_load_store_7 <= io_in_r_bypass_18_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_3_df_is_ws_7 <= io_in_r_bypass_18_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_3_stall_7 <= io_in_r_bypass_18_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_0_data_7 <= io_in_r_bypass_19_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_0_load_store_7 <= io_in_r_bypass_19_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_0_df_is_ws_7 <= io_in_r_bypass_19_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_0_stall_7 <= io_in_r_bypass_19_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_1_data_7 <= io_in_r_bypass_19_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_1_load_store_7 <= io_in_r_bypass_19_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_1_df_is_ws_7 <= io_in_r_bypass_19_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_1_stall_7 <= io_in_r_bypass_19_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_2_data_7 <= io_in_r_bypass_19_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_2_load_store_7 <= io_in_r_bypass_19_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_2_df_is_ws_7 <= io_in_r_bypass_19_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_2_stall_7 <= io_in_r_bypass_19_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_3_data_7 <= io_in_r_bypass_19_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_3_load_store_7 <= io_in_r_bypass_19_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_3_df_is_ws_7 <= io_in_r_bypass_19_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_3_stall_7 <= io_in_r_bypass_19_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_0_data_7 <= io_in_r_bypass_20_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_0_load_store_7 <= io_in_r_bypass_20_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_0_df_is_ws_7 <= io_in_r_bypass_20_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_0_stall_7 <= io_in_r_bypass_20_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_1_data_7 <= io_in_r_bypass_20_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_1_load_store_7 <= io_in_r_bypass_20_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_1_df_is_ws_7 <= io_in_r_bypass_20_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_1_stall_7 <= io_in_r_bypass_20_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_2_data_7 <= io_in_r_bypass_20_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_2_load_store_7 <= io_in_r_bypass_20_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_2_df_is_ws_7 <= io_in_r_bypass_20_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_2_stall_7 <= io_in_r_bypass_20_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_3_data_7 <= io_in_r_bypass_20_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_3_load_store_7 <= io_in_r_bypass_20_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_3_df_is_ws_7 <= io_in_r_bypass_20_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_3_stall_7 <= io_in_r_bypass_20_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_0_data_7 <= io_in_r_bypass_21_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_0_load_store_7 <= io_in_r_bypass_21_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_0_df_is_ws_7 <= io_in_r_bypass_21_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_0_stall_7 <= io_in_r_bypass_21_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_1_data_7 <= io_in_r_bypass_21_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_1_load_store_7 <= io_in_r_bypass_21_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_1_df_is_ws_7 <= io_in_r_bypass_21_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_1_stall_7 <= io_in_r_bypass_21_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_2_data_7 <= io_in_r_bypass_21_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_2_load_store_7 <= io_in_r_bypass_21_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_2_df_is_ws_7 <= io_in_r_bypass_21_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_2_stall_7 <= io_in_r_bypass_21_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_3_data_7 <= io_in_r_bypass_21_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_3_load_store_7 <= io_in_r_bypass_21_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_3_df_is_ws_7 <= io_in_r_bypass_21_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_3_stall_7 <= io_in_r_bypass_21_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_0_data_7 <= io_in_r_bypass_22_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_0_load_store_7 <= io_in_r_bypass_22_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_0_df_is_ws_7 <= io_in_r_bypass_22_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_0_stall_7 <= io_in_r_bypass_22_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_1_data_7 <= io_in_r_bypass_22_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_1_load_store_7 <= io_in_r_bypass_22_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_1_df_is_ws_7 <= io_in_r_bypass_22_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_1_stall_7 <= io_in_r_bypass_22_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_2_data_7 <= io_in_r_bypass_22_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_2_load_store_7 <= io_in_r_bypass_22_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_2_df_is_ws_7 <= io_in_r_bypass_22_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_2_stall_7 <= io_in_r_bypass_22_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_3_data_7 <= io_in_r_bypass_22_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_3_load_store_7 <= io_in_r_bypass_22_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_3_df_is_ws_7 <= io_in_r_bypass_22_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_3_stall_7 <= io_in_r_bypass_22_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_0_data_7 <= io_in_r_bypass_23_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_0_load_store_7 <= io_in_r_bypass_23_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_0_df_is_ws_7 <= io_in_r_bypass_23_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_0_stall_7 <= io_in_r_bypass_23_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_1_data_7 <= io_in_r_bypass_23_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_1_load_store_7 <= io_in_r_bypass_23_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_1_df_is_ws_7 <= io_in_r_bypass_23_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_1_stall_7 <= io_in_r_bypass_23_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_2_data_7 <= io_in_r_bypass_23_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_2_load_store_7 <= io_in_r_bypass_23_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_2_df_is_ws_7 <= io_in_r_bypass_23_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_2_stall_7 <= io_in_r_bypass_23_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_3_data_7 <= io_in_r_bypass_23_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_3_load_store_7 <= io_in_r_bypass_23_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_3_df_is_ws_7 <= io_in_r_bypass_23_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_3_stall_7 <= io_in_r_bypass_23_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_0_data_7 <= io_in_r_bypass_24_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_0_load_store_7 <= io_in_r_bypass_24_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_0_df_is_ws_7 <= io_in_r_bypass_24_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_0_stall_7 <= io_in_r_bypass_24_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_1_data_7 <= io_in_r_bypass_24_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_1_load_store_7 <= io_in_r_bypass_24_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_1_df_is_ws_7 <= io_in_r_bypass_24_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_1_stall_7 <= io_in_r_bypass_24_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_2_data_7 <= io_in_r_bypass_24_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_2_load_store_7 <= io_in_r_bypass_24_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_2_df_is_ws_7 <= io_in_r_bypass_24_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_2_stall_7 <= io_in_r_bypass_24_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_3_data_7 <= io_in_r_bypass_24_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_3_load_store_7 <= io_in_r_bypass_24_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_3_df_is_ws_7 <= io_in_r_bypass_24_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_3_stall_7 <= io_in_r_bypass_24_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_0_data_7 <= io_in_r_bypass_25_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_0_load_store_7 <= io_in_r_bypass_25_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_0_df_is_ws_7 <= io_in_r_bypass_25_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_0_stall_7 <= io_in_r_bypass_25_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_1_data_7 <= io_in_r_bypass_25_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_1_load_store_7 <= io_in_r_bypass_25_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_1_df_is_ws_7 <= io_in_r_bypass_25_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_1_stall_7 <= io_in_r_bypass_25_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_2_data_7 <= io_in_r_bypass_25_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_2_load_store_7 <= io_in_r_bypass_25_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_2_df_is_ws_7 <= io_in_r_bypass_25_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_2_stall_7 <= io_in_r_bypass_25_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_3_data_7 <= io_in_r_bypass_25_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_3_load_store_7 <= io_in_r_bypass_25_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_3_df_is_ws_7 <= io_in_r_bypass_25_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_3_stall_7 <= io_in_r_bypass_25_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_0_data_7 <= io_in_r_bypass_26_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_0_load_store_7 <= io_in_r_bypass_26_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_0_df_is_ws_7 <= io_in_r_bypass_26_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_0_stall_7 <= io_in_r_bypass_26_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_1_data_7 <= io_in_r_bypass_26_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_1_load_store_7 <= io_in_r_bypass_26_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_1_df_is_ws_7 <= io_in_r_bypass_26_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_1_stall_7 <= io_in_r_bypass_26_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_2_data_7 <= io_in_r_bypass_26_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_2_load_store_7 <= io_in_r_bypass_26_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_2_df_is_ws_7 <= io_in_r_bypass_26_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_2_stall_7 <= io_in_r_bypass_26_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_3_data_7 <= io_in_r_bypass_26_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_3_load_store_7 <= io_in_r_bypass_26_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_3_df_is_ws_7 <= io_in_r_bypass_26_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_3_stall_7 <= io_in_r_bypass_26_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_0_data_7 <= io_in_r_bypass_27_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_0_load_store_7 <= io_in_r_bypass_27_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_0_df_is_ws_7 <= io_in_r_bypass_27_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_0_stall_7 <= io_in_r_bypass_27_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_1_data_7 <= io_in_r_bypass_27_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_1_load_store_7 <= io_in_r_bypass_27_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_1_df_is_ws_7 <= io_in_r_bypass_27_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_1_stall_7 <= io_in_r_bypass_27_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_2_data_7 <= io_in_r_bypass_27_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_2_load_store_7 <= io_in_r_bypass_27_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_2_df_is_ws_7 <= io_in_r_bypass_27_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_2_stall_7 <= io_in_r_bypass_27_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_3_data_7 <= io_in_r_bypass_27_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_3_load_store_7 <= io_in_r_bypass_27_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_3_df_is_ws_7 <= io_in_r_bypass_27_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_3_stall_7 <= io_in_r_bypass_27_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_0_data_7 <= io_in_r_bypass_28_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_0_load_store_7 <= io_in_r_bypass_28_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_0_df_is_ws_7 <= io_in_r_bypass_28_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_0_stall_7 <= io_in_r_bypass_28_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_1_data_7 <= io_in_r_bypass_28_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_1_load_store_7 <= io_in_r_bypass_28_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_1_df_is_ws_7 <= io_in_r_bypass_28_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_1_stall_7 <= io_in_r_bypass_28_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_2_data_7 <= io_in_r_bypass_28_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_2_load_store_7 <= io_in_r_bypass_28_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_2_df_is_ws_7 <= io_in_r_bypass_28_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_2_stall_7 <= io_in_r_bypass_28_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_3_data_7 <= io_in_r_bypass_28_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_3_load_store_7 <= io_in_r_bypass_28_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_3_df_is_ws_7 <= io_in_r_bypass_28_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_3_stall_7 <= io_in_r_bypass_28_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_0_data_7 <= io_in_r_bypass_29_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_0_load_store_7 <= io_in_r_bypass_29_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_0_df_is_ws_7 <= io_in_r_bypass_29_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_0_stall_7 <= io_in_r_bypass_29_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_1_data_7 <= io_in_r_bypass_29_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_1_load_store_7 <= io_in_r_bypass_29_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_1_df_is_ws_7 <= io_in_r_bypass_29_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_1_stall_7 <= io_in_r_bypass_29_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_2_data_7 <= io_in_r_bypass_29_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_2_load_store_7 <= io_in_r_bypass_29_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_2_df_is_ws_7 <= io_in_r_bypass_29_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_2_stall_7 <= io_in_r_bypass_29_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_3_data_7 <= io_in_r_bypass_29_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_3_load_store_7 <= io_in_r_bypass_29_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_3_df_is_ws_7 <= io_in_r_bypass_29_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_3_stall_7 <= io_in_r_bypass_29_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_0_data_7 <= io_in_r_bypass_30_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_0_load_store_7 <= io_in_r_bypass_30_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_0_df_is_ws_7 <= io_in_r_bypass_30_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_0_stall_7 <= io_in_r_bypass_30_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_1_data_7 <= io_in_r_bypass_30_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_1_load_store_7 <= io_in_r_bypass_30_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_1_df_is_ws_7 <= io_in_r_bypass_30_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_1_stall_7 <= io_in_r_bypass_30_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_2_data_7 <= io_in_r_bypass_30_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_2_load_store_7 <= io_in_r_bypass_30_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_2_df_is_ws_7 <= io_in_r_bypass_30_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_2_stall_7 <= io_in_r_bypass_30_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_3_data_7 <= io_in_r_bypass_30_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_3_load_store_7 <= io_in_r_bypass_30_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_3_df_is_ws_7 <= io_in_r_bypass_30_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_3_stall_7 <= io_in_r_bypass_30_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_0_data_7 <= io_in_r_bypass_31_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_0_load_store_7 <= io_in_r_bypass_31_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_0_df_is_ws_7 <= io_in_r_bypass_31_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_0_stall_7 <= io_in_r_bypass_31_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_1_data_7 <= io_in_r_bypass_31_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_1_load_store_7 <= io_in_r_bypass_31_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_1_df_is_ws_7 <= io_in_r_bypass_31_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_1_stall_7 <= io_in_r_bypass_31_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_2_data_7 <= io_in_r_bypass_31_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_2_load_store_7 <= io_in_r_bypass_31_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_2_df_is_ws_7 <= io_in_r_bypass_31_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_2_stall_7 <= io_in_r_bypass_31_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_3_data_7 <= io_in_r_bypass_31_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_3_load_store_7 <= io_in_r_bypass_31_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_3_df_is_ws_7 <= io_in_r_bypass_31_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_3_stall_7 <= io_in_r_bypass_31_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_0_data_8 <= io_in_r_bypass_0_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_0_load_store_8 <= io_in_r_bypass_0_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_0_df_is_ws_8 <= io_in_r_bypass_0_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_0_stall_8 <= io_in_r_bypass_0_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_1_data_8 <= io_in_r_bypass_0_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_1_load_store_8 <= io_in_r_bypass_0_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_1_df_is_ws_8 <= io_in_r_bypass_0_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_1_stall_8 <= io_in_r_bypass_0_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_2_data_8 <= io_in_r_bypass_0_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_2_load_store_8 <= io_in_r_bypass_0_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_2_df_is_ws_8 <= io_in_r_bypass_0_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_2_stall_8 <= io_in_r_bypass_0_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_3_data_8 <= io_in_r_bypass_0_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_3_load_store_8 <= io_in_r_bypass_0_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_3_df_is_ws_8 <= io_in_r_bypass_0_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_3_stall_8 <= io_in_r_bypass_0_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_0_data_8 <= io_in_r_bypass_1_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_0_load_store_8 <= io_in_r_bypass_1_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_0_df_is_ws_8 <= io_in_r_bypass_1_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_0_stall_8 <= io_in_r_bypass_1_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_1_data_8 <= io_in_r_bypass_1_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_1_load_store_8 <= io_in_r_bypass_1_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_1_df_is_ws_8 <= io_in_r_bypass_1_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_1_stall_8 <= io_in_r_bypass_1_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_2_data_8 <= io_in_r_bypass_1_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_2_load_store_8 <= io_in_r_bypass_1_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_2_df_is_ws_8 <= io_in_r_bypass_1_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_2_stall_8 <= io_in_r_bypass_1_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_3_data_8 <= io_in_r_bypass_1_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_3_load_store_8 <= io_in_r_bypass_1_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_3_df_is_ws_8 <= io_in_r_bypass_1_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_3_stall_8 <= io_in_r_bypass_1_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_0_data_8 <= io_in_r_bypass_2_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_0_load_store_8 <= io_in_r_bypass_2_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_0_df_is_ws_8 <= io_in_r_bypass_2_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_0_stall_8 <= io_in_r_bypass_2_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_1_data_8 <= io_in_r_bypass_2_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_1_load_store_8 <= io_in_r_bypass_2_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_1_df_is_ws_8 <= io_in_r_bypass_2_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_1_stall_8 <= io_in_r_bypass_2_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_2_data_8 <= io_in_r_bypass_2_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_2_load_store_8 <= io_in_r_bypass_2_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_2_df_is_ws_8 <= io_in_r_bypass_2_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_2_stall_8 <= io_in_r_bypass_2_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_3_data_8 <= io_in_r_bypass_2_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_3_load_store_8 <= io_in_r_bypass_2_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_3_df_is_ws_8 <= io_in_r_bypass_2_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_3_stall_8 <= io_in_r_bypass_2_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_0_data_8 <= io_in_r_bypass_3_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_0_load_store_8 <= io_in_r_bypass_3_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_0_df_is_ws_8 <= io_in_r_bypass_3_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_0_stall_8 <= io_in_r_bypass_3_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_1_data_8 <= io_in_r_bypass_3_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_1_load_store_8 <= io_in_r_bypass_3_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_1_df_is_ws_8 <= io_in_r_bypass_3_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_1_stall_8 <= io_in_r_bypass_3_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_2_data_8 <= io_in_r_bypass_3_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_2_load_store_8 <= io_in_r_bypass_3_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_2_df_is_ws_8 <= io_in_r_bypass_3_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_2_stall_8 <= io_in_r_bypass_3_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_3_data_8 <= io_in_r_bypass_3_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_3_load_store_8 <= io_in_r_bypass_3_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_3_df_is_ws_8 <= io_in_r_bypass_3_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_3_stall_8 <= io_in_r_bypass_3_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_0_data_8 <= io_in_r_bypass_4_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_0_load_store_8 <= io_in_r_bypass_4_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_0_df_is_ws_8 <= io_in_r_bypass_4_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_0_stall_8 <= io_in_r_bypass_4_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_1_data_8 <= io_in_r_bypass_4_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_1_load_store_8 <= io_in_r_bypass_4_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_1_df_is_ws_8 <= io_in_r_bypass_4_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_1_stall_8 <= io_in_r_bypass_4_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_2_data_8 <= io_in_r_bypass_4_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_2_load_store_8 <= io_in_r_bypass_4_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_2_df_is_ws_8 <= io_in_r_bypass_4_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_2_stall_8 <= io_in_r_bypass_4_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_3_data_8 <= io_in_r_bypass_4_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_3_load_store_8 <= io_in_r_bypass_4_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_3_df_is_ws_8 <= io_in_r_bypass_4_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_3_stall_8 <= io_in_r_bypass_4_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_0_data_8 <= io_in_r_bypass_5_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_0_load_store_8 <= io_in_r_bypass_5_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_0_df_is_ws_8 <= io_in_r_bypass_5_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_0_stall_8 <= io_in_r_bypass_5_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_1_data_8 <= io_in_r_bypass_5_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_1_load_store_8 <= io_in_r_bypass_5_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_1_df_is_ws_8 <= io_in_r_bypass_5_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_1_stall_8 <= io_in_r_bypass_5_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_2_data_8 <= io_in_r_bypass_5_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_2_load_store_8 <= io_in_r_bypass_5_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_2_df_is_ws_8 <= io_in_r_bypass_5_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_2_stall_8 <= io_in_r_bypass_5_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_3_data_8 <= io_in_r_bypass_5_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_3_load_store_8 <= io_in_r_bypass_5_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_3_df_is_ws_8 <= io_in_r_bypass_5_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_3_stall_8 <= io_in_r_bypass_5_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_0_data_8 <= io_in_r_bypass_6_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_0_load_store_8 <= io_in_r_bypass_6_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_0_df_is_ws_8 <= io_in_r_bypass_6_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_0_stall_8 <= io_in_r_bypass_6_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_1_data_8 <= io_in_r_bypass_6_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_1_load_store_8 <= io_in_r_bypass_6_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_1_df_is_ws_8 <= io_in_r_bypass_6_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_1_stall_8 <= io_in_r_bypass_6_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_2_data_8 <= io_in_r_bypass_6_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_2_load_store_8 <= io_in_r_bypass_6_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_2_df_is_ws_8 <= io_in_r_bypass_6_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_2_stall_8 <= io_in_r_bypass_6_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_3_data_8 <= io_in_r_bypass_6_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_3_load_store_8 <= io_in_r_bypass_6_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_3_df_is_ws_8 <= io_in_r_bypass_6_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_3_stall_8 <= io_in_r_bypass_6_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_0_data_8 <= io_in_r_bypass_7_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_0_load_store_8 <= io_in_r_bypass_7_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_0_df_is_ws_8 <= io_in_r_bypass_7_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_0_stall_8 <= io_in_r_bypass_7_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_1_data_8 <= io_in_r_bypass_7_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_1_load_store_8 <= io_in_r_bypass_7_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_1_df_is_ws_8 <= io_in_r_bypass_7_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_1_stall_8 <= io_in_r_bypass_7_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_2_data_8 <= io_in_r_bypass_7_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_2_load_store_8 <= io_in_r_bypass_7_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_2_df_is_ws_8 <= io_in_r_bypass_7_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_2_stall_8 <= io_in_r_bypass_7_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_3_data_8 <= io_in_r_bypass_7_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_3_load_store_8 <= io_in_r_bypass_7_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_3_df_is_ws_8 <= io_in_r_bypass_7_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_3_stall_8 <= io_in_r_bypass_7_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_0_data_8 <= io_in_r_bypass_8_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_0_load_store_8 <= io_in_r_bypass_8_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_0_df_is_ws_8 <= io_in_r_bypass_8_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_0_stall_8 <= io_in_r_bypass_8_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_1_data_8 <= io_in_r_bypass_8_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_1_load_store_8 <= io_in_r_bypass_8_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_1_df_is_ws_8 <= io_in_r_bypass_8_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_1_stall_8 <= io_in_r_bypass_8_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_2_data_8 <= io_in_r_bypass_8_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_2_load_store_8 <= io_in_r_bypass_8_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_2_df_is_ws_8 <= io_in_r_bypass_8_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_2_stall_8 <= io_in_r_bypass_8_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_3_data_8 <= io_in_r_bypass_8_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_3_load_store_8 <= io_in_r_bypass_8_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_3_df_is_ws_8 <= io_in_r_bypass_8_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_3_stall_8 <= io_in_r_bypass_8_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_0_data_8 <= io_in_r_bypass_9_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_0_load_store_8 <= io_in_r_bypass_9_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_0_df_is_ws_8 <= io_in_r_bypass_9_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_0_stall_8 <= io_in_r_bypass_9_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_1_data_8 <= io_in_r_bypass_9_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_1_load_store_8 <= io_in_r_bypass_9_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_1_df_is_ws_8 <= io_in_r_bypass_9_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_1_stall_8 <= io_in_r_bypass_9_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_2_data_8 <= io_in_r_bypass_9_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_2_load_store_8 <= io_in_r_bypass_9_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_2_df_is_ws_8 <= io_in_r_bypass_9_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_2_stall_8 <= io_in_r_bypass_9_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_3_data_8 <= io_in_r_bypass_9_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_3_load_store_8 <= io_in_r_bypass_9_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_3_df_is_ws_8 <= io_in_r_bypass_9_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_3_stall_8 <= io_in_r_bypass_9_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_0_data_8 <= io_in_r_bypass_10_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_0_load_store_8 <= io_in_r_bypass_10_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_0_df_is_ws_8 <= io_in_r_bypass_10_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_0_stall_8 <= io_in_r_bypass_10_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_1_data_8 <= io_in_r_bypass_10_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_1_load_store_8 <= io_in_r_bypass_10_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_1_df_is_ws_8 <= io_in_r_bypass_10_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_1_stall_8 <= io_in_r_bypass_10_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_2_data_8 <= io_in_r_bypass_10_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_2_load_store_8 <= io_in_r_bypass_10_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_2_df_is_ws_8 <= io_in_r_bypass_10_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_2_stall_8 <= io_in_r_bypass_10_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_3_data_8 <= io_in_r_bypass_10_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_3_load_store_8 <= io_in_r_bypass_10_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_3_df_is_ws_8 <= io_in_r_bypass_10_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_3_stall_8 <= io_in_r_bypass_10_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_0_data_8 <= io_in_r_bypass_11_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_0_load_store_8 <= io_in_r_bypass_11_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_0_df_is_ws_8 <= io_in_r_bypass_11_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_0_stall_8 <= io_in_r_bypass_11_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_1_data_8 <= io_in_r_bypass_11_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_1_load_store_8 <= io_in_r_bypass_11_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_1_df_is_ws_8 <= io_in_r_bypass_11_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_1_stall_8 <= io_in_r_bypass_11_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_2_data_8 <= io_in_r_bypass_11_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_2_load_store_8 <= io_in_r_bypass_11_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_2_df_is_ws_8 <= io_in_r_bypass_11_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_2_stall_8 <= io_in_r_bypass_11_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_3_data_8 <= io_in_r_bypass_11_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_3_load_store_8 <= io_in_r_bypass_11_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_3_df_is_ws_8 <= io_in_r_bypass_11_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_3_stall_8 <= io_in_r_bypass_11_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_0_data_8 <= io_in_r_bypass_12_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_0_load_store_8 <= io_in_r_bypass_12_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_0_df_is_ws_8 <= io_in_r_bypass_12_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_0_stall_8 <= io_in_r_bypass_12_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_1_data_8 <= io_in_r_bypass_12_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_1_load_store_8 <= io_in_r_bypass_12_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_1_df_is_ws_8 <= io_in_r_bypass_12_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_1_stall_8 <= io_in_r_bypass_12_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_2_data_8 <= io_in_r_bypass_12_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_2_load_store_8 <= io_in_r_bypass_12_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_2_df_is_ws_8 <= io_in_r_bypass_12_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_2_stall_8 <= io_in_r_bypass_12_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_3_data_8 <= io_in_r_bypass_12_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_3_load_store_8 <= io_in_r_bypass_12_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_3_df_is_ws_8 <= io_in_r_bypass_12_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_3_stall_8 <= io_in_r_bypass_12_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_0_data_8 <= io_in_r_bypass_13_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_0_load_store_8 <= io_in_r_bypass_13_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_0_df_is_ws_8 <= io_in_r_bypass_13_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_0_stall_8 <= io_in_r_bypass_13_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_1_data_8 <= io_in_r_bypass_13_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_1_load_store_8 <= io_in_r_bypass_13_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_1_df_is_ws_8 <= io_in_r_bypass_13_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_1_stall_8 <= io_in_r_bypass_13_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_2_data_8 <= io_in_r_bypass_13_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_2_load_store_8 <= io_in_r_bypass_13_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_2_df_is_ws_8 <= io_in_r_bypass_13_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_2_stall_8 <= io_in_r_bypass_13_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_3_data_8 <= io_in_r_bypass_13_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_3_load_store_8 <= io_in_r_bypass_13_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_3_df_is_ws_8 <= io_in_r_bypass_13_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_3_stall_8 <= io_in_r_bypass_13_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_0_data_8 <= io_in_r_bypass_14_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_0_load_store_8 <= io_in_r_bypass_14_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_0_df_is_ws_8 <= io_in_r_bypass_14_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_0_stall_8 <= io_in_r_bypass_14_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_1_data_8 <= io_in_r_bypass_14_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_1_load_store_8 <= io_in_r_bypass_14_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_1_df_is_ws_8 <= io_in_r_bypass_14_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_1_stall_8 <= io_in_r_bypass_14_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_2_data_8 <= io_in_r_bypass_14_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_2_load_store_8 <= io_in_r_bypass_14_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_2_df_is_ws_8 <= io_in_r_bypass_14_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_2_stall_8 <= io_in_r_bypass_14_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_3_data_8 <= io_in_r_bypass_14_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_3_load_store_8 <= io_in_r_bypass_14_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_3_df_is_ws_8 <= io_in_r_bypass_14_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_3_stall_8 <= io_in_r_bypass_14_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_0_data_8 <= io_in_r_bypass_15_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_0_load_store_8 <= io_in_r_bypass_15_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_0_df_is_ws_8 <= io_in_r_bypass_15_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_0_stall_8 <= io_in_r_bypass_15_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_1_data_8 <= io_in_r_bypass_15_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_1_load_store_8 <= io_in_r_bypass_15_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_1_df_is_ws_8 <= io_in_r_bypass_15_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_1_stall_8 <= io_in_r_bypass_15_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_2_data_8 <= io_in_r_bypass_15_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_2_load_store_8 <= io_in_r_bypass_15_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_2_df_is_ws_8 <= io_in_r_bypass_15_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_2_stall_8 <= io_in_r_bypass_15_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_3_data_8 <= io_in_r_bypass_15_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_3_load_store_8 <= io_in_r_bypass_15_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_3_df_is_ws_8 <= io_in_r_bypass_15_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_3_stall_8 <= io_in_r_bypass_15_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_0_data_8 <= io_in_r_bypass_16_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_0_load_store_8 <= io_in_r_bypass_16_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_0_df_is_ws_8 <= io_in_r_bypass_16_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_0_stall_8 <= io_in_r_bypass_16_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_1_data_8 <= io_in_r_bypass_16_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_1_load_store_8 <= io_in_r_bypass_16_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_1_df_is_ws_8 <= io_in_r_bypass_16_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_1_stall_8 <= io_in_r_bypass_16_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_2_data_8 <= io_in_r_bypass_16_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_2_load_store_8 <= io_in_r_bypass_16_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_2_df_is_ws_8 <= io_in_r_bypass_16_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_2_stall_8 <= io_in_r_bypass_16_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_3_data_8 <= io_in_r_bypass_16_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_3_load_store_8 <= io_in_r_bypass_16_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_3_df_is_ws_8 <= io_in_r_bypass_16_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_3_stall_8 <= io_in_r_bypass_16_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_0_data_8 <= io_in_r_bypass_17_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_0_load_store_8 <= io_in_r_bypass_17_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_0_df_is_ws_8 <= io_in_r_bypass_17_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_0_stall_8 <= io_in_r_bypass_17_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_1_data_8 <= io_in_r_bypass_17_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_1_load_store_8 <= io_in_r_bypass_17_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_1_df_is_ws_8 <= io_in_r_bypass_17_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_1_stall_8 <= io_in_r_bypass_17_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_2_data_8 <= io_in_r_bypass_17_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_2_load_store_8 <= io_in_r_bypass_17_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_2_df_is_ws_8 <= io_in_r_bypass_17_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_2_stall_8 <= io_in_r_bypass_17_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_3_data_8 <= io_in_r_bypass_17_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_3_load_store_8 <= io_in_r_bypass_17_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_3_df_is_ws_8 <= io_in_r_bypass_17_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_3_stall_8 <= io_in_r_bypass_17_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_0_data_8 <= io_in_r_bypass_18_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_0_load_store_8 <= io_in_r_bypass_18_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_0_df_is_ws_8 <= io_in_r_bypass_18_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_0_stall_8 <= io_in_r_bypass_18_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_1_data_8 <= io_in_r_bypass_18_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_1_load_store_8 <= io_in_r_bypass_18_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_1_df_is_ws_8 <= io_in_r_bypass_18_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_1_stall_8 <= io_in_r_bypass_18_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_2_data_8 <= io_in_r_bypass_18_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_2_load_store_8 <= io_in_r_bypass_18_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_2_df_is_ws_8 <= io_in_r_bypass_18_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_2_stall_8 <= io_in_r_bypass_18_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_3_data_8 <= io_in_r_bypass_18_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_3_load_store_8 <= io_in_r_bypass_18_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_3_df_is_ws_8 <= io_in_r_bypass_18_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_3_stall_8 <= io_in_r_bypass_18_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_0_data_8 <= io_in_r_bypass_19_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_0_load_store_8 <= io_in_r_bypass_19_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_0_df_is_ws_8 <= io_in_r_bypass_19_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_0_stall_8 <= io_in_r_bypass_19_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_1_data_8 <= io_in_r_bypass_19_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_1_load_store_8 <= io_in_r_bypass_19_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_1_df_is_ws_8 <= io_in_r_bypass_19_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_1_stall_8 <= io_in_r_bypass_19_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_2_data_8 <= io_in_r_bypass_19_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_2_load_store_8 <= io_in_r_bypass_19_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_2_df_is_ws_8 <= io_in_r_bypass_19_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_2_stall_8 <= io_in_r_bypass_19_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_3_data_8 <= io_in_r_bypass_19_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_3_load_store_8 <= io_in_r_bypass_19_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_3_df_is_ws_8 <= io_in_r_bypass_19_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_3_stall_8 <= io_in_r_bypass_19_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_0_data_8 <= io_in_r_bypass_20_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_0_load_store_8 <= io_in_r_bypass_20_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_0_df_is_ws_8 <= io_in_r_bypass_20_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_0_stall_8 <= io_in_r_bypass_20_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_1_data_8 <= io_in_r_bypass_20_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_1_load_store_8 <= io_in_r_bypass_20_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_1_df_is_ws_8 <= io_in_r_bypass_20_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_1_stall_8 <= io_in_r_bypass_20_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_2_data_8 <= io_in_r_bypass_20_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_2_load_store_8 <= io_in_r_bypass_20_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_2_df_is_ws_8 <= io_in_r_bypass_20_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_2_stall_8 <= io_in_r_bypass_20_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_3_data_8 <= io_in_r_bypass_20_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_3_load_store_8 <= io_in_r_bypass_20_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_3_df_is_ws_8 <= io_in_r_bypass_20_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_3_stall_8 <= io_in_r_bypass_20_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_0_data_8 <= io_in_r_bypass_21_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_0_load_store_8 <= io_in_r_bypass_21_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_0_df_is_ws_8 <= io_in_r_bypass_21_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_0_stall_8 <= io_in_r_bypass_21_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_1_data_8 <= io_in_r_bypass_21_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_1_load_store_8 <= io_in_r_bypass_21_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_1_df_is_ws_8 <= io_in_r_bypass_21_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_1_stall_8 <= io_in_r_bypass_21_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_2_data_8 <= io_in_r_bypass_21_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_2_load_store_8 <= io_in_r_bypass_21_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_2_df_is_ws_8 <= io_in_r_bypass_21_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_2_stall_8 <= io_in_r_bypass_21_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_3_data_8 <= io_in_r_bypass_21_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_3_load_store_8 <= io_in_r_bypass_21_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_3_df_is_ws_8 <= io_in_r_bypass_21_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_3_stall_8 <= io_in_r_bypass_21_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_0_data_8 <= io_in_r_bypass_22_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_0_load_store_8 <= io_in_r_bypass_22_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_0_df_is_ws_8 <= io_in_r_bypass_22_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_0_stall_8 <= io_in_r_bypass_22_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_1_data_8 <= io_in_r_bypass_22_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_1_load_store_8 <= io_in_r_bypass_22_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_1_df_is_ws_8 <= io_in_r_bypass_22_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_1_stall_8 <= io_in_r_bypass_22_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_2_data_8 <= io_in_r_bypass_22_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_2_load_store_8 <= io_in_r_bypass_22_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_2_df_is_ws_8 <= io_in_r_bypass_22_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_2_stall_8 <= io_in_r_bypass_22_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_3_data_8 <= io_in_r_bypass_22_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_3_load_store_8 <= io_in_r_bypass_22_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_3_df_is_ws_8 <= io_in_r_bypass_22_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_3_stall_8 <= io_in_r_bypass_22_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_0_data_8 <= io_in_r_bypass_23_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_0_load_store_8 <= io_in_r_bypass_23_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_0_df_is_ws_8 <= io_in_r_bypass_23_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_0_stall_8 <= io_in_r_bypass_23_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_1_data_8 <= io_in_r_bypass_23_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_1_load_store_8 <= io_in_r_bypass_23_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_1_df_is_ws_8 <= io_in_r_bypass_23_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_1_stall_8 <= io_in_r_bypass_23_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_2_data_8 <= io_in_r_bypass_23_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_2_load_store_8 <= io_in_r_bypass_23_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_2_df_is_ws_8 <= io_in_r_bypass_23_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_2_stall_8 <= io_in_r_bypass_23_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_3_data_8 <= io_in_r_bypass_23_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_3_load_store_8 <= io_in_r_bypass_23_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_3_df_is_ws_8 <= io_in_r_bypass_23_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_3_stall_8 <= io_in_r_bypass_23_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_0_data_8 <= io_in_r_bypass_24_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_0_load_store_8 <= io_in_r_bypass_24_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_0_df_is_ws_8 <= io_in_r_bypass_24_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_0_stall_8 <= io_in_r_bypass_24_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_1_data_8 <= io_in_r_bypass_24_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_1_load_store_8 <= io_in_r_bypass_24_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_1_df_is_ws_8 <= io_in_r_bypass_24_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_1_stall_8 <= io_in_r_bypass_24_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_2_data_8 <= io_in_r_bypass_24_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_2_load_store_8 <= io_in_r_bypass_24_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_2_df_is_ws_8 <= io_in_r_bypass_24_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_2_stall_8 <= io_in_r_bypass_24_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_3_data_8 <= io_in_r_bypass_24_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_3_load_store_8 <= io_in_r_bypass_24_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_3_df_is_ws_8 <= io_in_r_bypass_24_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_3_stall_8 <= io_in_r_bypass_24_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_0_data_8 <= io_in_r_bypass_25_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_0_load_store_8 <= io_in_r_bypass_25_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_0_df_is_ws_8 <= io_in_r_bypass_25_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_0_stall_8 <= io_in_r_bypass_25_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_1_data_8 <= io_in_r_bypass_25_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_1_load_store_8 <= io_in_r_bypass_25_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_1_df_is_ws_8 <= io_in_r_bypass_25_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_1_stall_8 <= io_in_r_bypass_25_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_2_data_8 <= io_in_r_bypass_25_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_2_load_store_8 <= io_in_r_bypass_25_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_2_df_is_ws_8 <= io_in_r_bypass_25_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_2_stall_8 <= io_in_r_bypass_25_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_3_data_8 <= io_in_r_bypass_25_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_3_load_store_8 <= io_in_r_bypass_25_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_3_df_is_ws_8 <= io_in_r_bypass_25_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_3_stall_8 <= io_in_r_bypass_25_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_0_data_8 <= io_in_r_bypass_26_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_0_load_store_8 <= io_in_r_bypass_26_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_0_df_is_ws_8 <= io_in_r_bypass_26_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_0_stall_8 <= io_in_r_bypass_26_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_1_data_8 <= io_in_r_bypass_26_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_1_load_store_8 <= io_in_r_bypass_26_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_1_df_is_ws_8 <= io_in_r_bypass_26_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_1_stall_8 <= io_in_r_bypass_26_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_2_data_8 <= io_in_r_bypass_26_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_2_load_store_8 <= io_in_r_bypass_26_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_2_df_is_ws_8 <= io_in_r_bypass_26_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_2_stall_8 <= io_in_r_bypass_26_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_3_data_8 <= io_in_r_bypass_26_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_3_load_store_8 <= io_in_r_bypass_26_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_3_df_is_ws_8 <= io_in_r_bypass_26_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_3_stall_8 <= io_in_r_bypass_26_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_0_data_8 <= io_in_r_bypass_27_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_0_load_store_8 <= io_in_r_bypass_27_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_0_df_is_ws_8 <= io_in_r_bypass_27_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_0_stall_8 <= io_in_r_bypass_27_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_1_data_8 <= io_in_r_bypass_27_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_1_load_store_8 <= io_in_r_bypass_27_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_1_df_is_ws_8 <= io_in_r_bypass_27_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_1_stall_8 <= io_in_r_bypass_27_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_2_data_8 <= io_in_r_bypass_27_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_2_load_store_8 <= io_in_r_bypass_27_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_2_df_is_ws_8 <= io_in_r_bypass_27_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_2_stall_8 <= io_in_r_bypass_27_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_3_data_8 <= io_in_r_bypass_27_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_3_load_store_8 <= io_in_r_bypass_27_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_3_df_is_ws_8 <= io_in_r_bypass_27_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_3_stall_8 <= io_in_r_bypass_27_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_0_data_8 <= io_in_r_bypass_28_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_0_load_store_8 <= io_in_r_bypass_28_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_0_df_is_ws_8 <= io_in_r_bypass_28_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_0_stall_8 <= io_in_r_bypass_28_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_1_data_8 <= io_in_r_bypass_28_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_1_load_store_8 <= io_in_r_bypass_28_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_1_df_is_ws_8 <= io_in_r_bypass_28_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_1_stall_8 <= io_in_r_bypass_28_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_2_data_8 <= io_in_r_bypass_28_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_2_load_store_8 <= io_in_r_bypass_28_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_2_df_is_ws_8 <= io_in_r_bypass_28_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_2_stall_8 <= io_in_r_bypass_28_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_3_data_8 <= io_in_r_bypass_28_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_3_load_store_8 <= io_in_r_bypass_28_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_3_df_is_ws_8 <= io_in_r_bypass_28_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_3_stall_8 <= io_in_r_bypass_28_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_0_data_8 <= io_in_r_bypass_29_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_0_load_store_8 <= io_in_r_bypass_29_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_0_df_is_ws_8 <= io_in_r_bypass_29_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_0_stall_8 <= io_in_r_bypass_29_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_1_data_8 <= io_in_r_bypass_29_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_1_load_store_8 <= io_in_r_bypass_29_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_1_df_is_ws_8 <= io_in_r_bypass_29_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_1_stall_8 <= io_in_r_bypass_29_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_2_data_8 <= io_in_r_bypass_29_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_2_load_store_8 <= io_in_r_bypass_29_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_2_df_is_ws_8 <= io_in_r_bypass_29_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_2_stall_8 <= io_in_r_bypass_29_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_3_data_8 <= io_in_r_bypass_29_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_3_load_store_8 <= io_in_r_bypass_29_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_3_df_is_ws_8 <= io_in_r_bypass_29_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_3_stall_8 <= io_in_r_bypass_29_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_0_data_8 <= io_in_r_bypass_30_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_0_load_store_8 <= io_in_r_bypass_30_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_0_df_is_ws_8 <= io_in_r_bypass_30_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_0_stall_8 <= io_in_r_bypass_30_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_1_data_8 <= io_in_r_bypass_30_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_1_load_store_8 <= io_in_r_bypass_30_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_1_df_is_ws_8 <= io_in_r_bypass_30_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_1_stall_8 <= io_in_r_bypass_30_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_2_data_8 <= io_in_r_bypass_30_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_2_load_store_8 <= io_in_r_bypass_30_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_2_df_is_ws_8 <= io_in_r_bypass_30_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_2_stall_8 <= io_in_r_bypass_30_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_3_data_8 <= io_in_r_bypass_30_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_3_load_store_8 <= io_in_r_bypass_30_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_3_df_is_ws_8 <= io_in_r_bypass_30_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_3_stall_8 <= io_in_r_bypass_30_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_0_data_8 <= io_in_r_bypass_31_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_0_load_store_8 <= io_in_r_bypass_31_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_0_df_is_ws_8 <= io_in_r_bypass_31_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_0_stall_8 <= io_in_r_bypass_31_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_1_data_8 <= io_in_r_bypass_31_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_1_load_store_8 <= io_in_r_bypass_31_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_1_df_is_ws_8 <= io_in_r_bypass_31_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_1_stall_8 <= io_in_r_bypass_31_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_2_data_8 <= io_in_r_bypass_31_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_2_load_store_8 <= io_in_r_bypass_31_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_2_df_is_ws_8 <= io_in_r_bypass_31_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_2_stall_8 <= io_in_r_bypass_31_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_3_data_8 <= io_in_r_bypass_31_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_3_load_store_8 <= io_in_r_bypass_31_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_3_df_is_ws_8 <= io_in_r_bypass_31_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_3_stall_8 <= io_in_r_bypass_31_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_0_data_9 <= io_in_r_bypass_0_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_0_load_store_9 <= io_in_r_bypass_0_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_0_df_is_ws_9 <= io_in_r_bypass_0_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_0_stall_9 <= io_in_r_bypass_0_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_1_data_9 <= io_in_r_bypass_0_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_1_load_store_9 <= io_in_r_bypass_0_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_1_df_is_ws_9 <= io_in_r_bypass_0_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_1_stall_9 <= io_in_r_bypass_0_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_2_data_9 <= io_in_r_bypass_0_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_2_load_store_9 <= io_in_r_bypass_0_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_2_df_is_ws_9 <= io_in_r_bypass_0_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_2_stall_9 <= io_in_r_bypass_0_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_3_data_9 <= io_in_r_bypass_0_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_3_load_store_9 <= io_in_r_bypass_0_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_3_df_is_ws_9 <= io_in_r_bypass_0_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_3_stall_9 <= io_in_r_bypass_0_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_0_data_9 <= io_in_r_bypass_1_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_0_load_store_9 <= io_in_r_bypass_1_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_0_df_is_ws_9 <= io_in_r_bypass_1_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_0_stall_9 <= io_in_r_bypass_1_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_1_data_9 <= io_in_r_bypass_1_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_1_load_store_9 <= io_in_r_bypass_1_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_1_df_is_ws_9 <= io_in_r_bypass_1_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_1_stall_9 <= io_in_r_bypass_1_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_2_data_9 <= io_in_r_bypass_1_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_2_load_store_9 <= io_in_r_bypass_1_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_2_df_is_ws_9 <= io_in_r_bypass_1_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_2_stall_9 <= io_in_r_bypass_1_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_3_data_9 <= io_in_r_bypass_1_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_3_load_store_9 <= io_in_r_bypass_1_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_3_df_is_ws_9 <= io_in_r_bypass_1_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_3_stall_9 <= io_in_r_bypass_1_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_0_data_9 <= io_in_r_bypass_2_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_0_load_store_9 <= io_in_r_bypass_2_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_0_df_is_ws_9 <= io_in_r_bypass_2_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_0_stall_9 <= io_in_r_bypass_2_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_1_data_9 <= io_in_r_bypass_2_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_1_load_store_9 <= io_in_r_bypass_2_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_1_df_is_ws_9 <= io_in_r_bypass_2_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_1_stall_9 <= io_in_r_bypass_2_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_2_data_9 <= io_in_r_bypass_2_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_2_load_store_9 <= io_in_r_bypass_2_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_2_df_is_ws_9 <= io_in_r_bypass_2_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_2_stall_9 <= io_in_r_bypass_2_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_3_data_9 <= io_in_r_bypass_2_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_3_load_store_9 <= io_in_r_bypass_2_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_3_df_is_ws_9 <= io_in_r_bypass_2_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_3_stall_9 <= io_in_r_bypass_2_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_0_data_9 <= io_in_r_bypass_3_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_0_load_store_9 <= io_in_r_bypass_3_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_0_df_is_ws_9 <= io_in_r_bypass_3_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_0_stall_9 <= io_in_r_bypass_3_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_1_data_9 <= io_in_r_bypass_3_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_1_load_store_9 <= io_in_r_bypass_3_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_1_df_is_ws_9 <= io_in_r_bypass_3_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_1_stall_9 <= io_in_r_bypass_3_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_2_data_9 <= io_in_r_bypass_3_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_2_load_store_9 <= io_in_r_bypass_3_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_2_df_is_ws_9 <= io_in_r_bypass_3_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_2_stall_9 <= io_in_r_bypass_3_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_3_data_9 <= io_in_r_bypass_3_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_3_load_store_9 <= io_in_r_bypass_3_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_3_df_is_ws_9 <= io_in_r_bypass_3_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_3_stall_9 <= io_in_r_bypass_3_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_0_data_9 <= io_in_r_bypass_4_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_0_load_store_9 <= io_in_r_bypass_4_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_0_df_is_ws_9 <= io_in_r_bypass_4_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_0_stall_9 <= io_in_r_bypass_4_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_1_data_9 <= io_in_r_bypass_4_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_1_load_store_9 <= io_in_r_bypass_4_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_1_df_is_ws_9 <= io_in_r_bypass_4_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_1_stall_9 <= io_in_r_bypass_4_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_2_data_9 <= io_in_r_bypass_4_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_2_load_store_9 <= io_in_r_bypass_4_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_2_df_is_ws_9 <= io_in_r_bypass_4_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_2_stall_9 <= io_in_r_bypass_4_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_3_data_9 <= io_in_r_bypass_4_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_3_load_store_9 <= io_in_r_bypass_4_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_3_df_is_ws_9 <= io_in_r_bypass_4_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_3_stall_9 <= io_in_r_bypass_4_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_0_data_9 <= io_in_r_bypass_5_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_0_load_store_9 <= io_in_r_bypass_5_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_0_df_is_ws_9 <= io_in_r_bypass_5_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_0_stall_9 <= io_in_r_bypass_5_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_1_data_9 <= io_in_r_bypass_5_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_1_load_store_9 <= io_in_r_bypass_5_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_1_df_is_ws_9 <= io_in_r_bypass_5_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_1_stall_9 <= io_in_r_bypass_5_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_2_data_9 <= io_in_r_bypass_5_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_2_load_store_9 <= io_in_r_bypass_5_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_2_df_is_ws_9 <= io_in_r_bypass_5_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_2_stall_9 <= io_in_r_bypass_5_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_3_data_9 <= io_in_r_bypass_5_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_3_load_store_9 <= io_in_r_bypass_5_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_3_df_is_ws_9 <= io_in_r_bypass_5_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_3_stall_9 <= io_in_r_bypass_5_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_0_data_9 <= io_in_r_bypass_6_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_0_load_store_9 <= io_in_r_bypass_6_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_0_df_is_ws_9 <= io_in_r_bypass_6_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_0_stall_9 <= io_in_r_bypass_6_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_1_data_9 <= io_in_r_bypass_6_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_1_load_store_9 <= io_in_r_bypass_6_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_1_df_is_ws_9 <= io_in_r_bypass_6_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_1_stall_9 <= io_in_r_bypass_6_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_2_data_9 <= io_in_r_bypass_6_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_2_load_store_9 <= io_in_r_bypass_6_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_2_df_is_ws_9 <= io_in_r_bypass_6_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_2_stall_9 <= io_in_r_bypass_6_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_3_data_9 <= io_in_r_bypass_6_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_3_load_store_9 <= io_in_r_bypass_6_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_3_df_is_ws_9 <= io_in_r_bypass_6_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_3_stall_9 <= io_in_r_bypass_6_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_0_data_9 <= io_in_r_bypass_7_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_0_load_store_9 <= io_in_r_bypass_7_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_0_df_is_ws_9 <= io_in_r_bypass_7_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_0_stall_9 <= io_in_r_bypass_7_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_1_data_9 <= io_in_r_bypass_7_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_1_load_store_9 <= io_in_r_bypass_7_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_1_df_is_ws_9 <= io_in_r_bypass_7_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_1_stall_9 <= io_in_r_bypass_7_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_2_data_9 <= io_in_r_bypass_7_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_2_load_store_9 <= io_in_r_bypass_7_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_2_df_is_ws_9 <= io_in_r_bypass_7_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_2_stall_9 <= io_in_r_bypass_7_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_3_data_9 <= io_in_r_bypass_7_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_3_load_store_9 <= io_in_r_bypass_7_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_3_df_is_ws_9 <= io_in_r_bypass_7_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_3_stall_9 <= io_in_r_bypass_7_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_0_data_9 <= io_in_r_bypass_8_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_0_load_store_9 <= io_in_r_bypass_8_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_0_df_is_ws_9 <= io_in_r_bypass_8_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_0_stall_9 <= io_in_r_bypass_8_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_1_data_9 <= io_in_r_bypass_8_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_1_load_store_9 <= io_in_r_bypass_8_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_1_df_is_ws_9 <= io_in_r_bypass_8_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_1_stall_9 <= io_in_r_bypass_8_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_2_data_9 <= io_in_r_bypass_8_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_2_load_store_9 <= io_in_r_bypass_8_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_2_df_is_ws_9 <= io_in_r_bypass_8_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_2_stall_9 <= io_in_r_bypass_8_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_3_data_9 <= io_in_r_bypass_8_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_3_load_store_9 <= io_in_r_bypass_8_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_3_df_is_ws_9 <= io_in_r_bypass_8_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_3_stall_9 <= io_in_r_bypass_8_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_0_data_9 <= io_in_r_bypass_9_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_0_load_store_9 <= io_in_r_bypass_9_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_0_df_is_ws_9 <= io_in_r_bypass_9_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_0_stall_9 <= io_in_r_bypass_9_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_1_data_9 <= io_in_r_bypass_9_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_1_load_store_9 <= io_in_r_bypass_9_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_1_df_is_ws_9 <= io_in_r_bypass_9_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_1_stall_9 <= io_in_r_bypass_9_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_2_data_9 <= io_in_r_bypass_9_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_2_load_store_9 <= io_in_r_bypass_9_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_2_df_is_ws_9 <= io_in_r_bypass_9_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_2_stall_9 <= io_in_r_bypass_9_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_3_data_9 <= io_in_r_bypass_9_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_3_load_store_9 <= io_in_r_bypass_9_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_3_df_is_ws_9 <= io_in_r_bypass_9_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_3_stall_9 <= io_in_r_bypass_9_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_0_data_9 <= io_in_r_bypass_10_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_0_load_store_9 <= io_in_r_bypass_10_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_0_df_is_ws_9 <= io_in_r_bypass_10_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_0_stall_9 <= io_in_r_bypass_10_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_1_data_9 <= io_in_r_bypass_10_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_1_load_store_9 <= io_in_r_bypass_10_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_1_df_is_ws_9 <= io_in_r_bypass_10_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_1_stall_9 <= io_in_r_bypass_10_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_2_data_9 <= io_in_r_bypass_10_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_2_load_store_9 <= io_in_r_bypass_10_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_2_df_is_ws_9 <= io_in_r_bypass_10_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_2_stall_9 <= io_in_r_bypass_10_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_3_data_9 <= io_in_r_bypass_10_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_3_load_store_9 <= io_in_r_bypass_10_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_3_df_is_ws_9 <= io_in_r_bypass_10_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_3_stall_9 <= io_in_r_bypass_10_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_0_data_9 <= io_in_r_bypass_11_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_0_load_store_9 <= io_in_r_bypass_11_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_0_df_is_ws_9 <= io_in_r_bypass_11_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_0_stall_9 <= io_in_r_bypass_11_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_1_data_9 <= io_in_r_bypass_11_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_1_load_store_9 <= io_in_r_bypass_11_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_1_df_is_ws_9 <= io_in_r_bypass_11_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_1_stall_9 <= io_in_r_bypass_11_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_2_data_9 <= io_in_r_bypass_11_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_2_load_store_9 <= io_in_r_bypass_11_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_2_df_is_ws_9 <= io_in_r_bypass_11_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_2_stall_9 <= io_in_r_bypass_11_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_3_data_9 <= io_in_r_bypass_11_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_3_load_store_9 <= io_in_r_bypass_11_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_3_df_is_ws_9 <= io_in_r_bypass_11_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_3_stall_9 <= io_in_r_bypass_11_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_0_data_9 <= io_in_r_bypass_12_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_0_load_store_9 <= io_in_r_bypass_12_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_0_df_is_ws_9 <= io_in_r_bypass_12_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_0_stall_9 <= io_in_r_bypass_12_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_1_data_9 <= io_in_r_bypass_12_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_1_load_store_9 <= io_in_r_bypass_12_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_1_df_is_ws_9 <= io_in_r_bypass_12_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_1_stall_9 <= io_in_r_bypass_12_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_2_data_9 <= io_in_r_bypass_12_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_2_load_store_9 <= io_in_r_bypass_12_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_2_df_is_ws_9 <= io_in_r_bypass_12_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_2_stall_9 <= io_in_r_bypass_12_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_3_data_9 <= io_in_r_bypass_12_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_3_load_store_9 <= io_in_r_bypass_12_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_3_df_is_ws_9 <= io_in_r_bypass_12_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_3_stall_9 <= io_in_r_bypass_12_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_0_data_9 <= io_in_r_bypass_13_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_0_load_store_9 <= io_in_r_bypass_13_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_0_df_is_ws_9 <= io_in_r_bypass_13_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_0_stall_9 <= io_in_r_bypass_13_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_1_data_9 <= io_in_r_bypass_13_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_1_load_store_9 <= io_in_r_bypass_13_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_1_df_is_ws_9 <= io_in_r_bypass_13_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_1_stall_9 <= io_in_r_bypass_13_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_2_data_9 <= io_in_r_bypass_13_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_2_load_store_9 <= io_in_r_bypass_13_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_2_df_is_ws_9 <= io_in_r_bypass_13_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_2_stall_9 <= io_in_r_bypass_13_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_3_data_9 <= io_in_r_bypass_13_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_3_load_store_9 <= io_in_r_bypass_13_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_3_df_is_ws_9 <= io_in_r_bypass_13_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_3_stall_9 <= io_in_r_bypass_13_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_0_data_9 <= io_in_r_bypass_14_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_0_load_store_9 <= io_in_r_bypass_14_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_0_df_is_ws_9 <= io_in_r_bypass_14_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_0_stall_9 <= io_in_r_bypass_14_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_1_data_9 <= io_in_r_bypass_14_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_1_load_store_9 <= io_in_r_bypass_14_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_1_df_is_ws_9 <= io_in_r_bypass_14_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_1_stall_9 <= io_in_r_bypass_14_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_2_data_9 <= io_in_r_bypass_14_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_2_load_store_9 <= io_in_r_bypass_14_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_2_df_is_ws_9 <= io_in_r_bypass_14_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_2_stall_9 <= io_in_r_bypass_14_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_3_data_9 <= io_in_r_bypass_14_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_3_load_store_9 <= io_in_r_bypass_14_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_3_df_is_ws_9 <= io_in_r_bypass_14_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_3_stall_9 <= io_in_r_bypass_14_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_0_data_9 <= io_in_r_bypass_15_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_0_load_store_9 <= io_in_r_bypass_15_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_0_df_is_ws_9 <= io_in_r_bypass_15_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_0_stall_9 <= io_in_r_bypass_15_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_1_data_9 <= io_in_r_bypass_15_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_1_load_store_9 <= io_in_r_bypass_15_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_1_df_is_ws_9 <= io_in_r_bypass_15_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_1_stall_9 <= io_in_r_bypass_15_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_2_data_9 <= io_in_r_bypass_15_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_2_load_store_9 <= io_in_r_bypass_15_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_2_df_is_ws_9 <= io_in_r_bypass_15_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_2_stall_9 <= io_in_r_bypass_15_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_3_data_9 <= io_in_r_bypass_15_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_3_load_store_9 <= io_in_r_bypass_15_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_3_df_is_ws_9 <= io_in_r_bypass_15_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_3_stall_9 <= io_in_r_bypass_15_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_0_data_9 <= io_in_r_bypass_16_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_0_load_store_9 <= io_in_r_bypass_16_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_0_df_is_ws_9 <= io_in_r_bypass_16_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_0_stall_9 <= io_in_r_bypass_16_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_1_data_9 <= io_in_r_bypass_16_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_1_load_store_9 <= io_in_r_bypass_16_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_1_df_is_ws_9 <= io_in_r_bypass_16_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_1_stall_9 <= io_in_r_bypass_16_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_2_data_9 <= io_in_r_bypass_16_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_2_load_store_9 <= io_in_r_bypass_16_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_2_df_is_ws_9 <= io_in_r_bypass_16_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_2_stall_9 <= io_in_r_bypass_16_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_3_data_9 <= io_in_r_bypass_16_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_3_load_store_9 <= io_in_r_bypass_16_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_3_df_is_ws_9 <= io_in_r_bypass_16_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_3_stall_9 <= io_in_r_bypass_16_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_0_data_9 <= io_in_r_bypass_17_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_0_load_store_9 <= io_in_r_bypass_17_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_0_df_is_ws_9 <= io_in_r_bypass_17_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_0_stall_9 <= io_in_r_bypass_17_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_1_data_9 <= io_in_r_bypass_17_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_1_load_store_9 <= io_in_r_bypass_17_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_1_df_is_ws_9 <= io_in_r_bypass_17_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_1_stall_9 <= io_in_r_bypass_17_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_2_data_9 <= io_in_r_bypass_17_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_2_load_store_9 <= io_in_r_bypass_17_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_2_df_is_ws_9 <= io_in_r_bypass_17_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_2_stall_9 <= io_in_r_bypass_17_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_3_data_9 <= io_in_r_bypass_17_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_3_load_store_9 <= io_in_r_bypass_17_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_3_df_is_ws_9 <= io_in_r_bypass_17_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_3_stall_9 <= io_in_r_bypass_17_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_0_data_9 <= io_in_r_bypass_18_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_0_load_store_9 <= io_in_r_bypass_18_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_0_df_is_ws_9 <= io_in_r_bypass_18_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_0_stall_9 <= io_in_r_bypass_18_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_1_data_9 <= io_in_r_bypass_18_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_1_load_store_9 <= io_in_r_bypass_18_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_1_df_is_ws_9 <= io_in_r_bypass_18_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_1_stall_9 <= io_in_r_bypass_18_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_2_data_9 <= io_in_r_bypass_18_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_2_load_store_9 <= io_in_r_bypass_18_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_2_df_is_ws_9 <= io_in_r_bypass_18_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_2_stall_9 <= io_in_r_bypass_18_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_3_data_9 <= io_in_r_bypass_18_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_3_load_store_9 <= io_in_r_bypass_18_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_3_df_is_ws_9 <= io_in_r_bypass_18_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_3_stall_9 <= io_in_r_bypass_18_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_0_data_9 <= io_in_r_bypass_19_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_0_load_store_9 <= io_in_r_bypass_19_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_0_df_is_ws_9 <= io_in_r_bypass_19_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_0_stall_9 <= io_in_r_bypass_19_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_1_data_9 <= io_in_r_bypass_19_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_1_load_store_9 <= io_in_r_bypass_19_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_1_df_is_ws_9 <= io_in_r_bypass_19_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_1_stall_9 <= io_in_r_bypass_19_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_2_data_9 <= io_in_r_bypass_19_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_2_load_store_9 <= io_in_r_bypass_19_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_2_df_is_ws_9 <= io_in_r_bypass_19_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_2_stall_9 <= io_in_r_bypass_19_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_3_data_9 <= io_in_r_bypass_19_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_3_load_store_9 <= io_in_r_bypass_19_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_3_df_is_ws_9 <= io_in_r_bypass_19_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_3_stall_9 <= io_in_r_bypass_19_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_0_data_9 <= io_in_r_bypass_20_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_0_load_store_9 <= io_in_r_bypass_20_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_0_df_is_ws_9 <= io_in_r_bypass_20_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_0_stall_9 <= io_in_r_bypass_20_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_1_data_9 <= io_in_r_bypass_20_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_1_load_store_9 <= io_in_r_bypass_20_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_1_df_is_ws_9 <= io_in_r_bypass_20_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_1_stall_9 <= io_in_r_bypass_20_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_2_data_9 <= io_in_r_bypass_20_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_2_load_store_9 <= io_in_r_bypass_20_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_2_df_is_ws_9 <= io_in_r_bypass_20_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_2_stall_9 <= io_in_r_bypass_20_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_3_data_9 <= io_in_r_bypass_20_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_3_load_store_9 <= io_in_r_bypass_20_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_3_df_is_ws_9 <= io_in_r_bypass_20_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_3_stall_9 <= io_in_r_bypass_20_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_0_data_9 <= io_in_r_bypass_21_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_0_load_store_9 <= io_in_r_bypass_21_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_0_df_is_ws_9 <= io_in_r_bypass_21_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_0_stall_9 <= io_in_r_bypass_21_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_1_data_9 <= io_in_r_bypass_21_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_1_load_store_9 <= io_in_r_bypass_21_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_1_df_is_ws_9 <= io_in_r_bypass_21_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_1_stall_9 <= io_in_r_bypass_21_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_2_data_9 <= io_in_r_bypass_21_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_2_load_store_9 <= io_in_r_bypass_21_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_2_df_is_ws_9 <= io_in_r_bypass_21_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_2_stall_9 <= io_in_r_bypass_21_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_3_data_9 <= io_in_r_bypass_21_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_3_load_store_9 <= io_in_r_bypass_21_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_3_df_is_ws_9 <= io_in_r_bypass_21_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_3_stall_9 <= io_in_r_bypass_21_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_0_data_9 <= io_in_r_bypass_22_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_0_load_store_9 <= io_in_r_bypass_22_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_0_df_is_ws_9 <= io_in_r_bypass_22_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_0_stall_9 <= io_in_r_bypass_22_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_1_data_9 <= io_in_r_bypass_22_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_1_load_store_9 <= io_in_r_bypass_22_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_1_df_is_ws_9 <= io_in_r_bypass_22_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_1_stall_9 <= io_in_r_bypass_22_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_2_data_9 <= io_in_r_bypass_22_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_2_load_store_9 <= io_in_r_bypass_22_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_2_df_is_ws_9 <= io_in_r_bypass_22_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_2_stall_9 <= io_in_r_bypass_22_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_3_data_9 <= io_in_r_bypass_22_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_3_load_store_9 <= io_in_r_bypass_22_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_3_df_is_ws_9 <= io_in_r_bypass_22_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_3_stall_9 <= io_in_r_bypass_22_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_0_data_9 <= io_in_r_bypass_23_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_0_load_store_9 <= io_in_r_bypass_23_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_0_df_is_ws_9 <= io_in_r_bypass_23_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_0_stall_9 <= io_in_r_bypass_23_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_1_data_9 <= io_in_r_bypass_23_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_1_load_store_9 <= io_in_r_bypass_23_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_1_df_is_ws_9 <= io_in_r_bypass_23_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_1_stall_9 <= io_in_r_bypass_23_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_2_data_9 <= io_in_r_bypass_23_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_2_load_store_9 <= io_in_r_bypass_23_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_2_df_is_ws_9 <= io_in_r_bypass_23_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_2_stall_9 <= io_in_r_bypass_23_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_3_data_9 <= io_in_r_bypass_23_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_3_load_store_9 <= io_in_r_bypass_23_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_3_df_is_ws_9 <= io_in_r_bypass_23_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_3_stall_9 <= io_in_r_bypass_23_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_0_data_9 <= io_in_r_bypass_24_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_0_load_store_9 <= io_in_r_bypass_24_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_0_df_is_ws_9 <= io_in_r_bypass_24_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_0_stall_9 <= io_in_r_bypass_24_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_1_data_9 <= io_in_r_bypass_24_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_1_load_store_9 <= io_in_r_bypass_24_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_1_df_is_ws_9 <= io_in_r_bypass_24_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_1_stall_9 <= io_in_r_bypass_24_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_2_data_9 <= io_in_r_bypass_24_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_2_load_store_9 <= io_in_r_bypass_24_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_2_df_is_ws_9 <= io_in_r_bypass_24_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_2_stall_9 <= io_in_r_bypass_24_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_3_data_9 <= io_in_r_bypass_24_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_3_load_store_9 <= io_in_r_bypass_24_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_3_df_is_ws_9 <= io_in_r_bypass_24_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_3_stall_9 <= io_in_r_bypass_24_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_0_data_9 <= io_in_r_bypass_25_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_0_load_store_9 <= io_in_r_bypass_25_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_0_df_is_ws_9 <= io_in_r_bypass_25_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_0_stall_9 <= io_in_r_bypass_25_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_1_data_9 <= io_in_r_bypass_25_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_1_load_store_9 <= io_in_r_bypass_25_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_1_df_is_ws_9 <= io_in_r_bypass_25_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_1_stall_9 <= io_in_r_bypass_25_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_2_data_9 <= io_in_r_bypass_25_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_2_load_store_9 <= io_in_r_bypass_25_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_2_df_is_ws_9 <= io_in_r_bypass_25_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_2_stall_9 <= io_in_r_bypass_25_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_3_data_9 <= io_in_r_bypass_25_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_3_load_store_9 <= io_in_r_bypass_25_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_3_df_is_ws_9 <= io_in_r_bypass_25_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_3_stall_9 <= io_in_r_bypass_25_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_0_data_9 <= io_in_r_bypass_26_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_0_load_store_9 <= io_in_r_bypass_26_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_0_df_is_ws_9 <= io_in_r_bypass_26_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_0_stall_9 <= io_in_r_bypass_26_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_1_data_9 <= io_in_r_bypass_26_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_1_load_store_9 <= io_in_r_bypass_26_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_1_df_is_ws_9 <= io_in_r_bypass_26_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_1_stall_9 <= io_in_r_bypass_26_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_2_data_9 <= io_in_r_bypass_26_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_2_load_store_9 <= io_in_r_bypass_26_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_2_df_is_ws_9 <= io_in_r_bypass_26_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_2_stall_9 <= io_in_r_bypass_26_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_3_data_9 <= io_in_r_bypass_26_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_3_load_store_9 <= io_in_r_bypass_26_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_3_df_is_ws_9 <= io_in_r_bypass_26_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_3_stall_9 <= io_in_r_bypass_26_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_0_data_9 <= io_in_r_bypass_27_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_0_load_store_9 <= io_in_r_bypass_27_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_0_df_is_ws_9 <= io_in_r_bypass_27_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_0_stall_9 <= io_in_r_bypass_27_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_1_data_9 <= io_in_r_bypass_27_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_1_load_store_9 <= io_in_r_bypass_27_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_1_df_is_ws_9 <= io_in_r_bypass_27_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_1_stall_9 <= io_in_r_bypass_27_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_2_data_9 <= io_in_r_bypass_27_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_2_load_store_9 <= io_in_r_bypass_27_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_2_df_is_ws_9 <= io_in_r_bypass_27_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_2_stall_9 <= io_in_r_bypass_27_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_3_data_9 <= io_in_r_bypass_27_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_3_load_store_9 <= io_in_r_bypass_27_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_3_df_is_ws_9 <= io_in_r_bypass_27_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_3_stall_9 <= io_in_r_bypass_27_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_0_data_9 <= io_in_r_bypass_28_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_0_load_store_9 <= io_in_r_bypass_28_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_0_df_is_ws_9 <= io_in_r_bypass_28_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_0_stall_9 <= io_in_r_bypass_28_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_1_data_9 <= io_in_r_bypass_28_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_1_load_store_9 <= io_in_r_bypass_28_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_1_df_is_ws_9 <= io_in_r_bypass_28_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_1_stall_9 <= io_in_r_bypass_28_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_2_data_9 <= io_in_r_bypass_28_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_2_load_store_9 <= io_in_r_bypass_28_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_2_df_is_ws_9 <= io_in_r_bypass_28_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_2_stall_9 <= io_in_r_bypass_28_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_3_data_9 <= io_in_r_bypass_28_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_3_load_store_9 <= io_in_r_bypass_28_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_3_df_is_ws_9 <= io_in_r_bypass_28_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_3_stall_9 <= io_in_r_bypass_28_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_0_data_9 <= io_in_r_bypass_29_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_0_load_store_9 <= io_in_r_bypass_29_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_0_df_is_ws_9 <= io_in_r_bypass_29_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_0_stall_9 <= io_in_r_bypass_29_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_1_data_9 <= io_in_r_bypass_29_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_1_load_store_9 <= io_in_r_bypass_29_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_1_df_is_ws_9 <= io_in_r_bypass_29_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_1_stall_9 <= io_in_r_bypass_29_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_2_data_9 <= io_in_r_bypass_29_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_2_load_store_9 <= io_in_r_bypass_29_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_2_df_is_ws_9 <= io_in_r_bypass_29_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_2_stall_9 <= io_in_r_bypass_29_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_3_data_9 <= io_in_r_bypass_29_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_3_load_store_9 <= io_in_r_bypass_29_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_3_df_is_ws_9 <= io_in_r_bypass_29_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_3_stall_9 <= io_in_r_bypass_29_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_0_data_9 <= io_in_r_bypass_30_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_0_load_store_9 <= io_in_r_bypass_30_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_0_df_is_ws_9 <= io_in_r_bypass_30_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_0_stall_9 <= io_in_r_bypass_30_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_1_data_9 <= io_in_r_bypass_30_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_1_load_store_9 <= io_in_r_bypass_30_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_1_df_is_ws_9 <= io_in_r_bypass_30_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_1_stall_9 <= io_in_r_bypass_30_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_2_data_9 <= io_in_r_bypass_30_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_2_load_store_9 <= io_in_r_bypass_30_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_2_df_is_ws_9 <= io_in_r_bypass_30_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_2_stall_9 <= io_in_r_bypass_30_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_3_data_9 <= io_in_r_bypass_30_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_3_load_store_9 <= io_in_r_bypass_30_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_3_df_is_ws_9 <= io_in_r_bypass_30_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_3_stall_9 <= io_in_r_bypass_30_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_0_data_9 <= io_in_r_bypass_31_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_0_load_store_9 <= io_in_r_bypass_31_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_0_df_is_ws_9 <= io_in_r_bypass_31_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_0_stall_9 <= io_in_r_bypass_31_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_1_data_9 <= io_in_r_bypass_31_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_1_load_store_9 <= io_in_r_bypass_31_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_1_df_is_ws_9 <= io_in_r_bypass_31_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_1_stall_9 <= io_in_r_bypass_31_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_2_data_9 <= io_in_r_bypass_31_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_2_load_store_9 <= io_in_r_bypass_31_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_2_df_is_ws_9 <= io_in_r_bypass_31_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_2_stall_9 <= io_in_r_bypass_31_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_3_data_9 <= io_in_r_bypass_31_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_3_load_store_9 <= io_in_r_bypass_31_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_3_df_is_ws_9 <= io_in_r_bypass_31_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_3_stall_9 <= io_in_r_bypass_31_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_0_data_10 <= io_in_r_bypass_0_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_0_load_store_10 <= io_in_r_bypass_0_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_0_df_is_ws_10 <= io_in_r_bypass_0_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_0_stall_10 <= io_in_r_bypass_0_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_1_data_10 <= io_in_r_bypass_0_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_1_load_store_10 <= io_in_r_bypass_0_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_1_df_is_ws_10 <= io_in_r_bypass_0_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_1_stall_10 <= io_in_r_bypass_0_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_2_data_10 <= io_in_r_bypass_0_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_2_load_store_10 <= io_in_r_bypass_0_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_2_df_is_ws_10 <= io_in_r_bypass_0_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_2_stall_10 <= io_in_r_bypass_0_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_3_data_10 <= io_in_r_bypass_0_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_3_load_store_10 <= io_in_r_bypass_0_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_3_df_is_ws_10 <= io_in_r_bypass_0_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_3_stall_10 <= io_in_r_bypass_0_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_0_data_10 <= io_in_r_bypass_1_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_0_load_store_10 <= io_in_r_bypass_1_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_0_df_is_ws_10 <= io_in_r_bypass_1_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_0_stall_10 <= io_in_r_bypass_1_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_1_data_10 <= io_in_r_bypass_1_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_1_load_store_10 <= io_in_r_bypass_1_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_1_df_is_ws_10 <= io_in_r_bypass_1_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_1_stall_10 <= io_in_r_bypass_1_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_2_data_10 <= io_in_r_bypass_1_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_2_load_store_10 <= io_in_r_bypass_1_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_2_df_is_ws_10 <= io_in_r_bypass_1_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_2_stall_10 <= io_in_r_bypass_1_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_3_data_10 <= io_in_r_bypass_1_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_3_load_store_10 <= io_in_r_bypass_1_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_3_df_is_ws_10 <= io_in_r_bypass_1_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_3_stall_10 <= io_in_r_bypass_1_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_0_data_10 <= io_in_r_bypass_2_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_0_load_store_10 <= io_in_r_bypass_2_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_0_df_is_ws_10 <= io_in_r_bypass_2_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_0_stall_10 <= io_in_r_bypass_2_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_1_data_10 <= io_in_r_bypass_2_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_1_load_store_10 <= io_in_r_bypass_2_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_1_df_is_ws_10 <= io_in_r_bypass_2_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_1_stall_10 <= io_in_r_bypass_2_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_2_data_10 <= io_in_r_bypass_2_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_2_load_store_10 <= io_in_r_bypass_2_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_2_df_is_ws_10 <= io_in_r_bypass_2_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_2_stall_10 <= io_in_r_bypass_2_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_3_data_10 <= io_in_r_bypass_2_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_3_load_store_10 <= io_in_r_bypass_2_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_3_df_is_ws_10 <= io_in_r_bypass_2_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_3_stall_10 <= io_in_r_bypass_2_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_0_data_10 <= io_in_r_bypass_3_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_0_load_store_10 <= io_in_r_bypass_3_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_0_df_is_ws_10 <= io_in_r_bypass_3_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_0_stall_10 <= io_in_r_bypass_3_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_1_data_10 <= io_in_r_bypass_3_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_1_load_store_10 <= io_in_r_bypass_3_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_1_df_is_ws_10 <= io_in_r_bypass_3_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_1_stall_10 <= io_in_r_bypass_3_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_2_data_10 <= io_in_r_bypass_3_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_2_load_store_10 <= io_in_r_bypass_3_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_2_df_is_ws_10 <= io_in_r_bypass_3_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_2_stall_10 <= io_in_r_bypass_3_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_3_data_10 <= io_in_r_bypass_3_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_3_load_store_10 <= io_in_r_bypass_3_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_3_df_is_ws_10 <= io_in_r_bypass_3_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_3_stall_10 <= io_in_r_bypass_3_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_0_data_10 <= io_in_r_bypass_4_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_0_load_store_10 <= io_in_r_bypass_4_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_0_df_is_ws_10 <= io_in_r_bypass_4_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_0_stall_10 <= io_in_r_bypass_4_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_1_data_10 <= io_in_r_bypass_4_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_1_load_store_10 <= io_in_r_bypass_4_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_1_df_is_ws_10 <= io_in_r_bypass_4_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_1_stall_10 <= io_in_r_bypass_4_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_2_data_10 <= io_in_r_bypass_4_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_2_load_store_10 <= io_in_r_bypass_4_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_2_df_is_ws_10 <= io_in_r_bypass_4_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_2_stall_10 <= io_in_r_bypass_4_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_3_data_10 <= io_in_r_bypass_4_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_3_load_store_10 <= io_in_r_bypass_4_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_3_df_is_ws_10 <= io_in_r_bypass_4_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_3_stall_10 <= io_in_r_bypass_4_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_0_data_10 <= io_in_r_bypass_5_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_0_load_store_10 <= io_in_r_bypass_5_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_0_df_is_ws_10 <= io_in_r_bypass_5_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_0_stall_10 <= io_in_r_bypass_5_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_1_data_10 <= io_in_r_bypass_5_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_1_load_store_10 <= io_in_r_bypass_5_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_1_df_is_ws_10 <= io_in_r_bypass_5_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_1_stall_10 <= io_in_r_bypass_5_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_2_data_10 <= io_in_r_bypass_5_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_2_load_store_10 <= io_in_r_bypass_5_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_2_df_is_ws_10 <= io_in_r_bypass_5_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_2_stall_10 <= io_in_r_bypass_5_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_3_data_10 <= io_in_r_bypass_5_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_3_load_store_10 <= io_in_r_bypass_5_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_3_df_is_ws_10 <= io_in_r_bypass_5_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_3_stall_10 <= io_in_r_bypass_5_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_0_data_10 <= io_in_r_bypass_6_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_0_load_store_10 <= io_in_r_bypass_6_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_0_df_is_ws_10 <= io_in_r_bypass_6_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_0_stall_10 <= io_in_r_bypass_6_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_1_data_10 <= io_in_r_bypass_6_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_1_load_store_10 <= io_in_r_bypass_6_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_1_df_is_ws_10 <= io_in_r_bypass_6_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_1_stall_10 <= io_in_r_bypass_6_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_2_data_10 <= io_in_r_bypass_6_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_2_load_store_10 <= io_in_r_bypass_6_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_2_df_is_ws_10 <= io_in_r_bypass_6_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_2_stall_10 <= io_in_r_bypass_6_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_3_data_10 <= io_in_r_bypass_6_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_3_load_store_10 <= io_in_r_bypass_6_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_3_df_is_ws_10 <= io_in_r_bypass_6_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_3_stall_10 <= io_in_r_bypass_6_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_0_data_10 <= io_in_r_bypass_7_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_0_load_store_10 <= io_in_r_bypass_7_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_0_df_is_ws_10 <= io_in_r_bypass_7_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_0_stall_10 <= io_in_r_bypass_7_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_1_data_10 <= io_in_r_bypass_7_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_1_load_store_10 <= io_in_r_bypass_7_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_1_df_is_ws_10 <= io_in_r_bypass_7_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_1_stall_10 <= io_in_r_bypass_7_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_2_data_10 <= io_in_r_bypass_7_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_2_load_store_10 <= io_in_r_bypass_7_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_2_df_is_ws_10 <= io_in_r_bypass_7_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_2_stall_10 <= io_in_r_bypass_7_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_3_data_10 <= io_in_r_bypass_7_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_3_load_store_10 <= io_in_r_bypass_7_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_3_df_is_ws_10 <= io_in_r_bypass_7_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_3_stall_10 <= io_in_r_bypass_7_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_0_data_10 <= io_in_r_bypass_8_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_0_load_store_10 <= io_in_r_bypass_8_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_0_df_is_ws_10 <= io_in_r_bypass_8_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_0_stall_10 <= io_in_r_bypass_8_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_1_data_10 <= io_in_r_bypass_8_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_1_load_store_10 <= io_in_r_bypass_8_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_1_df_is_ws_10 <= io_in_r_bypass_8_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_1_stall_10 <= io_in_r_bypass_8_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_2_data_10 <= io_in_r_bypass_8_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_2_load_store_10 <= io_in_r_bypass_8_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_2_df_is_ws_10 <= io_in_r_bypass_8_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_2_stall_10 <= io_in_r_bypass_8_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_3_data_10 <= io_in_r_bypass_8_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_3_load_store_10 <= io_in_r_bypass_8_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_3_df_is_ws_10 <= io_in_r_bypass_8_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_3_stall_10 <= io_in_r_bypass_8_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_0_data_10 <= io_in_r_bypass_9_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_0_load_store_10 <= io_in_r_bypass_9_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_0_df_is_ws_10 <= io_in_r_bypass_9_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_0_stall_10 <= io_in_r_bypass_9_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_1_data_10 <= io_in_r_bypass_9_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_1_load_store_10 <= io_in_r_bypass_9_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_1_df_is_ws_10 <= io_in_r_bypass_9_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_1_stall_10 <= io_in_r_bypass_9_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_2_data_10 <= io_in_r_bypass_9_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_2_load_store_10 <= io_in_r_bypass_9_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_2_df_is_ws_10 <= io_in_r_bypass_9_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_2_stall_10 <= io_in_r_bypass_9_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_3_data_10 <= io_in_r_bypass_9_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_3_load_store_10 <= io_in_r_bypass_9_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_3_df_is_ws_10 <= io_in_r_bypass_9_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_3_stall_10 <= io_in_r_bypass_9_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_0_data_10 <= io_in_r_bypass_10_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_0_load_store_10 <= io_in_r_bypass_10_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_0_df_is_ws_10 <= io_in_r_bypass_10_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_0_stall_10 <= io_in_r_bypass_10_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_1_data_10 <= io_in_r_bypass_10_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_1_load_store_10 <= io_in_r_bypass_10_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_1_df_is_ws_10 <= io_in_r_bypass_10_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_1_stall_10 <= io_in_r_bypass_10_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_2_data_10 <= io_in_r_bypass_10_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_2_load_store_10 <= io_in_r_bypass_10_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_2_df_is_ws_10 <= io_in_r_bypass_10_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_2_stall_10 <= io_in_r_bypass_10_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_3_data_10 <= io_in_r_bypass_10_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_3_load_store_10 <= io_in_r_bypass_10_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_3_df_is_ws_10 <= io_in_r_bypass_10_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_3_stall_10 <= io_in_r_bypass_10_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_0_data_10 <= io_in_r_bypass_11_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_0_load_store_10 <= io_in_r_bypass_11_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_0_df_is_ws_10 <= io_in_r_bypass_11_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_0_stall_10 <= io_in_r_bypass_11_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_1_data_10 <= io_in_r_bypass_11_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_1_load_store_10 <= io_in_r_bypass_11_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_1_df_is_ws_10 <= io_in_r_bypass_11_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_1_stall_10 <= io_in_r_bypass_11_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_2_data_10 <= io_in_r_bypass_11_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_2_load_store_10 <= io_in_r_bypass_11_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_2_df_is_ws_10 <= io_in_r_bypass_11_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_2_stall_10 <= io_in_r_bypass_11_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_3_data_10 <= io_in_r_bypass_11_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_3_load_store_10 <= io_in_r_bypass_11_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_3_df_is_ws_10 <= io_in_r_bypass_11_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_3_stall_10 <= io_in_r_bypass_11_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_0_data_10 <= io_in_r_bypass_12_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_0_load_store_10 <= io_in_r_bypass_12_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_0_df_is_ws_10 <= io_in_r_bypass_12_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_0_stall_10 <= io_in_r_bypass_12_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_1_data_10 <= io_in_r_bypass_12_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_1_load_store_10 <= io_in_r_bypass_12_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_1_df_is_ws_10 <= io_in_r_bypass_12_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_1_stall_10 <= io_in_r_bypass_12_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_2_data_10 <= io_in_r_bypass_12_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_2_load_store_10 <= io_in_r_bypass_12_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_2_df_is_ws_10 <= io_in_r_bypass_12_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_2_stall_10 <= io_in_r_bypass_12_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_3_data_10 <= io_in_r_bypass_12_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_3_load_store_10 <= io_in_r_bypass_12_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_3_df_is_ws_10 <= io_in_r_bypass_12_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_3_stall_10 <= io_in_r_bypass_12_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_0_data_10 <= io_in_r_bypass_13_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_0_load_store_10 <= io_in_r_bypass_13_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_0_df_is_ws_10 <= io_in_r_bypass_13_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_0_stall_10 <= io_in_r_bypass_13_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_1_data_10 <= io_in_r_bypass_13_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_1_load_store_10 <= io_in_r_bypass_13_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_1_df_is_ws_10 <= io_in_r_bypass_13_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_1_stall_10 <= io_in_r_bypass_13_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_2_data_10 <= io_in_r_bypass_13_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_2_load_store_10 <= io_in_r_bypass_13_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_2_df_is_ws_10 <= io_in_r_bypass_13_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_2_stall_10 <= io_in_r_bypass_13_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_3_data_10 <= io_in_r_bypass_13_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_3_load_store_10 <= io_in_r_bypass_13_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_3_df_is_ws_10 <= io_in_r_bypass_13_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_3_stall_10 <= io_in_r_bypass_13_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_0_data_10 <= io_in_r_bypass_14_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_0_load_store_10 <= io_in_r_bypass_14_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_0_df_is_ws_10 <= io_in_r_bypass_14_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_0_stall_10 <= io_in_r_bypass_14_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_1_data_10 <= io_in_r_bypass_14_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_1_load_store_10 <= io_in_r_bypass_14_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_1_df_is_ws_10 <= io_in_r_bypass_14_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_1_stall_10 <= io_in_r_bypass_14_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_2_data_10 <= io_in_r_bypass_14_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_2_load_store_10 <= io_in_r_bypass_14_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_2_df_is_ws_10 <= io_in_r_bypass_14_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_2_stall_10 <= io_in_r_bypass_14_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_3_data_10 <= io_in_r_bypass_14_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_3_load_store_10 <= io_in_r_bypass_14_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_3_df_is_ws_10 <= io_in_r_bypass_14_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_3_stall_10 <= io_in_r_bypass_14_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_0_data_10 <= io_in_r_bypass_15_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_0_load_store_10 <= io_in_r_bypass_15_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_0_df_is_ws_10 <= io_in_r_bypass_15_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_0_stall_10 <= io_in_r_bypass_15_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_1_data_10 <= io_in_r_bypass_15_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_1_load_store_10 <= io_in_r_bypass_15_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_1_df_is_ws_10 <= io_in_r_bypass_15_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_1_stall_10 <= io_in_r_bypass_15_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_2_data_10 <= io_in_r_bypass_15_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_2_load_store_10 <= io_in_r_bypass_15_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_2_df_is_ws_10 <= io_in_r_bypass_15_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_2_stall_10 <= io_in_r_bypass_15_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_3_data_10 <= io_in_r_bypass_15_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_3_load_store_10 <= io_in_r_bypass_15_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_3_df_is_ws_10 <= io_in_r_bypass_15_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_3_stall_10 <= io_in_r_bypass_15_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_0_data_10 <= io_in_r_bypass_16_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_0_load_store_10 <= io_in_r_bypass_16_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_0_df_is_ws_10 <= io_in_r_bypass_16_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_0_stall_10 <= io_in_r_bypass_16_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_1_data_10 <= io_in_r_bypass_16_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_1_load_store_10 <= io_in_r_bypass_16_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_1_df_is_ws_10 <= io_in_r_bypass_16_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_1_stall_10 <= io_in_r_bypass_16_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_2_data_10 <= io_in_r_bypass_16_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_2_load_store_10 <= io_in_r_bypass_16_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_2_df_is_ws_10 <= io_in_r_bypass_16_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_2_stall_10 <= io_in_r_bypass_16_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_3_data_10 <= io_in_r_bypass_16_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_3_load_store_10 <= io_in_r_bypass_16_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_3_df_is_ws_10 <= io_in_r_bypass_16_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_3_stall_10 <= io_in_r_bypass_16_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_0_data_10 <= io_in_r_bypass_17_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_0_load_store_10 <= io_in_r_bypass_17_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_0_df_is_ws_10 <= io_in_r_bypass_17_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_0_stall_10 <= io_in_r_bypass_17_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_1_data_10 <= io_in_r_bypass_17_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_1_load_store_10 <= io_in_r_bypass_17_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_1_df_is_ws_10 <= io_in_r_bypass_17_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_1_stall_10 <= io_in_r_bypass_17_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_2_data_10 <= io_in_r_bypass_17_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_2_load_store_10 <= io_in_r_bypass_17_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_2_df_is_ws_10 <= io_in_r_bypass_17_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_2_stall_10 <= io_in_r_bypass_17_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_3_data_10 <= io_in_r_bypass_17_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_3_load_store_10 <= io_in_r_bypass_17_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_3_df_is_ws_10 <= io_in_r_bypass_17_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_3_stall_10 <= io_in_r_bypass_17_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_0_data_10 <= io_in_r_bypass_18_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_0_load_store_10 <= io_in_r_bypass_18_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_0_df_is_ws_10 <= io_in_r_bypass_18_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_0_stall_10 <= io_in_r_bypass_18_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_1_data_10 <= io_in_r_bypass_18_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_1_load_store_10 <= io_in_r_bypass_18_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_1_df_is_ws_10 <= io_in_r_bypass_18_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_1_stall_10 <= io_in_r_bypass_18_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_2_data_10 <= io_in_r_bypass_18_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_2_load_store_10 <= io_in_r_bypass_18_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_2_df_is_ws_10 <= io_in_r_bypass_18_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_2_stall_10 <= io_in_r_bypass_18_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_3_data_10 <= io_in_r_bypass_18_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_3_load_store_10 <= io_in_r_bypass_18_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_3_df_is_ws_10 <= io_in_r_bypass_18_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_3_stall_10 <= io_in_r_bypass_18_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_0_data_10 <= io_in_r_bypass_19_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_0_load_store_10 <= io_in_r_bypass_19_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_0_df_is_ws_10 <= io_in_r_bypass_19_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_0_stall_10 <= io_in_r_bypass_19_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_1_data_10 <= io_in_r_bypass_19_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_1_load_store_10 <= io_in_r_bypass_19_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_1_df_is_ws_10 <= io_in_r_bypass_19_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_1_stall_10 <= io_in_r_bypass_19_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_2_data_10 <= io_in_r_bypass_19_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_2_load_store_10 <= io_in_r_bypass_19_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_2_df_is_ws_10 <= io_in_r_bypass_19_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_2_stall_10 <= io_in_r_bypass_19_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_3_data_10 <= io_in_r_bypass_19_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_3_load_store_10 <= io_in_r_bypass_19_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_3_df_is_ws_10 <= io_in_r_bypass_19_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_3_stall_10 <= io_in_r_bypass_19_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_0_data_10 <= io_in_r_bypass_20_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_0_load_store_10 <= io_in_r_bypass_20_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_0_df_is_ws_10 <= io_in_r_bypass_20_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_0_stall_10 <= io_in_r_bypass_20_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_1_data_10 <= io_in_r_bypass_20_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_1_load_store_10 <= io_in_r_bypass_20_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_1_df_is_ws_10 <= io_in_r_bypass_20_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_1_stall_10 <= io_in_r_bypass_20_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_2_data_10 <= io_in_r_bypass_20_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_2_load_store_10 <= io_in_r_bypass_20_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_2_df_is_ws_10 <= io_in_r_bypass_20_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_2_stall_10 <= io_in_r_bypass_20_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_3_data_10 <= io_in_r_bypass_20_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_3_load_store_10 <= io_in_r_bypass_20_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_3_df_is_ws_10 <= io_in_r_bypass_20_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_3_stall_10 <= io_in_r_bypass_20_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_0_data_10 <= io_in_r_bypass_21_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_0_load_store_10 <= io_in_r_bypass_21_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_0_df_is_ws_10 <= io_in_r_bypass_21_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_0_stall_10 <= io_in_r_bypass_21_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_1_data_10 <= io_in_r_bypass_21_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_1_load_store_10 <= io_in_r_bypass_21_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_1_df_is_ws_10 <= io_in_r_bypass_21_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_1_stall_10 <= io_in_r_bypass_21_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_2_data_10 <= io_in_r_bypass_21_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_2_load_store_10 <= io_in_r_bypass_21_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_2_df_is_ws_10 <= io_in_r_bypass_21_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_2_stall_10 <= io_in_r_bypass_21_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_3_data_10 <= io_in_r_bypass_21_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_3_load_store_10 <= io_in_r_bypass_21_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_3_df_is_ws_10 <= io_in_r_bypass_21_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_3_stall_10 <= io_in_r_bypass_21_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_0_data_10 <= io_in_r_bypass_22_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_0_load_store_10 <= io_in_r_bypass_22_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_0_df_is_ws_10 <= io_in_r_bypass_22_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_0_stall_10 <= io_in_r_bypass_22_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_1_data_10 <= io_in_r_bypass_22_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_1_load_store_10 <= io_in_r_bypass_22_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_1_df_is_ws_10 <= io_in_r_bypass_22_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_1_stall_10 <= io_in_r_bypass_22_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_2_data_10 <= io_in_r_bypass_22_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_2_load_store_10 <= io_in_r_bypass_22_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_2_df_is_ws_10 <= io_in_r_bypass_22_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_2_stall_10 <= io_in_r_bypass_22_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_3_data_10 <= io_in_r_bypass_22_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_3_load_store_10 <= io_in_r_bypass_22_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_3_df_is_ws_10 <= io_in_r_bypass_22_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_3_stall_10 <= io_in_r_bypass_22_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_0_data_10 <= io_in_r_bypass_23_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_0_load_store_10 <= io_in_r_bypass_23_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_0_df_is_ws_10 <= io_in_r_bypass_23_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_0_stall_10 <= io_in_r_bypass_23_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_1_data_10 <= io_in_r_bypass_23_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_1_load_store_10 <= io_in_r_bypass_23_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_1_df_is_ws_10 <= io_in_r_bypass_23_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_1_stall_10 <= io_in_r_bypass_23_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_2_data_10 <= io_in_r_bypass_23_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_2_load_store_10 <= io_in_r_bypass_23_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_2_df_is_ws_10 <= io_in_r_bypass_23_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_2_stall_10 <= io_in_r_bypass_23_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_3_data_10 <= io_in_r_bypass_23_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_3_load_store_10 <= io_in_r_bypass_23_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_3_df_is_ws_10 <= io_in_r_bypass_23_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_3_stall_10 <= io_in_r_bypass_23_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_0_data_10 <= io_in_r_bypass_24_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_0_load_store_10 <= io_in_r_bypass_24_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_0_df_is_ws_10 <= io_in_r_bypass_24_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_0_stall_10 <= io_in_r_bypass_24_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_1_data_10 <= io_in_r_bypass_24_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_1_load_store_10 <= io_in_r_bypass_24_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_1_df_is_ws_10 <= io_in_r_bypass_24_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_1_stall_10 <= io_in_r_bypass_24_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_2_data_10 <= io_in_r_bypass_24_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_2_load_store_10 <= io_in_r_bypass_24_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_2_df_is_ws_10 <= io_in_r_bypass_24_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_2_stall_10 <= io_in_r_bypass_24_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_3_data_10 <= io_in_r_bypass_24_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_3_load_store_10 <= io_in_r_bypass_24_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_3_df_is_ws_10 <= io_in_r_bypass_24_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_3_stall_10 <= io_in_r_bypass_24_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_0_data_10 <= io_in_r_bypass_25_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_0_load_store_10 <= io_in_r_bypass_25_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_0_df_is_ws_10 <= io_in_r_bypass_25_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_0_stall_10 <= io_in_r_bypass_25_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_1_data_10 <= io_in_r_bypass_25_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_1_load_store_10 <= io_in_r_bypass_25_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_1_df_is_ws_10 <= io_in_r_bypass_25_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_1_stall_10 <= io_in_r_bypass_25_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_2_data_10 <= io_in_r_bypass_25_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_2_load_store_10 <= io_in_r_bypass_25_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_2_df_is_ws_10 <= io_in_r_bypass_25_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_2_stall_10 <= io_in_r_bypass_25_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_3_data_10 <= io_in_r_bypass_25_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_3_load_store_10 <= io_in_r_bypass_25_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_3_df_is_ws_10 <= io_in_r_bypass_25_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_3_stall_10 <= io_in_r_bypass_25_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_0_data_10 <= io_in_r_bypass_26_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_0_load_store_10 <= io_in_r_bypass_26_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_0_df_is_ws_10 <= io_in_r_bypass_26_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_0_stall_10 <= io_in_r_bypass_26_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_1_data_10 <= io_in_r_bypass_26_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_1_load_store_10 <= io_in_r_bypass_26_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_1_df_is_ws_10 <= io_in_r_bypass_26_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_1_stall_10 <= io_in_r_bypass_26_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_2_data_10 <= io_in_r_bypass_26_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_2_load_store_10 <= io_in_r_bypass_26_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_2_df_is_ws_10 <= io_in_r_bypass_26_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_2_stall_10 <= io_in_r_bypass_26_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_3_data_10 <= io_in_r_bypass_26_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_3_load_store_10 <= io_in_r_bypass_26_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_3_df_is_ws_10 <= io_in_r_bypass_26_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_3_stall_10 <= io_in_r_bypass_26_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_0_data_10 <= io_in_r_bypass_27_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_0_load_store_10 <= io_in_r_bypass_27_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_0_df_is_ws_10 <= io_in_r_bypass_27_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_0_stall_10 <= io_in_r_bypass_27_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_1_data_10 <= io_in_r_bypass_27_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_1_load_store_10 <= io_in_r_bypass_27_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_1_df_is_ws_10 <= io_in_r_bypass_27_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_1_stall_10 <= io_in_r_bypass_27_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_2_data_10 <= io_in_r_bypass_27_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_2_load_store_10 <= io_in_r_bypass_27_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_2_df_is_ws_10 <= io_in_r_bypass_27_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_2_stall_10 <= io_in_r_bypass_27_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_3_data_10 <= io_in_r_bypass_27_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_3_load_store_10 <= io_in_r_bypass_27_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_3_df_is_ws_10 <= io_in_r_bypass_27_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_3_stall_10 <= io_in_r_bypass_27_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_0_data_10 <= io_in_r_bypass_28_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_0_load_store_10 <= io_in_r_bypass_28_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_0_df_is_ws_10 <= io_in_r_bypass_28_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_0_stall_10 <= io_in_r_bypass_28_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_1_data_10 <= io_in_r_bypass_28_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_1_load_store_10 <= io_in_r_bypass_28_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_1_df_is_ws_10 <= io_in_r_bypass_28_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_1_stall_10 <= io_in_r_bypass_28_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_2_data_10 <= io_in_r_bypass_28_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_2_load_store_10 <= io_in_r_bypass_28_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_2_df_is_ws_10 <= io_in_r_bypass_28_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_2_stall_10 <= io_in_r_bypass_28_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_3_data_10 <= io_in_r_bypass_28_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_3_load_store_10 <= io_in_r_bypass_28_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_3_df_is_ws_10 <= io_in_r_bypass_28_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_3_stall_10 <= io_in_r_bypass_28_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_0_data_10 <= io_in_r_bypass_29_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_0_load_store_10 <= io_in_r_bypass_29_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_0_df_is_ws_10 <= io_in_r_bypass_29_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_0_stall_10 <= io_in_r_bypass_29_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_1_data_10 <= io_in_r_bypass_29_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_1_load_store_10 <= io_in_r_bypass_29_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_1_df_is_ws_10 <= io_in_r_bypass_29_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_1_stall_10 <= io_in_r_bypass_29_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_2_data_10 <= io_in_r_bypass_29_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_2_load_store_10 <= io_in_r_bypass_29_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_2_df_is_ws_10 <= io_in_r_bypass_29_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_2_stall_10 <= io_in_r_bypass_29_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_3_data_10 <= io_in_r_bypass_29_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_3_load_store_10 <= io_in_r_bypass_29_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_3_df_is_ws_10 <= io_in_r_bypass_29_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_3_stall_10 <= io_in_r_bypass_29_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_0_data_10 <= io_in_r_bypass_30_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_0_load_store_10 <= io_in_r_bypass_30_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_0_df_is_ws_10 <= io_in_r_bypass_30_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_0_stall_10 <= io_in_r_bypass_30_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_1_data_10 <= io_in_r_bypass_30_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_1_load_store_10 <= io_in_r_bypass_30_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_1_df_is_ws_10 <= io_in_r_bypass_30_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_1_stall_10 <= io_in_r_bypass_30_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_2_data_10 <= io_in_r_bypass_30_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_2_load_store_10 <= io_in_r_bypass_30_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_2_df_is_ws_10 <= io_in_r_bypass_30_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_2_stall_10 <= io_in_r_bypass_30_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_3_data_10 <= io_in_r_bypass_30_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_3_load_store_10 <= io_in_r_bypass_30_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_3_df_is_ws_10 <= io_in_r_bypass_30_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_3_stall_10 <= io_in_r_bypass_30_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_0_data_10 <= io_in_r_bypass_31_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_0_load_store_10 <= io_in_r_bypass_31_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_0_df_is_ws_10 <= io_in_r_bypass_31_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_0_stall_10 <= io_in_r_bypass_31_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_1_data_10 <= io_in_r_bypass_31_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_1_load_store_10 <= io_in_r_bypass_31_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_1_df_is_ws_10 <= io_in_r_bypass_31_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_1_stall_10 <= io_in_r_bypass_31_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_2_data_10 <= io_in_r_bypass_31_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_2_load_store_10 <= io_in_r_bypass_31_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_2_df_is_ws_10 <= io_in_r_bypass_31_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_2_stall_10 <= io_in_r_bypass_31_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_3_data_10 <= io_in_r_bypass_31_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_3_load_store_10 <= io_in_r_bypass_31_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_3_df_is_ws_10 <= io_in_r_bypass_31_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_3_stall_10 <= io_in_r_bypass_31_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_0_data_11 <= io_in_r_bypass_0_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_0_load_store_11 <= io_in_r_bypass_0_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_0_df_is_ws_11 <= io_in_r_bypass_0_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_0_stall_11 <= io_in_r_bypass_0_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_1_data_11 <= io_in_r_bypass_0_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_1_load_store_11 <= io_in_r_bypass_0_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_1_df_is_ws_11 <= io_in_r_bypass_0_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_1_stall_11 <= io_in_r_bypass_0_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_2_data_11 <= io_in_r_bypass_0_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_2_load_store_11 <= io_in_r_bypass_0_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_2_df_is_ws_11 <= io_in_r_bypass_0_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_2_stall_11 <= io_in_r_bypass_0_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_3_data_11 <= io_in_r_bypass_0_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_3_load_store_11 <= io_in_r_bypass_0_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_3_df_is_ws_11 <= io_in_r_bypass_0_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_3_stall_11 <= io_in_r_bypass_0_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_0_data_11 <= io_in_r_bypass_1_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_0_load_store_11 <= io_in_r_bypass_1_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_0_df_is_ws_11 <= io_in_r_bypass_1_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_0_stall_11 <= io_in_r_bypass_1_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_1_data_11 <= io_in_r_bypass_1_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_1_load_store_11 <= io_in_r_bypass_1_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_1_df_is_ws_11 <= io_in_r_bypass_1_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_1_stall_11 <= io_in_r_bypass_1_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_2_data_11 <= io_in_r_bypass_1_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_2_load_store_11 <= io_in_r_bypass_1_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_2_df_is_ws_11 <= io_in_r_bypass_1_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_2_stall_11 <= io_in_r_bypass_1_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_3_data_11 <= io_in_r_bypass_1_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_3_load_store_11 <= io_in_r_bypass_1_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_3_df_is_ws_11 <= io_in_r_bypass_1_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_3_stall_11 <= io_in_r_bypass_1_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_0_data_11 <= io_in_r_bypass_2_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_0_load_store_11 <= io_in_r_bypass_2_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_0_df_is_ws_11 <= io_in_r_bypass_2_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_0_stall_11 <= io_in_r_bypass_2_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_1_data_11 <= io_in_r_bypass_2_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_1_load_store_11 <= io_in_r_bypass_2_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_1_df_is_ws_11 <= io_in_r_bypass_2_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_1_stall_11 <= io_in_r_bypass_2_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_2_data_11 <= io_in_r_bypass_2_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_2_load_store_11 <= io_in_r_bypass_2_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_2_df_is_ws_11 <= io_in_r_bypass_2_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_2_stall_11 <= io_in_r_bypass_2_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_3_data_11 <= io_in_r_bypass_2_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_3_load_store_11 <= io_in_r_bypass_2_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_3_df_is_ws_11 <= io_in_r_bypass_2_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_3_stall_11 <= io_in_r_bypass_2_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_0_data_11 <= io_in_r_bypass_3_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_0_load_store_11 <= io_in_r_bypass_3_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_0_df_is_ws_11 <= io_in_r_bypass_3_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_0_stall_11 <= io_in_r_bypass_3_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_1_data_11 <= io_in_r_bypass_3_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_1_load_store_11 <= io_in_r_bypass_3_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_1_df_is_ws_11 <= io_in_r_bypass_3_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_1_stall_11 <= io_in_r_bypass_3_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_2_data_11 <= io_in_r_bypass_3_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_2_load_store_11 <= io_in_r_bypass_3_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_2_df_is_ws_11 <= io_in_r_bypass_3_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_2_stall_11 <= io_in_r_bypass_3_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_3_data_11 <= io_in_r_bypass_3_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_3_load_store_11 <= io_in_r_bypass_3_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_3_df_is_ws_11 <= io_in_r_bypass_3_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_3_stall_11 <= io_in_r_bypass_3_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_0_data_11 <= io_in_r_bypass_4_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_0_load_store_11 <= io_in_r_bypass_4_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_0_df_is_ws_11 <= io_in_r_bypass_4_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_0_stall_11 <= io_in_r_bypass_4_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_1_data_11 <= io_in_r_bypass_4_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_1_load_store_11 <= io_in_r_bypass_4_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_1_df_is_ws_11 <= io_in_r_bypass_4_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_1_stall_11 <= io_in_r_bypass_4_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_2_data_11 <= io_in_r_bypass_4_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_2_load_store_11 <= io_in_r_bypass_4_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_2_df_is_ws_11 <= io_in_r_bypass_4_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_2_stall_11 <= io_in_r_bypass_4_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_3_data_11 <= io_in_r_bypass_4_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_3_load_store_11 <= io_in_r_bypass_4_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_3_df_is_ws_11 <= io_in_r_bypass_4_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_3_stall_11 <= io_in_r_bypass_4_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_0_data_11 <= io_in_r_bypass_5_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_0_load_store_11 <= io_in_r_bypass_5_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_0_df_is_ws_11 <= io_in_r_bypass_5_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_0_stall_11 <= io_in_r_bypass_5_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_1_data_11 <= io_in_r_bypass_5_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_1_load_store_11 <= io_in_r_bypass_5_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_1_df_is_ws_11 <= io_in_r_bypass_5_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_1_stall_11 <= io_in_r_bypass_5_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_2_data_11 <= io_in_r_bypass_5_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_2_load_store_11 <= io_in_r_bypass_5_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_2_df_is_ws_11 <= io_in_r_bypass_5_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_2_stall_11 <= io_in_r_bypass_5_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_3_data_11 <= io_in_r_bypass_5_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_3_load_store_11 <= io_in_r_bypass_5_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_3_df_is_ws_11 <= io_in_r_bypass_5_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_3_stall_11 <= io_in_r_bypass_5_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_0_data_11 <= io_in_r_bypass_6_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_0_load_store_11 <= io_in_r_bypass_6_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_0_df_is_ws_11 <= io_in_r_bypass_6_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_0_stall_11 <= io_in_r_bypass_6_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_1_data_11 <= io_in_r_bypass_6_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_1_load_store_11 <= io_in_r_bypass_6_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_1_df_is_ws_11 <= io_in_r_bypass_6_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_1_stall_11 <= io_in_r_bypass_6_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_2_data_11 <= io_in_r_bypass_6_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_2_load_store_11 <= io_in_r_bypass_6_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_2_df_is_ws_11 <= io_in_r_bypass_6_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_2_stall_11 <= io_in_r_bypass_6_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_3_data_11 <= io_in_r_bypass_6_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_3_load_store_11 <= io_in_r_bypass_6_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_3_df_is_ws_11 <= io_in_r_bypass_6_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_3_stall_11 <= io_in_r_bypass_6_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_0_data_11 <= io_in_r_bypass_7_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_0_load_store_11 <= io_in_r_bypass_7_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_0_df_is_ws_11 <= io_in_r_bypass_7_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_0_stall_11 <= io_in_r_bypass_7_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_1_data_11 <= io_in_r_bypass_7_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_1_load_store_11 <= io_in_r_bypass_7_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_1_df_is_ws_11 <= io_in_r_bypass_7_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_1_stall_11 <= io_in_r_bypass_7_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_2_data_11 <= io_in_r_bypass_7_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_2_load_store_11 <= io_in_r_bypass_7_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_2_df_is_ws_11 <= io_in_r_bypass_7_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_2_stall_11 <= io_in_r_bypass_7_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_3_data_11 <= io_in_r_bypass_7_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_3_load_store_11 <= io_in_r_bypass_7_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_3_df_is_ws_11 <= io_in_r_bypass_7_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_3_stall_11 <= io_in_r_bypass_7_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_0_data_11 <= io_in_r_bypass_8_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_0_load_store_11 <= io_in_r_bypass_8_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_0_df_is_ws_11 <= io_in_r_bypass_8_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_0_stall_11 <= io_in_r_bypass_8_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_1_data_11 <= io_in_r_bypass_8_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_1_load_store_11 <= io_in_r_bypass_8_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_1_df_is_ws_11 <= io_in_r_bypass_8_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_1_stall_11 <= io_in_r_bypass_8_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_2_data_11 <= io_in_r_bypass_8_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_2_load_store_11 <= io_in_r_bypass_8_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_2_df_is_ws_11 <= io_in_r_bypass_8_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_2_stall_11 <= io_in_r_bypass_8_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_3_data_11 <= io_in_r_bypass_8_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_3_load_store_11 <= io_in_r_bypass_8_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_3_df_is_ws_11 <= io_in_r_bypass_8_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_3_stall_11 <= io_in_r_bypass_8_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_0_data_11 <= io_in_r_bypass_9_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_0_load_store_11 <= io_in_r_bypass_9_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_0_df_is_ws_11 <= io_in_r_bypass_9_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_0_stall_11 <= io_in_r_bypass_9_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_1_data_11 <= io_in_r_bypass_9_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_1_load_store_11 <= io_in_r_bypass_9_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_1_df_is_ws_11 <= io_in_r_bypass_9_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_1_stall_11 <= io_in_r_bypass_9_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_2_data_11 <= io_in_r_bypass_9_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_2_load_store_11 <= io_in_r_bypass_9_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_2_df_is_ws_11 <= io_in_r_bypass_9_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_2_stall_11 <= io_in_r_bypass_9_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_3_data_11 <= io_in_r_bypass_9_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_3_load_store_11 <= io_in_r_bypass_9_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_3_df_is_ws_11 <= io_in_r_bypass_9_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_3_stall_11 <= io_in_r_bypass_9_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_0_data_11 <= io_in_r_bypass_10_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_0_load_store_11 <= io_in_r_bypass_10_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_0_df_is_ws_11 <= io_in_r_bypass_10_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_0_stall_11 <= io_in_r_bypass_10_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_1_data_11 <= io_in_r_bypass_10_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_1_load_store_11 <= io_in_r_bypass_10_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_1_df_is_ws_11 <= io_in_r_bypass_10_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_1_stall_11 <= io_in_r_bypass_10_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_2_data_11 <= io_in_r_bypass_10_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_2_load_store_11 <= io_in_r_bypass_10_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_2_df_is_ws_11 <= io_in_r_bypass_10_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_2_stall_11 <= io_in_r_bypass_10_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_3_data_11 <= io_in_r_bypass_10_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_3_load_store_11 <= io_in_r_bypass_10_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_3_df_is_ws_11 <= io_in_r_bypass_10_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_3_stall_11 <= io_in_r_bypass_10_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_0_data_11 <= io_in_r_bypass_11_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_0_load_store_11 <= io_in_r_bypass_11_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_0_df_is_ws_11 <= io_in_r_bypass_11_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_0_stall_11 <= io_in_r_bypass_11_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_1_data_11 <= io_in_r_bypass_11_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_1_load_store_11 <= io_in_r_bypass_11_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_1_df_is_ws_11 <= io_in_r_bypass_11_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_1_stall_11 <= io_in_r_bypass_11_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_2_data_11 <= io_in_r_bypass_11_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_2_load_store_11 <= io_in_r_bypass_11_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_2_df_is_ws_11 <= io_in_r_bypass_11_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_2_stall_11 <= io_in_r_bypass_11_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_3_data_11 <= io_in_r_bypass_11_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_3_load_store_11 <= io_in_r_bypass_11_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_3_df_is_ws_11 <= io_in_r_bypass_11_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_3_stall_11 <= io_in_r_bypass_11_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_0_data_11 <= io_in_r_bypass_12_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_0_load_store_11 <= io_in_r_bypass_12_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_0_df_is_ws_11 <= io_in_r_bypass_12_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_0_stall_11 <= io_in_r_bypass_12_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_1_data_11 <= io_in_r_bypass_12_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_1_load_store_11 <= io_in_r_bypass_12_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_1_df_is_ws_11 <= io_in_r_bypass_12_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_1_stall_11 <= io_in_r_bypass_12_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_2_data_11 <= io_in_r_bypass_12_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_2_load_store_11 <= io_in_r_bypass_12_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_2_df_is_ws_11 <= io_in_r_bypass_12_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_2_stall_11 <= io_in_r_bypass_12_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_3_data_11 <= io_in_r_bypass_12_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_3_load_store_11 <= io_in_r_bypass_12_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_3_df_is_ws_11 <= io_in_r_bypass_12_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_3_stall_11 <= io_in_r_bypass_12_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_0_data_11 <= io_in_r_bypass_13_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_0_load_store_11 <= io_in_r_bypass_13_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_0_df_is_ws_11 <= io_in_r_bypass_13_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_0_stall_11 <= io_in_r_bypass_13_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_1_data_11 <= io_in_r_bypass_13_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_1_load_store_11 <= io_in_r_bypass_13_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_1_df_is_ws_11 <= io_in_r_bypass_13_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_1_stall_11 <= io_in_r_bypass_13_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_2_data_11 <= io_in_r_bypass_13_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_2_load_store_11 <= io_in_r_bypass_13_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_2_df_is_ws_11 <= io_in_r_bypass_13_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_2_stall_11 <= io_in_r_bypass_13_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_3_data_11 <= io_in_r_bypass_13_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_3_load_store_11 <= io_in_r_bypass_13_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_3_df_is_ws_11 <= io_in_r_bypass_13_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_3_stall_11 <= io_in_r_bypass_13_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_0_data_11 <= io_in_r_bypass_14_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_0_load_store_11 <= io_in_r_bypass_14_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_0_df_is_ws_11 <= io_in_r_bypass_14_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_0_stall_11 <= io_in_r_bypass_14_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_1_data_11 <= io_in_r_bypass_14_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_1_load_store_11 <= io_in_r_bypass_14_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_1_df_is_ws_11 <= io_in_r_bypass_14_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_1_stall_11 <= io_in_r_bypass_14_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_2_data_11 <= io_in_r_bypass_14_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_2_load_store_11 <= io_in_r_bypass_14_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_2_df_is_ws_11 <= io_in_r_bypass_14_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_2_stall_11 <= io_in_r_bypass_14_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_3_data_11 <= io_in_r_bypass_14_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_3_load_store_11 <= io_in_r_bypass_14_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_3_df_is_ws_11 <= io_in_r_bypass_14_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_3_stall_11 <= io_in_r_bypass_14_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_0_data_11 <= io_in_r_bypass_15_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_0_load_store_11 <= io_in_r_bypass_15_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_0_df_is_ws_11 <= io_in_r_bypass_15_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_0_stall_11 <= io_in_r_bypass_15_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_1_data_11 <= io_in_r_bypass_15_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_1_load_store_11 <= io_in_r_bypass_15_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_1_df_is_ws_11 <= io_in_r_bypass_15_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_1_stall_11 <= io_in_r_bypass_15_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_2_data_11 <= io_in_r_bypass_15_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_2_load_store_11 <= io_in_r_bypass_15_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_2_df_is_ws_11 <= io_in_r_bypass_15_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_2_stall_11 <= io_in_r_bypass_15_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_3_data_11 <= io_in_r_bypass_15_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_3_load_store_11 <= io_in_r_bypass_15_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_3_df_is_ws_11 <= io_in_r_bypass_15_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_3_stall_11 <= io_in_r_bypass_15_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_0_data_11 <= io_in_r_bypass_16_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_0_load_store_11 <= io_in_r_bypass_16_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_0_df_is_ws_11 <= io_in_r_bypass_16_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_0_stall_11 <= io_in_r_bypass_16_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_1_data_11 <= io_in_r_bypass_16_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_1_load_store_11 <= io_in_r_bypass_16_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_1_df_is_ws_11 <= io_in_r_bypass_16_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_1_stall_11 <= io_in_r_bypass_16_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_2_data_11 <= io_in_r_bypass_16_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_2_load_store_11 <= io_in_r_bypass_16_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_2_df_is_ws_11 <= io_in_r_bypass_16_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_2_stall_11 <= io_in_r_bypass_16_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_3_data_11 <= io_in_r_bypass_16_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_3_load_store_11 <= io_in_r_bypass_16_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_3_df_is_ws_11 <= io_in_r_bypass_16_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_3_stall_11 <= io_in_r_bypass_16_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_0_data_11 <= io_in_r_bypass_17_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_0_load_store_11 <= io_in_r_bypass_17_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_0_df_is_ws_11 <= io_in_r_bypass_17_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_0_stall_11 <= io_in_r_bypass_17_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_1_data_11 <= io_in_r_bypass_17_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_1_load_store_11 <= io_in_r_bypass_17_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_1_df_is_ws_11 <= io_in_r_bypass_17_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_1_stall_11 <= io_in_r_bypass_17_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_2_data_11 <= io_in_r_bypass_17_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_2_load_store_11 <= io_in_r_bypass_17_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_2_df_is_ws_11 <= io_in_r_bypass_17_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_2_stall_11 <= io_in_r_bypass_17_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_3_data_11 <= io_in_r_bypass_17_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_3_load_store_11 <= io_in_r_bypass_17_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_3_df_is_ws_11 <= io_in_r_bypass_17_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_3_stall_11 <= io_in_r_bypass_17_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_0_data_11 <= io_in_r_bypass_18_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_0_load_store_11 <= io_in_r_bypass_18_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_0_df_is_ws_11 <= io_in_r_bypass_18_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_0_stall_11 <= io_in_r_bypass_18_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_1_data_11 <= io_in_r_bypass_18_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_1_load_store_11 <= io_in_r_bypass_18_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_1_df_is_ws_11 <= io_in_r_bypass_18_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_1_stall_11 <= io_in_r_bypass_18_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_2_data_11 <= io_in_r_bypass_18_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_2_load_store_11 <= io_in_r_bypass_18_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_2_df_is_ws_11 <= io_in_r_bypass_18_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_2_stall_11 <= io_in_r_bypass_18_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_3_data_11 <= io_in_r_bypass_18_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_3_load_store_11 <= io_in_r_bypass_18_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_3_df_is_ws_11 <= io_in_r_bypass_18_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_3_stall_11 <= io_in_r_bypass_18_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_0_data_11 <= io_in_r_bypass_19_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_0_load_store_11 <= io_in_r_bypass_19_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_0_df_is_ws_11 <= io_in_r_bypass_19_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_0_stall_11 <= io_in_r_bypass_19_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_1_data_11 <= io_in_r_bypass_19_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_1_load_store_11 <= io_in_r_bypass_19_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_1_df_is_ws_11 <= io_in_r_bypass_19_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_1_stall_11 <= io_in_r_bypass_19_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_2_data_11 <= io_in_r_bypass_19_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_2_load_store_11 <= io_in_r_bypass_19_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_2_df_is_ws_11 <= io_in_r_bypass_19_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_2_stall_11 <= io_in_r_bypass_19_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_3_data_11 <= io_in_r_bypass_19_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_3_load_store_11 <= io_in_r_bypass_19_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_3_df_is_ws_11 <= io_in_r_bypass_19_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_3_stall_11 <= io_in_r_bypass_19_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_0_data_11 <= io_in_r_bypass_20_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_0_load_store_11 <= io_in_r_bypass_20_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_0_df_is_ws_11 <= io_in_r_bypass_20_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_0_stall_11 <= io_in_r_bypass_20_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_1_data_11 <= io_in_r_bypass_20_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_1_load_store_11 <= io_in_r_bypass_20_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_1_df_is_ws_11 <= io_in_r_bypass_20_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_1_stall_11 <= io_in_r_bypass_20_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_2_data_11 <= io_in_r_bypass_20_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_2_load_store_11 <= io_in_r_bypass_20_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_2_df_is_ws_11 <= io_in_r_bypass_20_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_2_stall_11 <= io_in_r_bypass_20_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_3_data_11 <= io_in_r_bypass_20_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_3_load_store_11 <= io_in_r_bypass_20_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_3_df_is_ws_11 <= io_in_r_bypass_20_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_3_stall_11 <= io_in_r_bypass_20_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_0_data_11 <= io_in_r_bypass_21_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_0_load_store_11 <= io_in_r_bypass_21_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_0_df_is_ws_11 <= io_in_r_bypass_21_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_0_stall_11 <= io_in_r_bypass_21_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_1_data_11 <= io_in_r_bypass_21_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_1_load_store_11 <= io_in_r_bypass_21_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_1_df_is_ws_11 <= io_in_r_bypass_21_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_1_stall_11 <= io_in_r_bypass_21_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_2_data_11 <= io_in_r_bypass_21_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_2_load_store_11 <= io_in_r_bypass_21_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_2_df_is_ws_11 <= io_in_r_bypass_21_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_2_stall_11 <= io_in_r_bypass_21_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_3_data_11 <= io_in_r_bypass_21_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_3_load_store_11 <= io_in_r_bypass_21_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_3_df_is_ws_11 <= io_in_r_bypass_21_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_3_stall_11 <= io_in_r_bypass_21_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_0_data_11 <= io_in_r_bypass_22_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_0_load_store_11 <= io_in_r_bypass_22_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_0_df_is_ws_11 <= io_in_r_bypass_22_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_0_stall_11 <= io_in_r_bypass_22_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_1_data_11 <= io_in_r_bypass_22_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_1_load_store_11 <= io_in_r_bypass_22_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_1_df_is_ws_11 <= io_in_r_bypass_22_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_1_stall_11 <= io_in_r_bypass_22_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_2_data_11 <= io_in_r_bypass_22_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_2_load_store_11 <= io_in_r_bypass_22_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_2_df_is_ws_11 <= io_in_r_bypass_22_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_2_stall_11 <= io_in_r_bypass_22_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_3_data_11 <= io_in_r_bypass_22_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_3_load_store_11 <= io_in_r_bypass_22_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_3_df_is_ws_11 <= io_in_r_bypass_22_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_3_stall_11 <= io_in_r_bypass_22_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_0_data_11 <= io_in_r_bypass_23_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_0_load_store_11 <= io_in_r_bypass_23_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_0_df_is_ws_11 <= io_in_r_bypass_23_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_0_stall_11 <= io_in_r_bypass_23_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_1_data_11 <= io_in_r_bypass_23_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_1_load_store_11 <= io_in_r_bypass_23_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_1_df_is_ws_11 <= io_in_r_bypass_23_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_1_stall_11 <= io_in_r_bypass_23_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_2_data_11 <= io_in_r_bypass_23_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_2_load_store_11 <= io_in_r_bypass_23_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_2_df_is_ws_11 <= io_in_r_bypass_23_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_2_stall_11 <= io_in_r_bypass_23_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_3_data_11 <= io_in_r_bypass_23_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_3_load_store_11 <= io_in_r_bypass_23_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_3_df_is_ws_11 <= io_in_r_bypass_23_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_3_stall_11 <= io_in_r_bypass_23_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_0_data_11 <= io_in_r_bypass_24_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_0_load_store_11 <= io_in_r_bypass_24_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_0_df_is_ws_11 <= io_in_r_bypass_24_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_0_stall_11 <= io_in_r_bypass_24_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_1_data_11 <= io_in_r_bypass_24_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_1_load_store_11 <= io_in_r_bypass_24_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_1_df_is_ws_11 <= io_in_r_bypass_24_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_1_stall_11 <= io_in_r_bypass_24_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_2_data_11 <= io_in_r_bypass_24_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_2_load_store_11 <= io_in_r_bypass_24_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_2_df_is_ws_11 <= io_in_r_bypass_24_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_2_stall_11 <= io_in_r_bypass_24_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_3_data_11 <= io_in_r_bypass_24_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_3_load_store_11 <= io_in_r_bypass_24_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_3_df_is_ws_11 <= io_in_r_bypass_24_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_3_stall_11 <= io_in_r_bypass_24_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_0_data_11 <= io_in_r_bypass_25_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_0_load_store_11 <= io_in_r_bypass_25_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_0_df_is_ws_11 <= io_in_r_bypass_25_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_0_stall_11 <= io_in_r_bypass_25_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_1_data_11 <= io_in_r_bypass_25_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_1_load_store_11 <= io_in_r_bypass_25_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_1_df_is_ws_11 <= io_in_r_bypass_25_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_1_stall_11 <= io_in_r_bypass_25_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_2_data_11 <= io_in_r_bypass_25_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_2_load_store_11 <= io_in_r_bypass_25_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_2_df_is_ws_11 <= io_in_r_bypass_25_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_2_stall_11 <= io_in_r_bypass_25_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_3_data_11 <= io_in_r_bypass_25_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_3_load_store_11 <= io_in_r_bypass_25_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_3_df_is_ws_11 <= io_in_r_bypass_25_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_3_stall_11 <= io_in_r_bypass_25_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_0_data_11 <= io_in_r_bypass_26_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_0_load_store_11 <= io_in_r_bypass_26_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_0_df_is_ws_11 <= io_in_r_bypass_26_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_0_stall_11 <= io_in_r_bypass_26_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_1_data_11 <= io_in_r_bypass_26_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_1_load_store_11 <= io_in_r_bypass_26_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_1_df_is_ws_11 <= io_in_r_bypass_26_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_1_stall_11 <= io_in_r_bypass_26_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_2_data_11 <= io_in_r_bypass_26_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_2_load_store_11 <= io_in_r_bypass_26_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_2_df_is_ws_11 <= io_in_r_bypass_26_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_2_stall_11 <= io_in_r_bypass_26_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_3_data_11 <= io_in_r_bypass_26_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_3_load_store_11 <= io_in_r_bypass_26_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_3_df_is_ws_11 <= io_in_r_bypass_26_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_3_stall_11 <= io_in_r_bypass_26_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_0_data_11 <= io_in_r_bypass_27_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_0_load_store_11 <= io_in_r_bypass_27_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_0_df_is_ws_11 <= io_in_r_bypass_27_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_0_stall_11 <= io_in_r_bypass_27_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_1_data_11 <= io_in_r_bypass_27_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_1_load_store_11 <= io_in_r_bypass_27_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_1_df_is_ws_11 <= io_in_r_bypass_27_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_1_stall_11 <= io_in_r_bypass_27_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_2_data_11 <= io_in_r_bypass_27_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_2_load_store_11 <= io_in_r_bypass_27_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_2_df_is_ws_11 <= io_in_r_bypass_27_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_2_stall_11 <= io_in_r_bypass_27_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_3_data_11 <= io_in_r_bypass_27_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_3_load_store_11 <= io_in_r_bypass_27_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_3_df_is_ws_11 <= io_in_r_bypass_27_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_3_stall_11 <= io_in_r_bypass_27_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_0_data_11 <= io_in_r_bypass_28_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_0_load_store_11 <= io_in_r_bypass_28_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_0_df_is_ws_11 <= io_in_r_bypass_28_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_0_stall_11 <= io_in_r_bypass_28_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_1_data_11 <= io_in_r_bypass_28_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_1_load_store_11 <= io_in_r_bypass_28_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_1_df_is_ws_11 <= io_in_r_bypass_28_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_1_stall_11 <= io_in_r_bypass_28_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_2_data_11 <= io_in_r_bypass_28_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_2_load_store_11 <= io_in_r_bypass_28_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_2_df_is_ws_11 <= io_in_r_bypass_28_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_2_stall_11 <= io_in_r_bypass_28_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_3_data_11 <= io_in_r_bypass_28_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_3_load_store_11 <= io_in_r_bypass_28_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_3_df_is_ws_11 <= io_in_r_bypass_28_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_3_stall_11 <= io_in_r_bypass_28_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_0_data_11 <= io_in_r_bypass_29_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_0_load_store_11 <= io_in_r_bypass_29_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_0_df_is_ws_11 <= io_in_r_bypass_29_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_0_stall_11 <= io_in_r_bypass_29_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_1_data_11 <= io_in_r_bypass_29_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_1_load_store_11 <= io_in_r_bypass_29_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_1_df_is_ws_11 <= io_in_r_bypass_29_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_1_stall_11 <= io_in_r_bypass_29_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_2_data_11 <= io_in_r_bypass_29_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_2_load_store_11 <= io_in_r_bypass_29_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_2_df_is_ws_11 <= io_in_r_bypass_29_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_2_stall_11 <= io_in_r_bypass_29_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_3_data_11 <= io_in_r_bypass_29_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_3_load_store_11 <= io_in_r_bypass_29_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_3_df_is_ws_11 <= io_in_r_bypass_29_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_3_stall_11 <= io_in_r_bypass_29_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_0_data_11 <= io_in_r_bypass_30_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_0_load_store_11 <= io_in_r_bypass_30_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_0_df_is_ws_11 <= io_in_r_bypass_30_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_0_stall_11 <= io_in_r_bypass_30_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_1_data_11 <= io_in_r_bypass_30_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_1_load_store_11 <= io_in_r_bypass_30_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_1_df_is_ws_11 <= io_in_r_bypass_30_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_1_stall_11 <= io_in_r_bypass_30_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_2_data_11 <= io_in_r_bypass_30_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_2_load_store_11 <= io_in_r_bypass_30_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_2_df_is_ws_11 <= io_in_r_bypass_30_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_2_stall_11 <= io_in_r_bypass_30_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_3_data_11 <= io_in_r_bypass_30_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_3_load_store_11 <= io_in_r_bypass_30_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_3_df_is_ws_11 <= io_in_r_bypass_30_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_3_stall_11 <= io_in_r_bypass_30_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_0_data_11 <= io_in_r_bypass_31_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_0_load_store_11 <= io_in_r_bypass_31_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_0_df_is_ws_11 <= io_in_r_bypass_31_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_0_stall_11 <= io_in_r_bypass_31_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_1_data_11 <= io_in_r_bypass_31_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_1_load_store_11 <= io_in_r_bypass_31_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_1_df_is_ws_11 <= io_in_r_bypass_31_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_1_stall_11 <= io_in_r_bypass_31_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_2_data_11 <= io_in_r_bypass_31_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_2_load_store_11 <= io_in_r_bypass_31_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_2_df_is_ws_11 <= io_in_r_bypass_31_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_2_stall_11 <= io_in_r_bypass_31_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_3_data_11 <= io_in_r_bypass_31_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_3_load_store_11 <= io_in_r_bypass_31_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_3_df_is_ws_11 <= io_in_r_bypass_31_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_3_stall_11 <= io_in_r_bypass_31_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_0_data_12 <= io_in_r_bypass_0_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_0_load_store_12 <= io_in_r_bypass_0_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_0_df_is_ws_12 <= io_in_r_bypass_0_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_0_stall_12 <= io_in_r_bypass_0_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_1_data_12 <= io_in_r_bypass_0_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_1_load_store_12 <= io_in_r_bypass_0_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_1_df_is_ws_12 <= io_in_r_bypass_0_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_1_stall_12 <= io_in_r_bypass_0_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_2_data_12 <= io_in_r_bypass_0_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_2_load_store_12 <= io_in_r_bypass_0_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_2_df_is_ws_12 <= io_in_r_bypass_0_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_2_stall_12 <= io_in_r_bypass_0_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_3_data_12 <= io_in_r_bypass_0_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_3_load_store_12 <= io_in_r_bypass_0_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_3_df_is_ws_12 <= io_in_r_bypass_0_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_3_stall_12 <= io_in_r_bypass_0_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_0_data_12 <= io_in_r_bypass_1_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_0_load_store_12 <= io_in_r_bypass_1_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_0_df_is_ws_12 <= io_in_r_bypass_1_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_0_stall_12 <= io_in_r_bypass_1_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_1_data_12 <= io_in_r_bypass_1_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_1_load_store_12 <= io_in_r_bypass_1_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_1_df_is_ws_12 <= io_in_r_bypass_1_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_1_stall_12 <= io_in_r_bypass_1_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_2_data_12 <= io_in_r_bypass_1_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_2_load_store_12 <= io_in_r_bypass_1_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_2_df_is_ws_12 <= io_in_r_bypass_1_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_2_stall_12 <= io_in_r_bypass_1_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_3_data_12 <= io_in_r_bypass_1_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_3_load_store_12 <= io_in_r_bypass_1_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_3_df_is_ws_12 <= io_in_r_bypass_1_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_3_stall_12 <= io_in_r_bypass_1_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_0_data_12 <= io_in_r_bypass_2_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_0_load_store_12 <= io_in_r_bypass_2_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_0_df_is_ws_12 <= io_in_r_bypass_2_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_0_stall_12 <= io_in_r_bypass_2_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_1_data_12 <= io_in_r_bypass_2_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_1_load_store_12 <= io_in_r_bypass_2_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_1_df_is_ws_12 <= io_in_r_bypass_2_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_1_stall_12 <= io_in_r_bypass_2_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_2_data_12 <= io_in_r_bypass_2_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_2_load_store_12 <= io_in_r_bypass_2_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_2_df_is_ws_12 <= io_in_r_bypass_2_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_2_stall_12 <= io_in_r_bypass_2_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_3_data_12 <= io_in_r_bypass_2_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_3_load_store_12 <= io_in_r_bypass_2_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_3_df_is_ws_12 <= io_in_r_bypass_2_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_3_stall_12 <= io_in_r_bypass_2_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_0_data_12 <= io_in_r_bypass_3_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_0_load_store_12 <= io_in_r_bypass_3_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_0_df_is_ws_12 <= io_in_r_bypass_3_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_0_stall_12 <= io_in_r_bypass_3_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_1_data_12 <= io_in_r_bypass_3_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_1_load_store_12 <= io_in_r_bypass_3_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_1_df_is_ws_12 <= io_in_r_bypass_3_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_1_stall_12 <= io_in_r_bypass_3_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_2_data_12 <= io_in_r_bypass_3_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_2_load_store_12 <= io_in_r_bypass_3_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_2_df_is_ws_12 <= io_in_r_bypass_3_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_2_stall_12 <= io_in_r_bypass_3_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_3_data_12 <= io_in_r_bypass_3_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_3_load_store_12 <= io_in_r_bypass_3_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_3_df_is_ws_12 <= io_in_r_bypass_3_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_3_stall_12 <= io_in_r_bypass_3_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_0_data_12 <= io_in_r_bypass_4_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_0_load_store_12 <= io_in_r_bypass_4_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_0_df_is_ws_12 <= io_in_r_bypass_4_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_0_stall_12 <= io_in_r_bypass_4_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_1_data_12 <= io_in_r_bypass_4_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_1_load_store_12 <= io_in_r_bypass_4_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_1_df_is_ws_12 <= io_in_r_bypass_4_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_1_stall_12 <= io_in_r_bypass_4_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_2_data_12 <= io_in_r_bypass_4_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_2_load_store_12 <= io_in_r_bypass_4_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_2_df_is_ws_12 <= io_in_r_bypass_4_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_2_stall_12 <= io_in_r_bypass_4_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_3_data_12 <= io_in_r_bypass_4_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_3_load_store_12 <= io_in_r_bypass_4_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_3_df_is_ws_12 <= io_in_r_bypass_4_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_3_stall_12 <= io_in_r_bypass_4_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_0_data_12 <= io_in_r_bypass_5_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_0_load_store_12 <= io_in_r_bypass_5_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_0_df_is_ws_12 <= io_in_r_bypass_5_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_0_stall_12 <= io_in_r_bypass_5_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_1_data_12 <= io_in_r_bypass_5_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_1_load_store_12 <= io_in_r_bypass_5_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_1_df_is_ws_12 <= io_in_r_bypass_5_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_1_stall_12 <= io_in_r_bypass_5_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_2_data_12 <= io_in_r_bypass_5_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_2_load_store_12 <= io_in_r_bypass_5_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_2_df_is_ws_12 <= io_in_r_bypass_5_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_2_stall_12 <= io_in_r_bypass_5_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_3_data_12 <= io_in_r_bypass_5_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_3_load_store_12 <= io_in_r_bypass_5_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_3_df_is_ws_12 <= io_in_r_bypass_5_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_3_stall_12 <= io_in_r_bypass_5_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_0_data_12 <= io_in_r_bypass_6_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_0_load_store_12 <= io_in_r_bypass_6_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_0_df_is_ws_12 <= io_in_r_bypass_6_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_0_stall_12 <= io_in_r_bypass_6_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_1_data_12 <= io_in_r_bypass_6_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_1_load_store_12 <= io_in_r_bypass_6_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_1_df_is_ws_12 <= io_in_r_bypass_6_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_1_stall_12 <= io_in_r_bypass_6_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_2_data_12 <= io_in_r_bypass_6_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_2_load_store_12 <= io_in_r_bypass_6_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_2_df_is_ws_12 <= io_in_r_bypass_6_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_2_stall_12 <= io_in_r_bypass_6_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_3_data_12 <= io_in_r_bypass_6_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_3_load_store_12 <= io_in_r_bypass_6_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_3_df_is_ws_12 <= io_in_r_bypass_6_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_3_stall_12 <= io_in_r_bypass_6_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_0_data_12 <= io_in_r_bypass_7_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_0_load_store_12 <= io_in_r_bypass_7_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_0_df_is_ws_12 <= io_in_r_bypass_7_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_0_stall_12 <= io_in_r_bypass_7_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_1_data_12 <= io_in_r_bypass_7_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_1_load_store_12 <= io_in_r_bypass_7_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_1_df_is_ws_12 <= io_in_r_bypass_7_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_1_stall_12 <= io_in_r_bypass_7_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_2_data_12 <= io_in_r_bypass_7_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_2_load_store_12 <= io_in_r_bypass_7_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_2_df_is_ws_12 <= io_in_r_bypass_7_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_2_stall_12 <= io_in_r_bypass_7_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_3_data_12 <= io_in_r_bypass_7_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_3_load_store_12 <= io_in_r_bypass_7_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_3_df_is_ws_12 <= io_in_r_bypass_7_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_3_stall_12 <= io_in_r_bypass_7_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_0_data_12 <= io_in_r_bypass_8_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_0_load_store_12 <= io_in_r_bypass_8_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_0_df_is_ws_12 <= io_in_r_bypass_8_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_0_stall_12 <= io_in_r_bypass_8_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_1_data_12 <= io_in_r_bypass_8_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_1_load_store_12 <= io_in_r_bypass_8_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_1_df_is_ws_12 <= io_in_r_bypass_8_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_1_stall_12 <= io_in_r_bypass_8_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_2_data_12 <= io_in_r_bypass_8_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_2_load_store_12 <= io_in_r_bypass_8_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_2_df_is_ws_12 <= io_in_r_bypass_8_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_2_stall_12 <= io_in_r_bypass_8_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_3_data_12 <= io_in_r_bypass_8_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_3_load_store_12 <= io_in_r_bypass_8_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_3_df_is_ws_12 <= io_in_r_bypass_8_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_3_stall_12 <= io_in_r_bypass_8_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_0_data_12 <= io_in_r_bypass_9_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_0_load_store_12 <= io_in_r_bypass_9_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_0_df_is_ws_12 <= io_in_r_bypass_9_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_0_stall_12 <= io_in_r_bypass_9_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_1_data_12 <= io_in_r_bypass_9_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_1_load_store_12 <= io_in_r_bypass_9_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_1_df_is_ws_12 <= io_in_r_bypass_9_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_1_stall_12 <= io_in_r_bypass_9_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_2_data_12 <= io_in_r_bypass_9_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_2_load_store_12 <= io_in_r_bypass_9_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_2_df_is_ws_12 <= io_in_r_bypass_9_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_2_stall_12 <= io_in_r_bypass_9_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_3_data_12 <= io_in_r_bypass_9_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_3_load_store_12 <= io_in_r_bypass_9_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_3_df_is_ws_12 <= io_in_r_bypass_9_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_3_stall_12 <= io_in_r_bypass_9_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_0_data_12 <= io_in_r_bypass_10_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_0_load_store_12 <= io_in_r_bypass_10_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_0_df_is_ws_12 <= io_in_r_bypass_10_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_0_stall_12 <= io_in_r_bypass_10_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_1_data_12 <= io_in_r_bypass_10_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_1_load_store_12 <= io_in_r_bypass_10_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_1_df_is_ws_12 <= io_in_r_bypass_10_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_1_stall_12 <= io_in_r_bypass_10_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_2_data_12 <= io_in_r_bypass_10_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_2_load_store_12 <= io_in_r_bypass_10_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_2_df_is_ws_12 <= io_in_r_bypass_10_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_2_stall_12 <= io_in_r_bypass_10_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_3_data_12 <= io_in_r_bypass_10_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_3_load_store_12 <= io_in_r_bypass_10_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_3_df_is_ws_12 <= io_in_r_bypass_10_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_3_stall_12 <= io_in_r_bypass_10_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_0_data_12 <= io_in_r_bypass_11_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_0_load_store_12 <= io_in_r_bypass_11_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_0_df_is_ws_12 <= io_in_r_bypass_11_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_0_stall_12 <= io_in_r_bypass_11_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_1_data_12 <= io_in_r_bypass_11_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_1_load_store_12 <= io_in_r_bypass_11_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_1_df_is_ws_12 <= io_in_r_bypass_11_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_1_stall_12 <= io_in_r_bypass_11_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_2_data_12 <= io_in_r_bypass_11_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_2_load_store_12 <= io_in_r_bypass_11_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_2_df_is_ws_12 <= io_in_r_bypass_11_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_2_stall_12 <= io_in_r_bypass_11_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_3_data_12 <= io_in_r_bypass_11_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_3_load_store_12 <= io_in_r_bypass_11_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_3_df_is_ws_12 <= io_in_r_bypass_11_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_3_stall_12 <= io_in_r_bypass_11_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_0_data_12 <= io_in_r_bypass_12_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_0_load_store_12 <= io_in_r_bypass_12_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_0_df_is_ws_12 <= io_in_r_bypass_12_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_0_stall_12 <= io_in_r_bypass_12_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_1_data_12 <= io_in_r_bypass_12_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_1_load_store_12 <= io_in_r_bypass_12_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_1_df_is_ws_12 <= io_in_r_bypass_12_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_1_stall_12 <= io_in_r_bypass_12_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_2_data_12 <= io_in_r_bypass_12_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_2_load_store_12 <= io_in_r_bypass_12_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_2_df_is_ws_12 <= io_in_r_bypass_12_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_2_stall_12 <= io_in_r_bypass_12_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_3_data_12 <= io_in_r_bypass_12_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_3_load_store_12 <= io_in_r_bypass_12_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_3_df_is_ws_12 <= io_in_r_bypass_12_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_3_stall_12 <= io_in_r_bypass_12_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_0_data_12 <= io_in_r_bypass_13_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_0_load_store_12 <= io_in_r_bypass_13_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_0_df_is_ws_12 <= io_in_r_bypass_13_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_0_stall_12 <= io_in_r_bypass_13_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_1_data_12 <= io_in_r_bypass_13_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_1_load_store_12 <= io_in_r_bypass_13_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_1_df_is_ws_12 <= io_in_r_bypass_13_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_1_stall_12 <= io_in_r_bypass_13_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_2_data_12 <= io_in_r_bypass_13_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_2_load_store_12 <= io_in_r_bypass_13_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_2_df_is_ws_12 <= io_in_r_bypass_13_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_2_stall_12 <= io_in_r_bypass_13_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_3_data_12 <= io_in_r_bypass_13_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_3_load_store_12 <= io_in_r_bypass_13_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_3_df_is_ws_12 <= io_in_r_bypass_13_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_3_stall_12 <= io_in_r_bypass_13_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_0_data_12 <= io_in_r_bypass_14_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_0_load_store_12 <= io_in_r_bypass_14_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_0_df_is_ws_12 <= io_in_r_bypass_14_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_0_stall_12 <= io_in_r_bypass_14_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_1_data_12 <= io_in_r_bypass_14_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_1_load_store_12 <= io_in_r_bypass_14_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_1_df_is_ws_12 <= io_in_r_bypass_14_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_1_stall_12 <= io_in_r_bypass_14_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_2_data_12 <= io_in_r_bypass_14_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_2_load_store_12 <= io_in_r_bypass_14_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_2_df_is_ws_12 <= io_in_r_bypass_14_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_2_stall_12 <= io_in_r_bypass_14_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_3_data_12 <= io_in_r_bypass_14_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_3_load_store_12 <= io_in_r_bypass_14_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_3_df_is_ws_12 <= io_in_r_bypass_14_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_3_stall_12 <= io_in_r_bypass_14_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_0_data_12 <= io_in_r_bypass_15_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_0_load_store_12 <= io_in_r_bypass_15_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_0_df_is_ws_12 <= io_in_r_bypass_15_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_0_stall_12 <= io_in_r_bypass_15_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_1_data_12 <= io_in_r_bypass_15_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_1_load_store_12 <= io_in_r_bypass_15_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_1_df_is_ws_12 <= io_in_r_bypass_15_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_1_stall_12 <= io_in_r_bypass_15_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_2_data_12 <= io_in_r_bypass_15_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_2_load_store_12 <= io_in_r_bypass_15_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_2_df_is_ws_12 <= io_in_r_bypass_15_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_2_stall_12 <= io_in_r_bypass_15_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_3_data_12 <= io_in_r_bypass_15_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_3_load_store_12 <= io_in_r_bypass_15_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_3_df_is_ws_12 <= io_in_r_bypass_15_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_3_stall_12 <= io_in_r_bypass_15_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_0_data_12 <= io_in_r_bypass_16_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_0_load_store_12 <= io_in_r_bypass_16_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_0_df_is_ws_12 <= io_in_r_bypass_16_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_0_stall_12 <= io_in_r_bypass_16_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_1_data_12 <= io_in_r_bypass_16_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_1_load_store_12 <= io_in_r_bypass_16_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_1_df_is_ws_12 <= io_in_r_bypass_16_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_1_stall_12 <= io_in_r_bypass_16_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_2_data_12 <= io_in_r_bypass_16_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_2_load_store_12 <= io_in_r_bypass_16_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_2_df_is_ws_12 <= io_in_r_bypass_16_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_2_stall_12 <= io_in_r_bypass_16_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_3_data_12 <= io_in_r_bypass_16_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_3_load_store_12 <= io_in_r_bypass_16_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_3_df_is_ws_12 <= io_in_r_bypass_16_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_3_stall_12 <= io_in_r_bypass_16_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_0_data_12 <= io_in_r_bypass_17_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_0_load_store_12 <= io_in_r_bypass_17_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_0_df_is_ws_12 <= io_in_r_bypass_17_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_0_stall_12 <= io_in_r_bypass_17_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_1_data_12 <= io_in_r_bypass_17_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_1_load_store_12 <= io_in_r_bypass_17_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_1_df_is_ws_12 <= io_in_r_bypass_17_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_1_stall_12 <= io_in_r_bypass_17_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_2_data_12 <= io_in_r_bypass_17_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_2_load_store_12 <= io_in_r_bypass_17_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_2_df_is_ws_12 <= io_in_r_bypass_17_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_2_stall_12 <= io_in_r_bypass_17_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_3_data_12 <= io_in_r_bypass_17_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_3_load_store_12 <= io_in_r_bypass_17_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_3_df_is_ws_12 <= io_in_r_bypass_17_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_3_stall_12 <= io_in_r_bypass_17_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_0_data_12 <= io_in_r_bypass_18_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_0_load_store_12 <= io_in_r_bypass_18_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_0_df_is_ws_12 <= io_in_r_bypass_18_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_0_stall_12 <= io_in_r_bypass_18_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_1_data_12 <= io_in_r_bypass_18_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_1_load_store_12 <= io_in_r_bypass_18_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_1_df_is_ws_12 <= io_in_r_bypass_18_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_1_stall_12 <= io_in_r_bypass_18_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_2_data_12 <= io_in_r_bypass_18_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_2_load_store_12 <= io_in_r_bypass_18_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_2_df_is_ws_12 <= io_in_r_bypass_18_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_2_stall_12 <= io_in_r_bypass_18_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_3_data_12 <= io_in_r_bypass_18_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_3_load_store_12 <= io_in_r_bypass_18_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_3_df_is_ws_12 <= io_in_r_bypass_18_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_3_stall_12 <= io_in_r_bypass_18_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_0_data_12 <= io_in_r_bypass_19_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_0_load_store_12 <= io_in_r_bypass_19_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_0_df_is_ws_12 <= io_in_r_bypass_19_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_0_stall_12 <= io_in_r_bypass_19_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_1_data_12 <= io_in_r_bypass_19_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_1_load_store_12 <= io_in_r_bypass_19_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_1_df_is_ws_12 <= io_in_r_bypass_19_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_1_stall_12 <= io_in_r_bypass_19_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_2_data_12 <= io_in_r_bypass_19_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_2_load_store_12 <= io_in_r_bypass_19_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_2_df_is_ws_12 <= io_in_r_bypass_19_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_2_stall_12 <= io_in_r_bypass_19_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_3_data_12 <= io_in_r_bypass_19_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_3_load_store_12 <= io_in_r_bypass_19_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_3_df_is_ws_12 <= io_in_r_bypass_19_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_3_stall_12 <= io_in_r_bypass_19_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_0_data_12 <= io_in_r_bypass_20_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_0_load_store_12 <= io_in_r_bypass_20_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_0_df_is_ws_12 <= io_in_r_bypass_20_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_0_stall_12 <= io_in_r_bypass_20_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_1_data_12 <= io_in_r_bypass_20_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_1_load_store_12 <= io_in_r_bypass_20_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_1_df_is_ws_12 <= io_in_r_bypass_20_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_1_stall_12 <= io_in_r_bypass_20_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_2_data_12 <= io_in_r_bypass_20_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_2_load_store_12 <= io_in_r_bypass_20_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_2_df_is_ws_12 <= io_in_r_bypass_20_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_2_stall_12 <= io_in_r_bypass_20_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_3_data_12 <= io_in_r_bypass_20_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_3_load_store_12 <= io_in_r_bypass_20_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_3_df_is_ws_12 <= io_in_r_bypass_20_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_3_stall_12 <= io_in_r_bypass_20_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_0_data_12 <= io_in_r_bypass_21_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_0_load_store_12 <= io_in_r_bypass_21_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_0_df_is_ws_12 <= io_in_r_bypass_21_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_0_stall_12 <= io_in_r_bypass_21_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_1_data_12 <= io_in_r_bypass_21_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_1_load_store_12 <= io_in_r_bypass_21_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_1_df_is_ws_12 <= io_in_r_bypass_21_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_1_stall_12 <= io_in_r_bypass_21_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_2_data_12 <= io_in_r_bypass_21_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_2_load_store_12 <= io_in_r_bypass_21_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_2_df_is_ws_12 <= io_in_r_bypass_21_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_2_stall_12 <= io_in_r_bypass_21_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_3_data_12 <= io_in_r_bypass_21_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_3_load_store_12 <= io_in_r_bypass_21_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_3_df_is_ws_12 <= io_in_r_bypass_21_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_3_stall_12 <= io_in_r_bypass_21_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_0_data_12 <= io_in_r_bypass_22_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_0_load_store_12 <= io_in_r_bypass_22_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_0_df_is_ws_12 <= io_in_r_bypass_22_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_0_stall_12 <= io_in_r_bypass_22_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_1_data_12 <= io_in_r_bypass_22_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_1_load_store_12 <= io_in_r_bypass_22_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_1_df_is_ws_12 <= io_in_r_bypass_22_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_1_stall_12 <= io_in_r_bypass_22_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_2_data_12 <= io_in_r_bypass_22_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_2_load_store_12 <= io_in_r_bypass_22_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_2_df_is_ws_12 <= io_in_r_bypass_22_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_2_stall_12 <= io_in_r_bypass_22_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_3_data_12 <= io_in_r_bypass_22_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_3_load_store_12 <= io_in_r_bypass_22_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_3_df_is_ws_12 <= io_in_r_bypass_22_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_3_stall_12 <= io_in_r_bypass_22_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_0_data_12 <= io_in_r_bypass_23_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_0_load_store_12 <= io_in_r_bypass_23_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_0_df_is_ws_12 <= io_in_r_bypass_23_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_0_stall_12 <= io_in_r_bypass_23_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_1_data_12 <= io_in_r_bypass_23_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_1_load_store_12 <= io_in_r_bypass_23_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_1_df_is_ws_12 <= io_in_r_bypass_23_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_1_stall_12 <= io_in_r_bypass_23_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_2_data_12 <= io_in_r_bypass_23_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_2_load_store_12 <= io_in_r_bypass_23_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_2_df_is_ws_12 <= io_in_r_bypass_23_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_2_stall_12 <= io_in_r_bypass_23_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_3_data_12 <= io_in_r_bypass_23_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_3_load_store_12 <= io_in_r_bypass_23_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_3_df_is_ws_12 <= io_in_r_bypass_23_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_3_stall_12 <= io_in_r_bypass_23_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_0_data_12 <= io_in_r_bypass_24_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_0_load_store_12 <= io_in_r_bypass_24_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_0_df_is_ws_12 <= io_in_r_bypass_24_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_0_stall_12 <= io_in_r_bypass_24_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_1_data_12 <= io_in_r_bypass_24_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_1_load_store_12 <= io_in_r_bypass_24_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_1_df_is_ws_12 <= io_in_r_bypass_24_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_1_stall_12 <= io_in_r_bypass_24_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_2_data_12 <= io_in_r_bypass_24_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_2_load_store_12 <= io_in_r_bypass_24_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_2_df_is_ws_12 <= io_in_r_bypass_24_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_2_stall_12 <= io_in_r_bypass_24_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_3_data_12 <= io_in_r_bypass_24_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_3_load_store_12 <= io_in_r_bypass_24_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_3_df_is_ws_12 <= io_in_r_bypass_24_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_3_stall_12 <= io_in_r_bypass_24_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_0_data_12 <= io_in_r_bypass_25_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_0_load_store_12 <= io_in_r_bypass_25_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_0_df_is_ws_12 <= io_in_r_bypass_25_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_0_stall_12 <= io_in_r_bypass_25_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_1_data_12 <= io_in_r_bypass_25_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_1_load_store_12 <= io_in_r_bypass_25_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_1_df_is_ws_12 <= io_in_r_bypass_25_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_1_stall_12 <= io_in_r_bypass_25_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_2_data_12 <= io_in_r_bypass_25_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_2_load_store_12 <= io_in_r_bypass_25_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_2_df_is_ws_12 <= io_in_r_bypass_25_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_2_stall_12 <= io_in_r_bypass_25_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_3_data_12 <= io_in_r_bypass_25_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_3_load_store_12 <= io_in_r_bypass_25_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_3_df_is_ws_12 <= io_in_r_bypass_25_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_3_stall_12 <= io_in_r_bypass_25_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_0_data_12 <= io_in_r_bypass_26_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_0_load_store_12 <= io_in_r_bypass_26_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_0_df_is_ws_12 <= io_in_r_bypass_26_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_0_stall_12 <= io_in_r_bypass_26_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_1_data_12 <= io_in_r_bypass_26_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_1_load_store_12 <= io_in_r_bypass_26_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_1_df_is_ws_12 <= io_in_r_bypass_26_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_1_stall_12 <= io_in_r_bypass_26_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_2_data_12 <= io_in_r_bypass_26_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_2_load_store_12 <= io_in_r_bypass_26_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_2_df_is_ws_12 <= io_in_r_bypass_26_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_2_stall_12 <= io_in_r_bypass_26_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_3_data_12 <= io_in_r_bypass_26_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_3_load_store_12 <= io_in_r_bypass_26_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_3_df_is_ws_12 <= io_in_r_bypass_26_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_3_stall_12 <= io_in_r_bypass_26_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_0_data_12 <= io_in_r_bypass_27_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_0_load_store_12 <= io_in_r_bypass_27_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_0_df_is_ws_12 <= io_in_r_bypass_27_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_0_stall_12 <= io_in_r_bypass_27_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_1_data_12 <= io_in_r_bypass_27_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_1_load_store_12 <= io_in_r_bypass_27_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_1_df_is_ws_12 <= io_in_r_bypass_27_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_1_stall_12 <= io_in_r_bypass_27_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_2_data_12 <= io_in_r_bypass_27_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_2_load_store_12 <= io_in_r_bypass_27_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_2_df_is_ws_12 <= io_in_r_bypass_27_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_2_stall_12 <= io_in_r_bypass_27_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_3_data_12 <= io_in_r_bypass_27_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_3_load_store_12 <= io_in_r_bypass_27_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_3_df_is_ws_12 <= io_in_r_bypass_27_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_3_stall_12 <= io_in_r_bypass_27_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_0_data_12 <= io_in_r_bypass_28_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_0_load_store_12 <= io_in_r_bypass_28_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_0_df_is_ws_12 <= io_in_r_bypass_28_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_0_stall_12 <= io_in_r_bypass_28_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_1_data_12 <= io_in_r_bypass_28_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_1_load_store_12 <= io_in_r_bypass_28_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_1_df_is_ws_12 <= io_in_r_bypass_28_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_1_stall_12 <= io_in_r_bypass_28_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_2_data_12 <= io_in_r_bypass_28_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_2_load_store_12 <= io_in_r_bypass_28_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_2_df_is_ws_12 <= io_in_r_bypass_28_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_2_stall_12 <= io_in_r_bypass_28_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_3_data_12 <= io_in_r_bypass_28_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_3_load_store_12 <= io_in_r_bypass_28_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_3_df_is_ws_12 <= io_in_r_bypass_28_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_3_stall_12 <= io_in_r_bypass_28_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_0_data_12 <= io_in_r_bypass_29_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_0_load_store_12 <= io_in_r_bypass_29_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_0_df_is_ws_12 <= io_in_r_bypass_29_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_0_stall_12 <= io_in_r_bypass_29_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_1_data_12 <= io_in_r_bypass_29_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_1_load_store_12 <= io_in_r_bypass_29_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_1_df_is_ws_12 <= io_in_r_bypass_29_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_1_stall_12 <= io_in_r_bypass_29_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_2_data_12 <= io_in_r_bypass_29_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_2_load_store_12 <= io_in_r_bypass_29_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_2_df_is_ws_12 <= io_in_r_bypass_29_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_2_stall_12 <= io_in_r_bypass_29_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_3_data_12 <= io_in_r_bypass_29_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_3_load_store_12 <= io_in_r_bypass_29_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_3_df_is_ws_12 <= io_in_r_bypass_29_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_3_stall_12 <= io_in_r_bypass_29_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_0_data_12 <= io_in_r_bypass_30_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_0_load_store_12 <= io_in_r_bypass_30_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_0_df_is_ws_12 <= io_in_r_bypass_30_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_0_stall_12 <= io_in_r_bypass_30_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_1_data_12 <= io_in_r_bypass_30_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_1_load_store_12 <= io_in_r_bypass_30_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_1_df_is_ws_12 <= io_in_r_bypass_30_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_1_stall_12 <= io_in_r_bypass_30_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_2_data_12 <= io_in_r_bypass_30_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_2_load_store_12 <= io_in_r_bypass_30_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_2_df_is_ws_12 <= io_in_r_bypass_30_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_2_stall_12 <= io_in_r_bypass_30_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_3_data_12 <= io_in_r_bypass_30_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_3_load_store_12 <= io_in_r_bypass_30_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_3_df_is_ws_12 <= io_in_r_bypass_30_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_3_stall_12 <= io_in_r_bypass_30_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_0_data_12 <= io_in_r_bypass_31_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_0_load_store_12 <= io_in_r_bypass_31_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_0_df_is_ws_12 <= io_in_r_bypass_31_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_0_stall_12 <= io_in_r_bypass_31_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_1_data_12 <= io_in_r_bypass_31_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_1_load_store_12 <= io_in_r_bypass_31_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_1_df_is_ws_12 <= io_in_r_bypass_31_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_1_stall_12 <= io_in_r_bypass_31_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_2_data_12 <= io_in_r_bypass_31_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_2_load_store_12 <= io_in_r_bypass_31_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_2_df_is_ws_12 <= io_in_r_bypass_31_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_2_stall_12 <= io_in_r_bypass_31_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_3_data_12 <= io_in_r_bypass_31_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_3_load_store_12 <= io_in_r_bypass_31_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_3_df_is_ws_12 <= io_in_r_bypass_31_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_3_stall_12 <= io_in_r_bypass_31_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_0_data_13 <= io_in_r_bypass_0_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_0_load_store_13 <= io_in_r_bypass_0_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_0_df_is_ws_13 <= io_in_r_bypass_0_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_0_stall_13 <= io_in_r_bypass_0_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_1_data_13 <= io_in_r_bypass_0_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_1_load_store_13 <= io_in_r_bypass_0_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_1_df_is_ws_13 <= io_in_r_bypass_0_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_1_stall_13 <= io_in_r_bypass_0_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_2_data_13 <= io_in_r_bypass_0_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_2_load_store_13 <= io_in_r_bypass_0_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_2_df_is_ws_13 <= io_in_r_bypass_0_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_2_stall_13 <= io_in_r_bypass_0_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_3_data_13 <= io_in_r_bypass_0_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_3_load_store_13 <= io_in_r_bypass_0_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_3_df_is_ws_13 <= io_in_r_bypass_0_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_3_stall_13 <= io_in_r_bypass_0_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_0_data_13 <= io_in_r_bypass_1_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_0_load_store_13 <= io_in_r_bypass_1_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_0_df_is_ws_13 <= io_in_r_bypass_1_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_0_stall_13 <= io_in_r_bypass_1_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_1_data_13 <= io_in_r_bypass_1_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_1_load_store_13 <= io_in_r_bypass_1_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_1_df_is_ws_13 <= io_in_r_bypass_1_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_1_stall_13 <= io_in_r_bypass_1_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_2_data_13 <= io_in_r_bypass_1_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_2_load_store_13 <= io_in_r_bypass_1_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_2_df_is_ws_13 <= io_in_r_bypass_1_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_2_stall_13 <= io_in_r_bypass_1_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_3_data_13 <= io_in_r_bypass_1_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_3_load_store_13 <= io_in_r_bypass_1_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_3_df_is_ws_13 <= io_in_r_bypass_1_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_3_stall_13 <= io_in_r_bypass_1_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_0_data_13 <= io_in_r_bypass_2_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_0_load_store_13 <= io_in_r_bypass_2_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_0_df_is_ws_13 <= io_in_r_bypass_2_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_0_stall_13 <= io_in_r_bypass_2_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_1_data_13 <= io_in_r_bypass_2_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_1_load_store_13 <= io_in_r_bypass_2_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_1_df_is_ws_13 <= io_in_r_bypass_2_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_1_stall_13 <= io_in_r_bypass_2_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_2_data_13 <= io_in_r_bypass_2_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_2_load_store_13 <= io_in_r_bypass_2_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_2_df_is_ws_13 <= io_in_r_bypass_2_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_2_stall_13 <= io_in_r_bypass_2_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_3_data_13 <= io_in_r_bypass_2_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_3_load_store_13 <= io_in_r_bypass_2_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_3_df_is_ws_13 <= io_in_r_bypass_2_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_3_stall_13 <= io_in_r_bypass_2_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_0_data_13 <= io_in_r_bypass_3_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_0_load_store_13 <= io_in_r_bypass_3_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_0_df_is_ws_13 <= io_in_r_bypass_3_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_0_stall_13 <= io_in_r_bypass_3_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_1_data_13 <= io_in_r_bypass_3_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_1_load_store_13 <= io_in_r_bypass_3_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_1_df_is_ws_13 <= io_in_r_bypass_3_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_1_stall_13 <= io_in_r_bypass_3_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_2_data_13 <= io_in_r_bypass_3_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_2_load_store_13 <= io_in_r_bypass_3_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_2_df_is_ws_13 <= io_in_r_bypass_3_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_2_stall_13 <= io_in_r_bypass_3_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_3_data_13 <= io_in_r_bypass_3_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_3_load_store_13 <= io_in_r_bypass_3_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_3_df_is_ws_13 <= io_in_r_bypass_3_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_3_stall_13 <= io_in_r_bypass_3_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_0_data_13 <= io_in_r_bypass_4_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_0_load_store_13 <= io_in_r_bypass_4_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_0_df_is_ws_13 <= io_in_r_bypass_4_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_0_stall_13 <= io_in_r_bypass_4_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_1_data_13 <= io_in_r_bypass_4_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_1_load_store_13 <= io_in_r_bypass_4_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_1_df_is_ws_13 <= io_in_r_bypass_4_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_1_stall_13 <= io_in_r_bypass_4_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_2_data_13 <= io_in_r_bypass_4_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_2_load_store_13 <= io_in_r_bypass_4_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_2_df_is_ws_13 <= io_in_r_bypass_4_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_2_stall_13 <= io_in_r_bypass_4_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_3_data_13 <= io_in_r_bypass_4_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_3_load_store_13 <= io_in_r_bypass_4_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_3_df_is_ws_13 <= io_in_r_bypass_4_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_3_stall_13 <= io_in_r_bypass_4_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_0_data_13 <= io_in_r_bypass_5_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_0_load_store_13 <= io_in_r_bypass_5_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_0_df_is_ws_13 <= io_in_r_bypass_5_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_0_stall_13 <= io_in_r_bypass_5_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_1_data_13 <= io_in_r_bypass_5_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_1_load_store_13 <= io_in_r_bypass_5_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_1_df_is_ws_13 <= io_in_r_bypass_5_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_1_stall_13 <= io_in_r_bypass_5_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_2_data_13 <= io_in_r_bypass_5_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_2_load_store_13 <= io_in_r_bypass_5_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_2_df_is_ws_13 <= io_in_r_bypass_5_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_2_stall_13 <= io_in_r_bypass_5_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_3_data_13 <= io_in_r_bypass_5_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_3_load_store_13 <= io_in_r_bypass_5_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_3_df_is_ws_13 <= io_in_r_bypass_5_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_3_stall_13 <= io_in_r_bypass_5_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_0_data_13 <= io_in_r_bypass_6_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_0_load_store_13 <= io_in_r_bypass_6_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_0_df_is_ws_13 <= io_in_r_bypass_6_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_0_stall_13 <= io_in_r_bypass_6_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_1_data_13 <= io_in_r_bypass_6_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_1_load_store_13 <= io_in_r_bypass_6_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_1_df_is_ws_13 <= io_in_r_bypass_6_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_1_stall_13 <= io_in_r_bypass_6_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_2_data_13 <= io_in_r_bypass_6_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_2_load_store_13 <= io_in_r_bypass_6_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_2_df_is_ws_13 <= io_in_r_bypass_6_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_2_stall_13 <= io_in_r_bypass_6_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_3_data_13 <= io_in_r_bypass_6_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_3_load_store_13 <= io_in_r_bypass_6_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_3_df_is_ws_13 <= io_in_r_bypass_6_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_3_stall_13 <= io_in_r_bypass_6_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_0_data_13 <= io_in_r_bypass_7_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_0_load_store_13 <= io_in_r_bypass_7_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_0_df_is_ws_13 <= io_in_r_bypass_7_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_0_stall_13 <= io_in_r_bypass_7_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_1_data_13 <= io_in_r_bypass_7_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_1_load_store_13 <= io_in_r_bypass_7_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_1_df_is_ws_13 <= io_in_r_bypass_7_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_1_stall_13 <= io_in_r_bypass_7_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_2_data_13 <= io_in_r_bypass_7_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_2_load_store_13 <= io_in_r_bypass_7_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_2_df_is_ws_13 <= io_in_r_bypass_7_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_2_stall_13 <= io_in_r_bypass_7_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_3_data_13 <= io_in_r_bypass_7_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_3_load_store_13 <= io_in_r_bypass_7_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_3_df_is_ws_13 <= io_in_r_bypass_7_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_3_stall_13 <= io_in_r_bypass_7_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_0_data_13 <= io_in_r_bypass_8_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_0_load_store_13 <= io_in_r_bypass_8_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_0_df_is_ws_13 <= io_in_r_bypass_8_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_0_stall_13 <= io_in_r_bypass_8_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_1_data_13 <= io_in_r_bypass_8_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_1_load_store_13 <= io_in_r_bypass_8_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_1_df_is_ws_13 <= io_in_r_bypass_8_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_1_stall_13 <= io_in_r_bypass_8_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_2_data_13 <= io_in_r_bypass_8_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_2_load_store_13 <= io_in_r_bypass_8_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_2_df_is_ws_13 <= io_in_r_bypass_8_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_2_stall_13 <= io_in_r_bypass_8_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_3_data_13 <= io_in_r_bypass_8_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_3_load_store_13 <= io_in_r_bypass_8_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_3_df_is_ws_13 <= io_in_r_bypass_8_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_3_stall_13 <= io_in_r_bypass_8_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_0_data_13 <= io_in_r_bypass_9_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_0_load_store_13 <= io_in_r_bypass_9_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_0_df_is_ws_13 <= io_in_r_bypass_9_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_0_stall_13 <= io_in_r_bypass_9_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_1_data_13 <= io_in_r_bypass_9_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_1_load_store_13 <= io_in_r_bypass_9_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_1_df_is_ws_13 <= io_in_r_bypass_9_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_1_stall_13 <= io_in_r_bypass_9_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_2_data_13 <= io_in_r_bypass_9_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_2_load_store_13 <= io_in_r_bypass_9_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_2_df_is_ws_13 <= io_in_r_bypass_9_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_2_stall_13 <= io_in_r_bypass_9_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_3_data_13 <= io_in_r_bypass_9_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_3_load_store_13 <= io_in_r_bypass_9_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_3_df_is_ws_13 <= io_in_r_bypass_9_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_3_stall_13 <= io_in_r_bypass_9_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_0_data_13 <= io_in_r_bypass_10_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_0_load_store_13 <= io_in_r_bypass_10_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_0_df_is_ws_13 <= io_in_r_bypass_10_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_0_stall_13 <= io_in_r_bypass_10_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_1_data_13 <= io_in_r_bypass_10_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_1_load_store_13 <= io_in_r_bypass_10_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_1_df_is_ws_13 <= io_in_r_bypass_10_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_1_stall_13 <= io_in_r_bypass_10_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_2_data_13 <= io_in_r_bypass_10_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_2_load_store_13 <= io_in_r_bypass_10_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_2_df_is_ws_13 <= io_in_r_bypass_10_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_2_stall_13 <= io_in_r_bypass_10_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_3_data_13 <= io_in_r_bypass_10_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_3_load_store_13 <= io_in_r_bypass_10_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_3_df_is_ws_13 <= io_in_r_bypass_10_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_3_stall_13 <= io_in_r_bypass_10_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_0_data_13 <= io_in_r_bypass_11_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_0_load_store_13 <= io_in_r_bypass_11_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_0_df_is_ws_13 <= io_in_r_bypass_11_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_0_stall_13 <= io_in_r_bypass_11_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_1_data_13 <= io_in_r_bypass_11_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_1_load_store_13 <= io_in_r_bypass_11_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_1_df_is_ws_13 <= io_in_r_bypass_11_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_1_stall_13 <= io_in_r_bypass_11_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_2_data_13 <= io_in_r_bypass_11_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_2_load_store_13 <= io_in_r_bypass_11_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_2_df_is_ws_13 <= io_in_r_bypass_11_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_2_stall_13 <= io_in_r_bypass_11_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_3_data_13 <= io_in_r_bypass_11_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_3_load_store_13 <= io_in_r_bypass_11_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_3_df_is_ws_13 <= io_in_r_bypass_11_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_3_stall_13 <= io_in_r_bypass_11_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_0_data_13 <= io_in_r_bypass_12_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_0_load_store_13 <= io_in_r_bypass_12_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_0_df_is_ws_13 <= io_in_r_bypass_12_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_0_stall_13 <= io_in_r_bypass_12_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_1_data_13 <= io_in_r_bypass_12_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_1_load_store_13 <= io_in_r_bypass_12_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_1_df_is_ws_13 <= io_in_r_bypass_12_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_1_stall_13 <= io_in_r_bypass_12_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_2_data_13 <= io_in_r_bypass_12_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_2_load_store_13 <= io_in_r_bypass_12_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_2_df_is_ws_13 <= io_in_r_bypass_12_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_2_stall_13 <= io_in_r_bypass_12_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_3_data_13 <= io_in_r_bypass_12_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_3_load_store_13 <= io_in_r_bypass_12_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_3_df_is_ws_13 <= io_in_r_bypass_12_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_3_stall_13 <= io_in_r_bypass_12_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_0_data_13 <= io_in_r_bypass_13_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_0_load_store_13 <= io_in_r_bypass_13_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_0_df_is_ws_13 <= io_in_r_bypass_13_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_0_stall_13 <= io_in_r_bypass_13_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_1_data_13 <= io_in_r_bypass_13_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_1_load_store_13 <= io_in_r_bypass_13_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_1_df_is_ws_13 <= io_in_r_bypass_13_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_1_stall_13 <= io_in_r_bypass_13_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_2_data_13 <= io_in_r_bypass_13_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_2_load_store_13 <= io_in_r_bypass_13_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_2_df_is_ws_13 <= io_in_r_bypass_13_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_2_stall_13 <= io_in_r_bypass_13_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_3_data_13 <= io_in_r_bypass_13_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_3_load_store_13 <= io_in_r_bypass_13_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_3_df_is_ws_13 <= io_in_r_bypass_13_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_3_stall_13 <= io_in_r_bypass_13_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_0_data_13 <= io_in_r_bypass_14_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_0_load_store_13 <= io_in_r_bypass_14_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_0_df_is_ws_13 <= io_in_r_bypass_14_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_0_stall_13 <= io_in_r_bypass_14_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_1_data_13 <= io_in_r_bypass_14_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_1_load_store_13 <= io_in_r_bypass_14_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_1_df_is_ws_13 <= io_in_r_bypass_14_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_1_stall_13 <= io_in_r_bypass_14_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_2_data_13 <= io_in_r_bypass_14_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_2_load_store_13 <= io_in_r_bypass_14_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_2_df_is_ws_13 <= io_in_r_bypass_14_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_2_stall_13 <= io_in_r_bypass_14_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_3_data_13 <= io_in_r_bypass_14_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_3_load_store_13 <= io_in_r_bypass_14_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_3_df_is_ws_13 <= io_in_r_bypass_14_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_3_stall_13 <= io_in_r_bypass_14_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_0_data_13 <= io_in_r_bypass_15_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_0_load_store_13 <= io_in_r_bypass_15_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_0_df_is_ws_13 <= io_in_r_bypass_15_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_0_stall_13 <= io_in_r_bypass_15_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_1_data_13 <= io_in_r_bypass_15_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_1_load_store_13 <= io_in_r_bypass_15_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_1_df_is_ws_13 <= io_in_r_bypass_15_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_1_stall_13 <= io_in_r_bypass_15_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_2_data_13 <= io_in_r_bypass_15_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_2_load_store_13 <= io_in_r_bypass_15_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_2_df_is_ws_13 <= io_in_r_bypass_15_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_2_stall_13 <= io_in_r_bypass_15_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_3_data_13 <= io_in_r_bypass_15_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_3_load_store_13 <= io_in_r_bypass_15_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_3_df_is_ws_13 <= io_in_r_bypass_15_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_3_stall_13 <= io_in_r_bypass_15_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_0_data_13 <= io_in_r_bypass_16_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_0_load_store_13 <= io_in_r_bypass_16_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_0_df_is_ws_13 <= io_in_r_bypass_16_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_0_stall_13 <= io_in_r_bypass_16_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_1_data_13 <= io_in_r_bypass_16_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_1_load_store_13 <= io_in_r_bypass_16_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_1_df_is_ws_13 <= io_in_r_bypass_16_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_1_stall_13 <= io_in_r_bypass_16_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_2_data_13 <= io_in_r_bypass_16_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_2_load_store_13 <= io_in_r_bypass_16_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_2_df_is_ws_13 <= io_in_r_bypass_16_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_2_stall_13 <= io_in_r_bypass_16_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_3_data_13 <= io_in_r_bypass_16_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_3_load_store_13 <= io_in_r_bypass_16_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_3_df_is_ws_13 <= io_in_r_bypass_16_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_3_stall_13 <= io_in_r_bypass_16_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_0_data_13 <= io_in_r_bypass_17_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_0_load_store_13 <= io_in_r_bypass_17_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_0_df_is_ws_13 <= io_in_r_bypass_17_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_0_stall_13 <= io_in_r_bypass_17_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_1_data_13 <= io_in_r_bypass_17_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_1_load_store_13 <= io_in_r_bypass_17_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_1_df_is_ws_13 <= io_in_r_bypass_17_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_1_stall_13 <= io_in_r_bypass_17_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_2_data_13 <= io_in_r_bypass_17_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_2_load_store_13 <= io_in_r_bypass_17_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_2_df_is_ws_13 <= io_in_r_bypass_17_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_2_stall_13 <= io_in_r_bypass_17_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_3_data_13 <= io_in_r_bypass_17_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_3_load_store_13 <= io_in_r_bypass_17_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_3_df_is_ws_13 <= io_in_r_bypass_17_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_3_stall_13 <= io_in_r_bypass_17_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_0_data_13 <= io_in_r_bypass_18_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_0_load_store_13 <= io_in_r_bypass_18_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_0_df_is_ws_13 <= io_in_r_bypass_18_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_0_stall_13 <= io_in_r_bypass_18_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_1_data_13 <= io_in_r_bypass_18_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_1_load_store_13 <= io_in_r_bypass_18_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_1_df_is_ws_13 <= io_in_r_bypass_18_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_1_stall_13 <= io_in_r_bypass_18_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_2_data_13 <= io_in_r_bypass_18_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_2_load_store_13 <= io_in_r_bypass_18_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_2_df_is_ws_13 <= io_in_r_bypass_18_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_2_stall_13 <= io_in_r_bypass_18_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_3_data_13 <= io_in_r_bypass_18_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_3_load_store_13 <= io_in_r_bypass_18_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_3_df_is_ws_13 <= io_in_r_bypass_18_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_3_stall_13 <= io_in_r_bypass_18_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_0_data_13 <= io_in_r_bypass_19_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_0_load_store_13 <= io_in_r_bypass_19_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_0_df_is_ws_13 <= io_in_r_bypass_19_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_0_stall_13 <= io_in_r_bypass_19_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_1_data_13 <= io_in_r_bypass_19_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_1_load_store_13 <= io_in_r_bypass_19_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_1_df_is_ws_13 <= io_in_r_bypass_19_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_1_stall_13 <= io_in_r_bypass_19_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_2_data_13 <= io_in_r_bypass_19_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_2_load_store_13 <= io_in_r_bypass_19_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_2_df_is_ws_13 <= io_in_r_bypass_19_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_2_stall_13 <= io_in_r_bypass_19_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_3_data_13 <= io_in_r_bypass_19_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_3_load_store_13 <= io_in_r_bypass_19_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_3_df_is_ws_13 <= io_in_r_bypass_19_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_3_stall_13 <= io_in_r_bypass_19_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_0_data_13 <= io_in_r_bypass_20_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_0_load_store_13 <= io_in_r_bypass_20_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_0_df_is_ws_13 <= io_in_r_bypass_20_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_0_stall_13 <= io_in_r_bypass_20_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_1_data_13 <= io_in_r_bypass_20_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_1_load_store_13 <= io_in_r_bypass_20_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_1_df_is_ws_13 <= io_in_r_bypass_20_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_1_stall_13 <= io_in_r_bypass_20_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_2_data_13 <= io_in_r_bypass_20_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_2_load_store_13 <= io_in_r_bypass_20_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_2_df_is_ws_13 <= io_in_r_bypass_20_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_2_stall_13 <= io_in_r_bypass_20_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_3_data_13 <= io_in_r_bypass_20_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_3_load_store_13 <= io_in_r_bypass_20_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_3_df_is_ws_13 <= io_in_r_bypass_20_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_3_stall_13 <= io_in_r_bypass_20_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_0_data_13 <= io_in_r_bypass_21_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_0_load_store_13 <= io_in_r_bypass_21_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_0_df_is_ws_13 <= io_in_r_bypass_21_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_0_stall_13 <= io_in_r_bypass_21_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_1_data_13 <= io_in_r_bypass_21_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_1_load_store_13 <= io_in_r_bypass_21_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_1_df_is_ws_13 <= io_in_r_bypass_21_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_1_stall_13 <= io_in_r_bypass_21_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_2_data_13 <= io_in_r_bypass_21_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_2_load_store_13 <= io_in_r_bypass_21_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_2_df_is_ws_13 <= io_in_r_bypass_21_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_2_stall_13 <= io_in_r_bypass_21_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_3_data_13 <= io_in_r_bypass_21_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_3_load_store_13 <= io_in_r_bypass_21_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_3_df_is_ws_13 <= io_in_r_bypass_21_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_3_stall_13 <= io_in_r_bypass_21_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_0_data_13 <= io_in_r_bypass_22_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_0_load_store_13 <= io_in_r_bypass_22_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_0_df_is_ws_13 <= io_in_r_bypass_22_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_0_stall_13 <= io_in_r_bypass_22_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_1_data_13 <= io_in_r_bypass_22_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_1_load_store_13 <= io_in_r_bypass_22_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_1_df_is_ws_13 <= io_in_r_bypass_22_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_1_stall_13 <= io_in_r_bypass_22_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_2_data_13 <= io_in_r_bypass_22_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_2_load_store_13 <= io_in_r_bypass_22_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_2_df_is_ws_13 <= io_in_r_bypass_22_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_2_stall_13 <= io_in_r_bypass_22_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_3_data_13 <= io_in_r_bypass_22_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_3_load_store_13 <= io_in_r_bypass_22_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_3_df_is_ws_13 <= io_in_r_bypass_22_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_3_stall_13 <= io_in_r_bypass_22_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_0_data_13 <= io_in_r_bypass_23_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_0_load_store_13 <= io_in_r_bypass_23_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_0_df_is_ws_13 <= io_in_r_bypass_23_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_0_stall_13 <= io_in_r_bypass_23_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_1_data_13 <= io_in_r_bypass_23_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_1_load_store_13 <= io_in_r_bypass_23_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_1_df_is_ws_13 <= io_in_r_bypass_23_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_1_stall_13 <= io_in_r_bypass_23_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_2_data_13 <= io_in_r_bypass_23_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_2_load_store_13 <= io_in_r_bypass_23_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_2_df_is_ws_13 <= io_in_r_bypass_23_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_2_stall_13 <= io_in_r_bypass_23_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_3_data_13 <= io_in_r_bypass_23_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_3_load_store_13 <= io_in_r_bypass_23_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_3_df_is_ws_13 <= io_in_r_bypass_23_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_3_stall_13 <= io_in_r_bypass_23_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_0_data_13 <= io_in_r_bypass_24_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_0_load_store_13 <= io_in_r_bypass_24_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_0_df_is_ws_13 <= io_in_r_bypass_24_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_0_stall_13 <= io_in_r_bypass_24_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_1_data_13 <= io_in_r_bypass_24_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_1_load_store_13 <= io_in_r_bypass_24_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_1_df_is_ws_13 <= io_in_r_bypass_24_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_1_stall_13 <= io_in_r_bypass_24_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_2_data_13 <= io_in_r_bypass_24_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_2_load_store_13 <= io_in_r_bypass_24_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_2_df_is_ws_13 <= io_in_r_bypass_24_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_2_stall_13 <= io_in_r_bypass_24_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_3_data_13 <= io_in_r_bypass_24_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_3_load_store_13 <= io_in_r_bypass_24_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_3_df_is_ws_13 <= io_in_r_bypass_24_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_3_stall_13 <= io_in_r_bypass_24_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_0_data_13 <= io_in_r_bypass_25_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_0_load_store_13 <= io_in_r_bypass_25_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_0_df_is_ws_13 <= io_in_r_bypass_25_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_0_stall_13 <= io_in_r_bypass_25_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_1_data_13 <= io_in_r_bypass_25_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_1_load_store_13 <= io_in_r_bypass_25_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_1_df_is_ws_13 <= io_in_r_bypass_25_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_1_stall_13 <= io_in_r_bypass_25_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_2_data_13 <= io_in_r_bypass_25_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_2_load_store_13 <= io_in_r_bypass_25_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_2_df_is_ws_13 <= io_in_r_bypass_25_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_2_stall_13 <= io_in_r_bypass_25_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_3_data_13 <= io_in_r_bypass_25_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_3_load_store_13 <= io_in_r_bypass_25_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_3_df_is_ws_13 <= io_in_r_bypass_25_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_3_stall_13 <= io_in_r_bypass_25_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_0_data_13 <= io_in_r_bypass_26_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_0_load_store_13 <= io_in_r_bypass_26_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_0_df_is_ws_13 <= io_in_r_bypass_26_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_0_stall_13 <= io_in_r_bypass_26_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_1_data_13 <= io_in_r_bypass_26_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_1_load_store_13 <= io_in_r_bypass_26_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_1_df_is_ws_13 <= io_in_r_bypass_26_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_1_stall_13 <= io_in_r_bypass_26_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_2_data_13 <= io_in_r_bypass_26_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_2_load_store_13 <= io_in_r_bypass_26_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_2_df_is_ws_13 <= io_in_r_bypass_26_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_2_stall_13 <= io_in_r_bypass_26_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_3_data_13 <= io_in_r_bypass_26_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_3_load_store_13 <= io_in_r_bypass_26_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_3_df_is_ws_13 <= io_in_r_bypass_26_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_3_stall_13 <= io_in_r_bypass_26_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_0_data_13 <= io_in_r_bypass_27_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_0_load_store_13 <= io_in_r_bypass_27_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_0_df_is_ws_13 <= io_in_r_bypass_27_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_0_stall_13 <= io_in_r_bypass_27_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_1_data_13 <= io_in_r_bypass_27_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_1_load_store_13 <= io_in_r_bypass_27_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_1_df_is_ws_13 <= io_in_r_bypass_27_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_1_stall_13 <= io_in_r_bypass_27_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_2_data_13 <= io_in_r_bypass_27_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_2_load_store_13 <= io_in_r_bypass_27_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_2_df_is_ws_13 <= io_in_r_bypass_27_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_2_stall_13 <= io_in_r_bypass_27_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_3_data_13 <= io_in_r_bypass_27_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_3_load_store_13 <= io_in_r_bypass_27_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_3_df_is_ws_13 <= io_in_r_bypass_27_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_3_stall_13 <= io_in_r_bypass_27_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_0_data_13 <= io_in_r_bypass_28_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_0_load_store_13 <= io_in_r_bypass_28_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_0_df_is_ws_13 <= io_in_r_bypass_28_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_0_stall_13 <= io_in_r_bypass_28_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_1_data_13 <= io_in_r_bypass_28_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_1_load_store_13 <= io_in_r_bypass_28_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_1_df_is_ws_13 <= io_in_r_bypass_28_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_1_stall_13 <= io_in_r_bypass_28_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_2_data_13 <= io_in_r_bypass_28_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_2_load_store_13 <= io_in_r_bypass_28_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_2_df_is_ws_13 <= io_in_r_bypass_28_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_2_stall_13 <= io_in_r_bypass_28_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_3_data_13 <= io_in_r_bypass_28_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_3_load_store_13 <= io_in_r_bypass_28_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_3_df_is_ws_13 <= io_in_r_bypass_28_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_3_stall_13 <= io_in_r_bypass_28_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_0_data_13 <= io_in_r_bypass_29_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_0_load_store_13 <= io_in_r_bypass_29_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_0_df_is_ws_13 <= io_in_r_bypass_29_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_0_stall_13 <= io_in_r_bypass_29_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_1_data_13 <= io_in_r_bypass_29_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_1_load_store_13 <= io_in_r_bypass_29_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_1_df_is_ws_13 <= io_in_r_bypass_29_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_1_stall_13 <= io_in_r_bypass_29_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_2_data_13 <= io_in_r_bypass_29_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_2_load_store_13 <= io_in_r_bypass_29_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_2_df_is_ws_13 <= io_in_r_bypass_29_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_2_stall_13 <= io_in_r_bypass_29_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_3_data_13 <= io_in_r_bypass_29_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_3_load_store_13 <= io_in_r_bypass_29_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_3_df_is_ws_13 <= io_in_r_bypass_29_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_3_stall_13 <= io_in_r_bypass_29_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_0_data_13 <= io_in_r_bypass_30_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_0_load_store_13 <= io_in_r_bypass_30_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_0_df_is_ws_13 <= io_in_r_bypass_30_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_0_stall_13 <= io_in_r_bypass_30_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_1_data_13 <= io_in_r_bypass_30_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_1_load_store_13 <= io_in_r_bypass_30_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_1_df_is_ws_13 <= io_in_r_bypass_30_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_1_stall_13 <= io_in_r_bypass_30_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_2_data_13 <= io_in_r_bypass_30_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_2_load_store_13 <= io_in_r_bypass_30_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_2_df_is_ws_13 <= io_in_r_bypass_30_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_2_stall_13 <= io_in_r_bypass_30_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_3_data_13 <= io_in_r_bypass_30_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_3_load_store_13 <= io_in_r_bypass_30_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_3_df_is_ws_13 <= io_in_r_bypass_30_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_3_stall_13 <= io_in_r_bypass_30_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_0_data_13 <= io_in_r_bypass_31_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_0_load_store_13 <= io_in_r_bypass_31_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_0_df_is_ws_13 <= io_in_r_bypass_31_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_0_stall_13 <= io_in_r_bypass_31_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_1_data_13 <= io_in_r_bypass_31_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_1_load_store_13 <= io_in_r_bypass_31_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_1_df_is_ws_13 <= io_in_r_bypass_31_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_1_stall_13 <= io_in_r_bypass_31_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_2_data_13 <= io_in_r_bypass_31_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_2_load_store_13 <= io_in_r_bypass_31_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_2_df_is_ws_13 <= io_in_r_bypass_31_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_2_stall_13 <= io_in_r_bypass_31_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_3_data_13 <= io_in_r_bypass_31_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_3_load_store_13 <= io_in_r_bypass_31_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_3_df_is_ws_13 <= io_in_r_bypass_31_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_3_stall_13 <= io_in_r_bypass_31_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_0_data_14 <= io_in_r_bypass_0_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_0_load_store_14 <= io_in_r_bypass_0_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_0_df_is_ws_14 <= io_in_r_bypass_0_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_0_stall_14 <= io_in_r_bypass_0_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_1_data_14 <= io_in_r_bypass_0_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_1_load_store_14 <= io_in_r_bypass_0_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_1_df_is_ws_14 <= io_in_r_bypass_0_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_1_stall_14 <= io_in_r_bypass_0_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_2_data_14 <= io_in_r_bypass_0_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_2_load_store_14 <= io_in_r_bypass_0_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_2_df_is_ws_14 <= io_in_r_bypass_0_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_2_stall_14 <= io_in_r_bypass_0_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_3_data_14 <= io_in_r_bypass_0_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_3_load_store_14 <= io_in_r_bypass_0_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_3_df_is_ws_14 <= io_in_r_bypass_0_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_3_stall_14 <= io_in_r_bypass_0_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_0_data_14 <= io_in_r_bypass_1_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_0_load_store_14 <= io_in_r_bypass_1_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_0_df_is_ws_14 <= io_in_r_bypass_1_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_0_stall_14 <= io_in_r_bypass_1_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_1_data_14 <= io_in_r_bypass_1_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_1_load_store_14 <= io_in_r_bypass_1_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_1_df_is_ws_14 <= io_in_r_bypass_1_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_1_stall_14 <= io_in_r_bypass_1_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_2_data_14 <= io_in_r_bypass_1_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_2_load_store_14 <= io_in_r_bypass_1_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_2_df_is_ws_14 <= io_in_r_bypass_1_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_2_stall_14 <= io_in_r_bypass_1_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_3_data_14 <= io_in_r_bypass_1_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_3_load_store_14 <= io_in_r_bypass_1_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_3_df_is_ws_14 <= io_in_r_bypass_1_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_3_stall_14 <= io_in_r_bypass_1_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_0_data_14 <= io_in_r_bypass_2_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_0_load_store_14 <= io_in_r_bypass_2_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_0_df_is_ws_14 <= io_in_r_bypass_2_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_0_stall_14 <= io_in_r_bypass_2_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_1_data_14 <= io_in_r_bypass_2_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_1_load_store_14 <= io_in_r_bypass_2_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_1_df_is_ws_14 <= io_in_r_bypass_2_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_1_stall_14 <= io_in_r_bypass_2_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_2_data_14 <= io_in_r_bypass_2_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_2_load_store_14 <= io_in_r_bypass_2_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_2_df_is_ws_14 <= io_in_r_bypass_2_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_2_stall_14 <= io_in_r_bypass_2_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_3_data_14 <= io_in_r_bypass_2_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_3_load_store_14 <= io_in_r_bypass_2_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_3_df_is_ws_14 <= io_in_r_bypass_2_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_3_stall_14 <= io_in_r_bypass_2_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_0_data_14 <= io_in_r_bypass_3_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_0_load_store_14 <= io_in_r_bypass_3_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_0_df_is_ws_14 <= io_in_r_bypass_3_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_0_stall_14 <= io_in_r_bypass_3_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_1_data_14 <= io_in_r_bypass_3_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_1_load_store_14 <= io_in_r_bypass_3_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_1_df_is_ws_14 <= io_in_r_bypass_3_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_1_stall_14 <= io_in_r_bypass_3_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_2_data_14 <= io_in_r_bypass_3_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_2_load_store_14 <= io_in_r_bypass_3_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_2_df_is_ws_14 <= io_in_r_bypass_3_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_2_stall_14 <= io_in_r_bypass_3_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_3_data_14 <= io_in_r_bypass_3_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_3_load_store_14 <= io_in_r_bypass_3_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_3_df_is_ws_14 <= io_in_r_bypass_3_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_3_stall_14 <= io_in_r_bypass_3_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_0_data_14 <= io_in_r_bypass_4_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_0_load_store_14 <= io_in_r_bypass_4_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_0_df_is_ws_14 <= io_in_r_bypass_4_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_0_stall_14 <= io_in_r_bypass_4_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_1_data_14 <= io_in_r_bypass_4_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_1_load_store_14 <= io_in_r_bypass_4_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_1_df_is_ws_14 <= io_in_r_bypass_4_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_1_stall_14 <= io_in_r_bypass_4_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_2_data_14 <= io_in_r_bypass_4_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_2_load_store_14 <= io_in_r_bypass_4_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_2_df_is_ws_14 <= io_in_r_bypass_4_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_2_stall_14 <= io_in_r_bypass_4_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_3_data_14 <= io_in_r_bypass_4_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_3_load_store_14 <= io_in_r_bypass_4_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_3_df_is_ws_14 <= io_in_r_bypass_4_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_3_stall_14 <= io_in_r_bypass_4_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_0_data_14 <= io_in_r_bypass_5_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_0_load_store_14 <= io_in_r_bypass_5_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_0_df_is_ws_14 <= io_in_r_bypass_5_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_0_stall_14 <= io_in_r_bypass_5_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_1_data_14 <= io_in_r_bypass_5_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_1_load_store_14 <= io_in_r_bypass_5_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_1_df_is_ws_14 <= io_in_r_bypass_5_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_1_stall_14 <= io_in_r_bypass_5_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_2_data_14 <= io_in_r_bypass_5_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_2_load_store_14 <= io_in_r_bypass_5_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_2_df_is_ws_14 <= io_in_r_bypass_5_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_2_stall_14 <= io_in_r_bypass_5_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_3_data_14 <= io_in_r_bypass_5_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_3_load_store_14 <= io_in_r_bypass_5_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_3_df_is_ws_14 <= io_in_r_bypass_5_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_3_stall_14 <= io_in_r_bypass_5_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_0_data_14 <= io_in_r_bypass_6_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_0_load_store_14 <= io_in_r_bypass_6_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_0_df_is_ws_14 <= io_in_r_bypass_6_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_0_stall_14 <= io_in_r_bypass_6_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_1_data_14 <= io_in_r_bypass_6_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_1_load_store_14 <= io_in_r_bypass_6_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_1_df_is_ws_14 <= io_in_r_bypass_6_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_1_stall_14 <= io_in_r_bypass_6_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_2_data_14 <= io_in_r_bypass_6_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_2_load_store_14 <= io_in_r_bypass_6_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_2_df_is_ws_14 <= io_in_r_bypass_6_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_2_stall_14 <= io_in_r_bypass_6_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_3_data_14 <= io_in_r_bypass_6_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_3_load_store_14 <= io_in_r_bypass_6_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_3_df_is_ws_14 <= io_in_r_bypass_6_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_3_stall_14 <= io_in_r_bypass_6_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_0_data_14 <= io_in_r_bypass_7_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_0_load_store_14 <= io_in_r_bypass_7_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_0_df_is_ws_14 <= io_in_r_bypass_7_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_0_stall_14 <= io_in_r_bypass_7_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_1_data_14 <= io_in_r_bypass_7_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_1_load_store_14 <= io_in_r_bypass_7_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_1_df_is_ws_14 <= io_in_r_bypass_7_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_1_stall_14 <= io_in_r_bypass_7_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_2_data_14 <= io_in_r_bypass_7_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_2_load_store_14 <= io_in_r_bypass_7_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_2_df_is_ws_14 <= io_in_r_bypass_7_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_2_stall_14 <= io_in_r_bypass_7_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_3_data_14 <= io_in_r_bypass_7_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_3_load_store_14 <= io_in_r_bypass_7_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_3_df_is_ws_14 <= io_in_r_bypass_7_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_3_stall_14 <= io_in_r_bypass_7_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_0_data_14 <= io_in_r_bypass_8_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_0_load_store_14 <= io_in_r_bypass_8_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_0_df_is_ws_14 <= io_in_r_bypass_8_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_0_stall_14 <= io_in_r_bypass_8_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_1_data_14 <= io_in_r_bypass_8_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_1_load_store_14 <= io_in_r_bypass_8_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_1_df_is_ws_14 <= io_in_r_bypass_8_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_1_stall_14 <= io_in_r_bypass_8_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_2_data_14 <= io_in_r_bypass_8_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_2_load_store_14 <= io_in_r_bypass_8_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_2_df_is_ws_14 <= io_in_r_bypass_8_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_2_stall_14 <= io_in_r_bypass_8_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_3_data_14 <= io_in_r_bypass_8_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_3_load_store_14 <= io_in_r_bypass_8_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_3_df_is_ws_14 <= io_in_r_bypass_8_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_3_stall_14 <= io_in_r_bypass_8_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_0_data_14 <= io_in_r_bypass_9_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_0_load_store_14 <= io_in_r_bypass_9_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_0_df_is_ws_14 <= io_in_r_bypass_9_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_0_stall_14 <= io_in_r_bypass_9_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_1_data_14 <= io_in_r_bypass_9_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_1_load_store_14 <= io_in_r_bypass_9_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_1_df_is_ws_14 <= io_in_r_bypass_9_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_1_stall_14 <= io_in_r_bypass_9_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_2_data_14 <= io_in_r_bypass_9_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_2_load_store_14 <= io_in_r_bypass_9_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_2_df_is_ws_14 <= io_in_r_bypass_9_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_2_stall_14 <= io_in_r_bypass_9_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_3_data_14 <= io_in_r_bypass_9_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_3_load_store_14 <= io_in_r_bypass_9_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_3_df_is_ws_14 <= io_in_r_bypass_9_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_3_stall_14 <= io_in_r_bypass_9_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_0_data_14 <= io_in_r_bypass_10_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_0_load_store_14 <= io_in_r_bypass_10_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_0_df_is_ws_14 <= io_in_r_bypass_10_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_0_stall_14 <= io_in_r_bypass_10_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_1_data_14 <= io_in_r_bypass_10_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_1_load_store_14 <= io_in_r_bypass_10_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_1_df_is_ws_14 <= io_in_r_bypass_10_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_1_stall_14 <= io_in_r_bypass_10_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_2_data_14 <= io_in_r_bypass_10_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_2_load_store_14 <= io_in_r_bypass_10_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_2_df_is_ws_14 <= io_in_r_bypass_10_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_2_stall_14 <= io_in_r_bypass_10_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_3_data_14 <= io_in_r_bypass_10_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_3_load_store_14 <= io_in_r_bypass_10_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_3_df_is_ws_14 <= io_in_r_bypass_10_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_3_stall_14 <= io_in_r_bypass_10_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_0_data_14 <= io_in_r_bypass_11_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_0_load_store_14 <= io_in_r_bypass_11_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_0_df_is_ws_14 <= io_in_r_bypass_11_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_0_stall_14 <= io_in_r_bypass_11_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_1_data_14 <= io_in_r_bypass_11_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_1_load_store_14 <= io_in_r_bypass_11_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_1_df_is_ws_14 <= io_in_r_bypass_11_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_1_stall_14 <= io_in_r_bypass_11_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_2_data_14 <= io_in_r_bypass_11_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_2_load_store_14 <= io_in_r_bypass_11_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_2_df_is_ws_14 <= io_in_r_bypass_11_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_2_stall_14 <= io_in_r_bypass_11_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_3_data_14 <= io_in_r_bypass_11_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_3_load_store_14 <= io_in_r_bypass_11_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_3_df_is_ws_14 <= io_in_r_bypass_11_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_3_stall_14 <= io_in_r_bypass_11_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_0_data_14 <= io_in_r_bypass_12_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_0_load_store_14 <= io_in_r_bypass_12_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_0_df_is_ws_14 <= io_in_r_bypass_12_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_0_stall_14 <= io_in_r_bypass_12_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_1_data_14 <= io_in_r_bypass_12_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_1_load_store_14 <= io_in_r_bypass_12_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_1_df_is_ws_14 <= io_in_r_bypass_12_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_1_stall_14 <= io_in_r_bypass_12_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_2_data_14 <= io_in_r_bypass_12_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_2_load_store_14 <= io_in_r_bypass_12_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_2_df_is_ws_14 <= io_in_r_bypass_12_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_2_stall_14 <= io_in_r_bypass_12_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_3_data_14 <= io_in_r_bypass_12_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_3_load_store_14 <= io_in_r_bypass_12_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_3_df_is_ws_14 <= io_in_r_bypass_12_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_3_stall_14 <= io_in_r_bypass_12_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_0_data_14 <= io_in_r_bypass_13_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_0_load_store_14 <= io_in_r_bypass_13_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_0_df_is_ws_14 <= io_in_r_bypass_13_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_0_stall_14 <= io_in_r_bypass_13_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_1_data_14 <= io_in_r_bypass_13_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_1_load_store_14 <= io_in_r_bypass_13_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_1_df_is_ws_14 <= io_in_r_bypass_13_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_1_stall_14 <= io_in_r_bypass_13_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_2_data_14 <= io_in_r_bypass_13_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_2_load_store_14 <= io_in_r_bypass_13_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_2_df_is_ws_14 <= io_in_r_bypass_13_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_2_stall_14 <= io_in_r_bypass_13_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_3_data_14 <= io_in_r_bypass_13_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_3_load_store_14 <= io_in_r_bypass_13_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_3_df_is_ws_14 <= io_in_r_bypass_13_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_3_stall_14 <= io_in_r_bypass_13_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_0_data_14 <= io_in_r_bypass_14_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_0_load_store_14 <= io_in_r_bypass_14_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_0_df_is_ws_14 <= io_in_r_bypass_14_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_0_stall_14 <= io_in_r_bypass_14_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_1_data_14 <= io_in_r_bypass_14_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_1_load_store_14 <= io_in_r_bypass_14_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_1_df_is_ws_14 <= io_in_r_bypass_14_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_1_stall_14 <= io_in_r_bypass_14_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_2_data_14 <= io_in_r_bypass_14_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_2_load_store_14 <= io_in_r_bypass_14_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_2_df_is_ws_14 <= io_in_r_bypass_14_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_2_stall_14 <= io_in_r_bypass_14_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_3_data_14 <= io_in_r_bypass_14_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_3_load_store_14 <= io_in_r_bypass_14_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_3_df_is_ws_14 <= io_in_r_bypass_14_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_3_stall_14 <= io_in_r_bypass_14_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_0_data_14 <= io_in_r_bypass_15_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_0_load_store_14 <= io_in_r_bypass_15_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_0_df_is_ws_14 <= io_in_r_bypass_15_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_0_stall_14 <= io_in_r_bypass_15_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_1_data_14 <= io_in_r_bypass_15_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_1_load_store_14 <= io_in_r_bypass_15_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_1_df_is_ws_14 <= io_in_r_bypass_15_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_1_stall_14 <= io_in_r_bypass_15_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_2_data_14 <= io_in_r_bypass_15_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_2_load_store_14 <= io_in_r_bypass_15_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_2_df_is_ws_14 <= io_in_r_bypass_15_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_2_stall_14 <= io_in_r_bypass_15_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_3_data_14 <= io_in_r_bypass_15_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_3_load_store_14 <= io_in_r_bypass_15_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_3_df_is_ws_14 <= io_in_r_bypass_15_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_3_stall_14 <= io_in_r_bypass_15_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_0_data_14 <= io_in_r_bypass_16_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_0_load_store_14 <= io_in_r_bypass_16_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_0_df_is_ws_14 <= io_in_r_bypass_16_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_0_stall_14 <= io_in_r_bypass_16_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_1_data_14 <= io_in_r_bypass_16_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_1_load_store_14 <= io_in_r_bypass_16_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_1_df_is_ws_14 <= io_in_r_bypass_16_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_1_stall_14 <= io_in_r_bypass_16_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_2_data_14 <= io_in_r_bypass_16_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_2_load_store_14 <= io_in_r_bypass_16_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_2_df_is_ws_14 <= io_in_r_bypass_16_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_2_stall_14 <= io_in_r_bypass_16_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_3_data_14 <= io_in_r_bypass_16_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_3_load_store_14 <= io_in_r_bypass_16_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_3_df_is_ws_14 <= io_in_r_bypass_16_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_3_stall_14 <= io_in_r_bypass_16_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_0_data_14 <= io_in_r_bypass_17_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_0_load_store_14 <= io_in_r_bypass_17_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_0_df_is_ws_14 <= io_in_r_bypass_17_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_0_stall_14 <= io_in_r_bypass_17_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_1_data_14 <= io_in_r_bypass_17_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_1_load_store_14 <= io_in_r_bypass_17_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_1_df_is_ws_14 <= io_in_r_bypass_17_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_1_stall_14 <= io_in_r_bypass_17_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_2_data_14 <= io_in_r_bypass_17_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_2_load_store_14 <= io_in_r_bypass_17_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_2_df_is_ws_14 <= io_in_r_bypass_17_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_2_stall_14 <= io_in_r_bypass_17_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_3_data_14 <= io_in_r_bypass_17_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_3_load_store_14 <= io_in_r_bypass_17_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_3_df_is_ws_14 <= io_in_r_bypass_17_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_3_stall_14 <= io_in_r_bypass_17_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_0_data_14 <= io_in_r_bypass_18_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_0_load_store_14 <= io_in_r_bypass_18_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_0_df_is_ws_14 <= io_in_r_bypass_18_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_0_stall_14 <= io_in_r_bypass_18_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_1_data_14 <= io_in_r_bypass_18_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_1_load_store_14 <= io_in_r_bypass_18_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_1_df_is_ws_14 <= io_in_r_bypass_18_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_1_stall_14 <= io_in_r_bypass_18_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_2_data_14 <= io_in_r_bypass_18_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_2_load_store_14 <= io_in_r_bypass_18_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_2_df_is_ws_14 <= io_in_r_bypass_18_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_2_stall_14 <= io_in_r_bypass_18_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_3_data_14 <= io_in_r_bypass_18_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_3_load_store_14 <= io_in_r_bypass_18_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_3_df_is_ws_14 <= io_in_r_bypass_18_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_3_stall_14 <= io_in_r_bypass_18_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_0_data_14 <= io_in_r_bypass_19_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_0_load_store_14 <= io_in_r_bypass_19_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_0_df_is_ws_14 <= io_in_r_bypass_19_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_0_stall_14 <= io_in_r_bypass_19_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_1_data_14 <= io_in_r_bypass_19_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_1_load_store_14 <= io_in_r_bypass_19_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_1_df_is_ws_14 <= io_in_r_bypass_19_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_1_stall_14 <= io_in_r_bypass_19_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_2_data_14 <= io_in_r_bypass_19_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_2_load_store_14 <= io_in_r_bypass_19_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_2_df_is_ws_14 <= io_in_r_bypass_19_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_2_stall_14 <= io_in_r_bypass_19_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_3_data_14 <= io_in_r_bypass_19_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_3_load_store_14 <= io_in_r_bypass_19_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_3_df_is_ws_14 <= io_in_r_bypass_19_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_3_stall_14 <= io_in_r_bypass_19_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_0_data_14 <= io_in_r_bypass_20_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_0_load_store_14 <= io_in_r_bypass_20_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_0_df_is_ws_14 <= io_in_r_bypass_20_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_0_stall_14 <= io_in_r_bypass_20_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_1_data_14 <= io_in_r_bypass_20_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_1_load_store_14 <= io_in_r_bypass_20_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_1_df_is_ws_14 <= io_in_r_bypass_20_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_1_stall_14 <= io_in_r_bypass_20_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_2_data_14 <= io_in_r_bypass_20_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_2_load_store_14 <= io_in_r_bypass_20_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_2_df_is_ws_14 <= io_in_r_bypass_20_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_2_stall_14 <= io_in_r_bypass_20_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_3_data_14 <= io_in_r_bypass_20_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_3_load_store_14 <= io_in_r_bypass_20_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_3_df_is_ws_14 <= io_in_r_bypass_20_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_3_stall_14 <= io_in_r_bypass_20_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_0_data_14 <= io_in_r_bypass_21_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_0_load_store_14 <= io_in_r_bypass_21_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_0_df_is_ws_14 <= io_in_r_bypass_21_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_0_stall_14 <= io_in_r_bypass_21_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_1_data_14 <= io_in_r_bypass_21_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_1_load_store_14 <= io_in_r_bypass_21_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_1_df_is_ws_14 <= io_in_r_bypass_21_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_1_stall_14 <= io_in_r_bypass_21_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_2_data_14 <= io_in_r_bypass_21_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_2_load_store_14 <= io_in_r_bypass_21_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_2_df_is_ws_14 <= io_in_r_bypass_21_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_2_stall_14 <= io_in_r_bypass_21_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_3_data_14 <= io_in_r_bypass_21_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_3_load_store_14 <= io_in_r_bypass_21_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_3_df_is_ws_14 <= io_in_r_bypass_21_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_3_stall_14 <= io_in_r_bypass_21_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_0_data_14 <= io_in_r_bypass_22_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_0_load_store_14 <= io_in_r_bypass_22_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_0_df_is_ws_14 <= io_in_r_bypass_22_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_0_stall_14 <= io_in_r_bypass_22_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_1_data_14 <= io_in_r_bypass_22_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_1_load_store_14 <= io_in_r_bypass_22_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_1_df_is_ws_14 <= io_in_r_bypass_22_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_1_stall_14 <= io_in_r_bypass_22_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_2_data_14 <= io_in_r_bypass_22_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_2_load_store_14 <= io_in_r_bypass_22_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_2_df_is_ws_14 <= io_in_r_bypass_22_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_2_stall_14 <= io_in_r_bypass_22_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_3_data_14 <= io_in_r_bypass_22_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_3_load_store_14 <= io_in_r_bypass_22_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_3_df_is_ws_14 <= io_in_r_bypass_22_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_3_stall_14 <= io_in_r_bypass_22_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_0_data_14 <= io_in_r_bypass_23_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_0_load_store_14 <= io_in_r_bypass_23_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_0_df_is_ws_14 <= io_in_r_bypass_23_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_0_stall_14 <= io_in_r_bypass_23_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_1_data_14 <= io_in_r_bypass_23_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_1_load_store_14 <= io_in_r_bypass_23_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_1_df_is_ws_14 <= io_in_r_bypass_23_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_1_stall_14 <= io_in_r_bypass_23_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_2_data_14 <= io_in_r_bypass_23_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_2_load_store_14 <= io_in_r_bypass_23_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_2_df_is_ws_14 <= io_in_r_bypass_23_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_2_stall_14 <= io_in_r_bypass_23_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_3_data_14 <= io_in_r_bypass_23_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_3_load_store_14 <= io_in_r_bypass_23_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_3_df_is_ws_14 <= io_in_r_bypass_23_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_3_stall_14 <= io_in_r_bypass_23_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_0_data_14 <= io_in_r_bypass_24_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_0_load_store_14 <= io_in_r_bypass_24_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_0_df_is_ws_14 <= io_in_r_bypass_24_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_0_stall_14 <= io_in_r_bypass_24_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_1_data_14 <= io_in_r_bypass_24_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_1_load_store_14 <= io_in_r_bypass_24_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_1_df_is_ws_14 <= io_in_r_bypass_24_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_1_stall_14 <= io_in_r_bypass_24_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_2_data_14 <= io_in_r_bypass_24_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_2_load_store_14 <= io_in_r_bypass_24_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_2_df_is_ws_14 <= io_in_r_bypass_24_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_2_stall_14 <= io_in_r_bypass_24_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_3_data_14 <= io_in_r_bypass_24_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_3_load_store_14 <= io_in_r_bypass_24_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_3_df_is_ws_14 <= io_in_r_bypass_24_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_3_stall_14 <= io_in_r_bypass_24_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_0_data_14 <= io_in_r_bypass_25_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_0_load_store_14 <= io_in_r_bypass_25_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_0_df_is_ws_14 <= io_in_r_bypass_25_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_0_stall_14 <= io_in_r_bypass_25_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_1_data_14 <= io_in_r_bypass_25_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_1_load_store_14 <= io_in_r_bypass_25_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_1_df_is_ws_14 <= io_in_r_bypass_25_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_1_stall_14 <= io_in_r_bypass_25_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_2_data_14 <= io_in_r_bypass_25_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_2_load_store_14 <= io_in_r_bypass_25_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_2_df_is_ws_14 <= io_in_r_bypass_25_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_2_stall_14 <= io_in_r_bypass_25_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_3_data_14 <= io_in_r_bypass_25_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_3_load_store_14 <= io_in_r_bypass_25_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_3_df_is_ws_14 <= io_in_r_bypass_25_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_3_stall_14 <= io_in_r_bypass_25_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_0_data_14 <= io_in_r_bypass_26_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_0_load_store_14 <= io_in_r_bypass_26_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_0_df_is_ws_14 <= io_in_r_bypass_26_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_0_stall_14 <= io_in_r_bypass_26_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_1_data_14 <= io_in_r_bypass_26_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_1_load_store_14 <= io_in_r_bypass_26_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_1_df_is_ws_14 <= io_in_r_bypass_26_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_1_stall_14 <= io_in_r_bypass_26_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_2_data_14 <= io_in_r_bypass_26_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_2_load_store_14 <= io_in_r_bypass_26_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_2_df_is_ws_14 <= io_in_r_bypass_26_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_2_stall_14 <= io_in_r_bypass_26_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_3_data_14 <= io_in_r_bypass_26_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_3_load_store_14 <= io_in_r_bypass_26_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_3_df_is_ws_14 <= io_in_r_bypass_26_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_3_stall_14 <= io_in_r_bypass_26_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_0_data_14 <= io_in_r_bypass_27_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_0_load_store_14 <= io_in_r_bypass_27_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_0_df_is_ws_14 <= io_in_r_bypass_27_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_0_stall_14 <= io_in_r_bypass_27_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_1_data_14 <= io_in_r_bypass_27_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_1_load_store_14 <= io_in_r_bypass_27_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_1_df_is_ws_14 <= io_in_r_bypass_27_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_1_stall_14 <= io_in_r_bypass_27_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_2_data_14 <= io_in_r_bypass_27_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_2_load_store_14 <= io_in_r_bypass_27_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_2_df_is_ws_14 <= io_in_r_bypass_27_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_2_stall_14 <= io_in_r_bypass_27_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_3_data_14 <= io_in_r_bypass_27_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_3_load_store_14 <= io_in_r_bypass_27_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_3_df_is_ws_14 <= io_in_r_bypass_27_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_3_stall_14 <= io_in_r_bypass_27_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_0_data_14 <= io_in_r_bypass_28_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_0_load_store_14 <= io_in_r_bypass_28_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_0_df_is_ws_14 <= io_in_r_bypass_28_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_0_stall_14 <= io_in_r_bypass_28_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_1_data_14 <= io_in_r_bypass_28_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_1_load_store_14 <= io_in_r_bypass_28_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_1_df_is_ws_14 <= io_in_r_bypass_28_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_1_stall_14 <= io_in_r_bypass_28_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_2_data_14 <= io_in_r_bypass_28_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_2_load_store_14 <= io_in_r_bypass_28_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_2_df_is_ws_14 <= io_in_r_bypass_28_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_2_stall_14 <= io_in_r_bypass_28_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_3_data_14 <= io_in_r_bypass_28_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_3_load_store_14 <= io_in_r_bypass_28_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_3_df_is_ws_14 <= io_in_r_bypass_28_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_3_stall_14 <= io_in_r_bypass_28_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_0_data_14 <= io_in_r_bypass_29_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_0_load_store_14 <= io_in_r_bypass_29_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_0_df_is_ws_14 <= io_in_r_bypass_29_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_0_stall_14 <= io_in_r_bypass_29_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_1_data_14 <= io_in_r_bypass_29_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_1_load_store_14 <= io_in_r_bypass_29_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_1_df_is_ws_14 <= io_in_r_bypass_29_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_1_stall_14 <= io_in_r_bypass_29_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_2_data_14 <= io_in_r_bypass_29_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_2_load_store_14 <= io_in_r_bypass_29_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_2_df_is_ws_14 <= io_in_r_bypass_29_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_2_stall_14 <= io_in_r_bypass_29_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_3_data_14 <= io_in_r_bypass_29_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_3_load_store_14 <= io_in_r_bypass_29_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_3_df_is_ws_14 <= io_in_r_bypass_29_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_3_stall_14 <= io_in_r_bypass_29_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_0_data_14 <= io_in_r_bypass_30_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_0_load_store_14 <= io_in_r_bypass_30_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_0_df_is_ws_14 <= io_in_r_bypass_30_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_0_stall_14 <= io_in_r_bypass_30_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_1_data_14 <= io_in_r_bypass_30_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_1_load_store_14 <= io_in_r_bypass_30_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_1_df_is_ws_14 <= io_in_r_bypass_30_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_1_stall_14 <= io_in_r_bypass_30_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_2_data_14 <= io_in_r_bypass_30_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_2_load_store_14 <= io_in_r_bypass_30_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_2_df_is_ws_14 <= io_in_r_bypass_30_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_2_stall_14 <= io_in_r_bypass_30_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_3_data_14 <= io_in_r_bypass_30_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_3_load_store_14 <= io_in_r_bypass_30_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_3_df_is_ws_14 <= io_in_r_bypass_30_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_3_stall_14 <= io_in_r_bypass_30_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_0_data_14 <= io_in_r_bypass_31_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_0_load_store_14 <= io_in_r_bypass_31_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_0_df_is_ws_14 <= io_in_r_bypass_31_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_0_stall_14 <= io_in_r_bypass_31_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_1_data_14 <= io_in_r_bypass_31_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_1_load_store_14 <= io_in_r_bypass_31_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_1_df_is_ws_14 <= io_in_r_bypass_31_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_1_stall_14 <= io_in_r_bypass_31_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_2_data_14 <= io_in_r_bypass_31_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_2_load_store_14 <= io_in_r_bypass_31_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_2_df_is_ws_14 <= io_in_r_bypass_31_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_2_stall_14 <= io_in_r_bypass_31_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_3_data_14 <= io_in_r_bypass_31_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_3_load_store_14 <= io_in_r_bypass_31_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_3_df_is_ws_14 <= io_in_r_bypass_31_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_3_stall_14 <= io_in_r_bypass_31_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_0_data_15 <= io_in_r_bypass_0_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_0_load_store_15 <= io_in_r_bypass_0_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_0_df_is_ws_15 <= io_in_r_bypass_0_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_0_stall_15 <= io_in_r_bypass_0_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_1_data_15 <= io_in_r_bypass_0_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_1_load_store_15 <= io_in_r_bypass_0_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_1_df_is_ws_15 <= io_in_r_bypass_0_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_1_stall_15 <= io_in_r_bypass_0_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_2_data_15 <= io_in_r_bypass_0_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_2_load_store_15 <= io_in_r_bypass_0_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_2_df_is_ws_15 <= io_in_r_bypass_0_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_2_stall_15 <= io_in_r_bypass_0_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_3_data_15 <= io_in_r_bypass_0_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_3_load_store_15 <= io_in_r_bypass_0_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_3_df_is_ws_15 <= io_in_r_bypass_0_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_3_stall_15 <= io_in_r_bypass_0_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_0_data_15 <= io_in_r_bypass_1_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_0_load_store_15 <= io_in_r_bypass_1_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_0_df_is_ws_15 <= io_in_r_bypass_1_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_0_stall_15 <= io_in_r_bypass_1_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_1_data_15 <= io_in_r_bypass_1_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_1_load_store_15 <= io_in_r_bypass_1_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_1_df_is_ws_15 <= io_in_r_bypass_1_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_1_stall_15 <= io_in_r_bypass_1_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_2_data_15 <= io_in_r_bypass_1_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_2_load_store_15 <= io_in_r_bypass_1_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_2_df_is_ws_15 <= io_in_r_bypass_1_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_2_stall_15 <= io_in_r_bypass_1_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_3_data_15 <= io_in_r_bypass_1_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_3_load_store_15 <= io_in_r_bypass_1_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_3_df_is_ws_15 <= io_in_r_bypass_1_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_3_stall_15 <= io_in_r_bypass_1_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_0_data_15 <= io_in_r_bypass_2_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_0_load_store_15 <= io_in_r_bypass_2_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_0_df_is_ws_15 <= io_in_r_bypass_2_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_0_stall_15 <= io_in_r_bypass_2_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_1_data_15 <= io_in_r_bypass_2_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_1_load_store_15 <= io_in_r_bypass_2_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_1_df_is_ws_15 <= io_in_r_bypass_2_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_1_stall_15 <= io_in_r_bypass_2_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_2_data_15 <= io_in_r_bypass_2_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_2_load_store_15 <= io_in_r_bypass_2_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_2_df_is_ws_15 <= io_in_r_bypass_2_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_2_stall_15 <= io_in_r_bypass_2_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_3_data_15 <= io_in_r_bypass_2_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_3_load_store_15 <= io_in_r_bypass_2_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_3_df_is_ws_15 <= io_in_r_bypass_2_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_3_stall_15 <= io_in_r_bypass_2_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_0_data_15 <= io_in_r_bypass_3_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_0_load_store_15 <= io_in_r_bypass_3_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_0_df_is_ws_15 <= io_in_r_bypass_3_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_0_stall_15 <= io_in_r_bypass_3_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_1_data_15 <= io_in_r_bypass_3_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_1_load_store_15 <= io_in_r_bypass_3_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_1_df_is_ws_15 <= io_in_r_bypass_3_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_1_stall_15 <= io_in_r_bypass_3_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_2_data_15 <= io_in_r_bypass_3_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_2_load_store_15 <= io_in_r_bypass_3_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_2_df_is_ws_15 <= io_in_r_bypass_3_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_2_stall_15 <= io_in_r_bypass_3_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_3_data_15 <= io_in_r_bypass_3_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_3_load_store_15 <= io_in_r_bypass_3_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_3_df_is_ws_15 <= io_in_r_bypass_3_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_3_stall_15 <= io_in_r_bypass_3_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_0_data_15 <= io_in_r_bypass_4_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_0_load_store_15 <= io_in_r_bypass_4_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_0_df_is_ws_15 <= io_in_r_bypass_4_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_0_stall_15 <= io_in_r_bypass_4_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_1_data_15 <= io_in_r_bypass_4_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_1_load_store_15 <= io_in_r_bypass_4_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_1_df_is_ws_15 <= io_in_r_bypass_4_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_1_stall_15 <= io_in_r_bypass_4_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_2_data_15 <= io_in_r_bypass_4_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_2_load_store_15 <= io_in_r_bypass_4_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_2_df_is_ws_15 <= io_in_r_bypass_4_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_2_stall_15 <= io_in_r_bypass_4_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_3_data_15 <= io_in_r_bypass_4_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_3_load_store_15 <= io_in_r_bypass_4_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_3_df_is_ws_15 <= io_in_r_bypass_4_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_3_stall_15 <= io_in_r_bypass_4_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_0_data_15 <= io_in_r_bypass_5_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_0_load_store_15 <= io_in_r_bypass_5_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_0_df_is_ws_15 <= io_in_r_bypass_5_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_0_stall_15 <= io_in_r_bypass_5_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_1_data_15 <= io_in_r_bypass_5_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_1_load_store_15 <= io_in_r_bypass_5_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_1_df_is_ws_15 <= io_in_r_bypass_5_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_1_stall_15 <= io_in_r_bypass_5_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_2_data_15 <= io_in_r_bypass_5_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_2_load_store_15 <= io_in_r_bypass_5_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_2_df_is_ws_15 <= io_in_r_bypass_5_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_2_stall_15 <= io_in_r_bypass_5_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_3_data_15 <= io_in_r_bypass_5_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_3_load_store_15 <= io_in_r_bypass_5_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_3_df_is_ws_15 <= io_in_r_bypass_5_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_3_stall_15 <= io_in_r_bypass_5_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_0_data_15 <= io_in_r_bypass_6_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_0_load_store_15 <= io_in_r_bypass_6_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_0_df_is_ws_15 <= io_in_r_bypass_6_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_0_stall_15 <= io_in_r_bypass_6_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_1_data_15 <= io_in_r_bypass_6_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_1_load_store_15 <= io_in_r_bypass_6_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_1_df_is_ws_15 <= io_in_r_bypass_6_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_1_stall_15 <= io_in_r_bypass_6_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_2_data_15 <= io_in_r_bypass_6_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_2_load_store_15 <= io_in_r_bypass_6_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_2_df_is_ws_15 <= io_in_r_bypass_6_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_2_stall_15 <= io_in_r_bypass_6_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_3_data_15 <= io_in_r_bypass_6_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_3_load_store_15 <= io_in_r_bypass_6_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_3_df_is_ws_15 <= io_in_r_bypass_6_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_3_stall_15 <= io_in_r_bypass_6_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_0_data_15 <= io_in_r_bypass_7_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_0_load_store_15 <= io_in_r_bypass_7_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_0_df_is_ws_15 <= io_in_r_bypass_7_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_0_stall_15 <= io_in_r_bypass_7_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_1_data_15 <= io_in_r_bypass_7_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_1_load_store_15 <= io_in_r_bypass_7_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_1_df_is_ws_15 <= io_in_r_bypass_7_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_1_stall_15 <= io_in_r_bypass_7_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_2_data_15 <= io_in_r_bypass_7_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_2_load_store_15 <= io_in_r_bypass_7_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_2_df_is_ws_15 <= io_in_r_bypass_7_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_2_stall_15 <= io_in_r_bypass_7_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_3_data_15 <= io_in_r_bypass_7_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_3_load_store_15 <= io_in_r_bypass_7_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_3_df_is_ws_15 <= io_in_r_bypass_7_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_3_stall_15 <= io_in_r_bypass_7_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_0_data_15 <= io_in_r_bypass_8_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_0_load_store_15 <= io_in_r_bypass_8_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_0_df_is_ws_15 <= io_in_r_bypass_8_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_0_stall_15 <= io_in_r_bypass_8_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_1_data_15 <= io_in_r_bypass_8_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_1_load_store_15 <= io_in_r_bypass_8_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_1_df_is_ws_15 <= io_in_r_bypass_8_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_1_stall_15 <= io_in_r_bypass_8_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_2_data_15 <= io_in_r_bypass_8_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_2_load_store_15 <= io_in_r_bypass_8_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_2_df_is_ws_15 <= io_in_r_bypass_8_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_2_stall_15 <= io_in_r_bypass_8_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_3_data_15 <= io_in_r_bypass_8_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_3_load_store_15 <= io_in_r_bypass_8_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_3_df_is_ws_15 <= io_in_r_bypass_8_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_3_stall_15 <= io_in_r_bypass_8_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_0_data_15 <= io_in_r_bypass_9_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_0_load_store_15 <= io_in_r_bypass_9_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_0_df_is_ws_15 <= io_in_r_bypass_9_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_0_stall_15 <= io_in_r_bypass_9_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_1_data_15 <= io_in_r_bypass_9_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_1_load_store_15 <= io_in_r_bypass_9_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_1_df_is_ws_15 <= io_in_r_bypass_9_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_1_stall_15 <= io_in_r_bypass_9_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_2_data_15 <= io_in_r_bypass_9_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_2_load_store_15 <= io_in_r_bypass_9_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_2_df_is_ws_15 <= io_in_r_bypass_9_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_2_stall_15 <= io_in_r_bypass_9_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_3_data_15 <= io_in_r_bypass_9_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_3_load_store_15 <= io_in_r_bypass_9_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_3_df_is_ws_15 <= io_in_r_bypass_9_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_3_stall_15 <= io_in_r_bypass_9_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_0_data_15 <= io_in_r_bypass_10_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_0_load_store_15 <= io_in_r_bypass_10_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_0_df_is_ws_15 <= io_in_r_bypass_10_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_0_stall_15 <= io_in_r_bypass_10_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_1_data_15 <= io_in_r_bypass_10_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_1_load_store_15 <= io_in_r_bypass_10_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_1_df_is_ws_15 <= io_in_r_bypass_10_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_1_stall_15 <= io_in_r_bypass_10_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_2_data_15 <= io_in_r_bypass_10_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_2_load_store_15 <= io_in_r_bypass_10_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_2_df_is_ws_15 <= io_in_r_bypass_10_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_2_stall_15 <= io_in_r_bypass_10_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_3_data_15 <= io_in_r_bypass_10_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_3_load_store_15 <= io_in_r_bypass_10_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_3_df_is_ws_15 <= io_in_r_bypass_10_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_3_stall_15 <= io_in_r_bypass_10_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_0_data_15 <= io_in_r_bypass_11_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_0_load_store_15 <= io_in_r_bypass_11_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_0_df_is_ws_15 <= io_in_r_bypass_11_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_0_stall_15 <= io_in_r_bypass_11_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_1_data_15 <= io_in_r_bypass_11_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_1_load_store_15 <= io_in_r_bypass_11_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_1_df_is_ws_15 <= io_in_r_bypass_11_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_1_stall_15 <= io_in_r_bypass_11_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_2_data_15 <= io_in_r_bypass_11_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_2_load_store_15 <= io_in_r_bypass_11_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_2_df_is_ws_15 <= io_in_r_bypass_11_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_2_stall_15 <= io_in_r_bypass_11_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_3_data_15 <= io_in_r_bypass_11_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_3_load_store_15 <= io_in_r_bypass_11_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_3_df_is_ws_15 <= io_in_r_bypass_11_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_3_stall_15 <= io_in_r_bypass_11_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_0_data_15 <= io_in_r_bypass_12_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_0_load_store_15 <= io_in_r_bypass_12_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_0_df_is_ws_15 <= io_in_r_bypass_12_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_0_stall_15 <= io_in_r_bypass_12_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_1_data_15 <= io_in_r_bypass_12_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_1_load_store_15 <= io_in_r_bypass_12_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_1_df_is_ws_15 <= io_in_r_bypass_12_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_1_stall_15 <= io_in_r_bypass_12_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_2_data_15 <= io_in_r_bypass_12_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_2_load_store_15 <= io_in_r_bypass_12_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_2_df_is_ws_15 <= io_in_r_bypass_12_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_2_stall_15 <= io_in_r_bypass_12_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_3_data_15 <= io_in_r_bypass_12_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_3_load_store_15 <= io_in_r_bypass_12_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_3_df_is_ws_15 <= io_in_r_bypass_12_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_3_stall_15 <= io_in_r_bypass_12_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_0_data_15 <= io_in_r_bypass_13_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_0_load_store_15 <= io_in_r_bypass_13_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_0_df_is_ws_15 <= io_in_r_bypass_13_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_0_stall_15 <= io_in_r_bypass_13_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_1_data_15 <= io_in_r_bypass_13_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_1_load_store_15 <= io_in_r_bypass_13_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_1_df_is_ws_15 <= io_in_r_bypass_13_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_1_stall_15 <= io_in_r_bypass_13_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_2_data_15 <= io_in_r_bypass_13_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_2_load_store_15 <= io_in_r_bypass_13_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_2_df_is_ws_15 <= io_in_r_bypass_13_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_2_stall_15 <= io_in_r_bypass_13_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_3_data_15 <= io_in_r_bypass_13_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_3_load_store_15 <= io_in_r_bypass_13_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_3_df_is_ws_15 <= io_in_r_bypass_13_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_3_stall_15 <= io_in_r_bypass_13_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_0_data_15 <= io_in_r_bypass_14_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_0_load_store_15 <= io_in_r_bypass_14_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_0_df_is_ws_15 <= io_in_r_bypass_14_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_0_stall_15 <= io_in_r_bypass_14_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_1_data_15 <= io_in_r_bypass_14_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_1_load_store_15 <= io_in_r_bypass_14_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_1_df_is_ws_15 <= io_in_r_bypass_14_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_1_stall_15 <= io_in_r_bypass_14_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_2_data_15 <= io_in_r_bypass_14_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_2_load_store_15 <= io_in_r_bypass_14_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_2_df_is_ws_15 <= io_in_r_bypass_14_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_2_stall_15 <= io_in_r_bypass_14_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_3_data_15 <= io_in_r_bypass_14_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_3_load_store_15 <= io_in_r_bypass_14_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_3_df_is_ws_15 <= io_in_r_bypass_14_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_3_stall_15 <= io_in_r_bypass_14_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_0_data_15 <= io_in_r_bypass_15_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_0_load_store_15 <= io_in_r_bypass_15_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_0_df_is_ws_15 <= io_in_r_bypass_15_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_0_stall_15 <= io_in_r_bypass_15_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_1_data_15 <= io_in_r_bypass_15_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_1_load_store_15 <= io_in_r_bypass_15_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_1_df_is_ws_15 <= io_in_r_bypass_15_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_1_stall_15 <= io_in_r_bypass_15_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_2_data_15 <= io_in_r_bypass_15_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_2_load_store_15 <= io_in_r_bypass_15_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_2_df_is_ws_15 <= io_in_r_bypass_15_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_2_stall_15 <= io_in_r_bypass_15_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_3_data_15 <= io_in_r_bypass_15_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_3_load_store_15 <= io_in_r_bypass_15_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_3_df_is_ws_15 <= io_in_r_bypass_15_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_3_stall_15 <= io_in_r_bypass_15_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_0_data_15 <= io_in_r_bypass_16_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_0_load_store_15 <= io_in_r_bypass_16_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_0_df_is_ws_15 <= io_in_r_bypass_16_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_0_stall_15 <= io_in_r_bypass_16_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_1_data_15 <= io_in_r_bypass_16_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_1_load_store_15 <= io_in_r_bypass_16_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_1_df_is_ws_15 <= io_in_r_bypass_16_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_1_stall_15 <= io_in_r_bypass_16_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_2_data_15 <= io_in_r_bypass_16_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_2_load_store_15 <= io_in_r_bypass_16_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_2_df_is_ws_15 <= io_in_r_bypass_16_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_2_stall_15 <= io_in_r_bypass_16_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_3_data_15 <= io_in_r_bypass_16_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_3_load_store_15 <= io_in_r_bypass_16_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_3_df_is_ws_15 <= io_in_r_bypass_16_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_3_stall_15 <= io_in_r_bypass_16_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_0_data_15 <= io_in_r_bypass_17_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_0_load_store_15 <= io_in_r_bypass_17_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_0_df_is_ws_15 <= io_in_r_bypass_17_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_0_stall_15 <= io_in_r_bypass_17_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_1_data_15 <= io_in_r_bypass_17_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_1_load_store_15 <= io_in_r_bypass_17_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_1_df_is_ws_15 <= io_in_r_bypass_17_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_1_stall_15 <= io_in_r_bypass_17_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_2_data_15 <= io_in_r_bypass_17_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_2_load_store_15 <= io_in_r_bypass_17_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_2_df_is_ws_15 <= io_in_r_bypass_17_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_2_stall_15 <= io_in_r_bypass_17_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_3_data_15 <= io_in_r_bypass_17_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_3_load_store_15 <= io_in_r_bypass_17_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_3_df_is_ws_15 <= io_in_r_bypass_17_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_3_stall_15 <= io_in_r_bypass_17_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_0_data_15 <= io_in_r_bypass_18_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_0_load_store_15 <= io_in_r_bypass_18_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_0_df_is_ws_15 <= io_in_r_bypass_18_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_0_stall_15 <= io_in_r_bypass_18_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_1_data_15 <= io_in_r_bypass_18_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_1_load_store_15 <= io_in_r_bypass_18_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_1_df_is_ws_15 <= io_in_r_bypass_18_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_1_stall_15 <= io_in_r_bypass_18_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_2_data_15 <= io_in_r_bypass_18_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_2_load_store_15 <= io_in_r_bypass_18_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_2_df_is_ws_15 <= io_in_r_bypass_18_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_2_stall_15 <= io_in_r_bypass_18_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_3_data_15 <= io_in_r_bypass_18_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_3_load_store_15 <= io_in_r_bypass_18_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_3_df_is_ws_15 <= io_in_r_bypass_18_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_3_stall_15 <= io_in_r_bypass_18_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_0_data_15 <= io_in_r_bypass_19_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_0_load_store_15 <= io_in_r_bypass_19_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_0_df_is_ws_15 <= io_in_r_bypass_19_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_0_stall_15 <= io_in_r_bypass_19_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_1_data_15 <= io_in_r_bypass_19_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_1_load_store_15 <= io_in_r_bypass_19_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_1_df_is_ws_15 <= io_in_r_bypass_19_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_1_stall_15 <= io_in_r_bypass_19_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_2_data_15 <= io_in_r_bypass_19_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_2_load_store_15 <= io_in_r_bypass_19_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_2_df_is_ws_15 <= io_in_r_bypass_19_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_2_stall_15 <= io_in_r_bypass_19_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_3_data_15 <= io_in_r_bypass_19_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_3_load_store_15 <= io_in_r_bypass_19_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_3_df_is_ws_15 <= io_in_r_bypass_19_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_3_stall_15 <= io_in_r_bypass_19_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_0_data_15 <= io_in_r_bypass_20_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_0_load_store_15 <= io_in_r_bypass_20_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_0_df_is_ws_15 <= io_in_r_bypass_20_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_0_stall_15 <= io_in_r_bypass_20_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_1_data_15 <= io_in_r_bypass_20_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_1_load_store_15 <= io_in_r_bypass_20_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_1_df_is_ws_15 <= io_in_r_bypass_20_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_1_stall_15 <= io_in_r_bypass_20_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_2_data_15 <= io_in_r_bypass_20_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_2_load_store_15 <= io_in_r_bypass_20_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_2_df_is_ws_15 <= io_in_r_bypass_20_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_2_stall_15 <= io_in_r_bypass_20_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_3_data_15 <= io_in_r_bypass_20_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_3_load_store_15 <= io_in_r_bypass_20_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_3_df_is_ws_15 <= io_in_r_bypass_20_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_3_stall_15 <= io_in_r_bypass_20_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_0_data_15 <= io_in_r_bypass_21_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_0_load_store_15 <= io_in_r_bypass_21_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_0_df_is_ws_15 <= io_in_r_bypass_21_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_0_stall_15 <= io_in_r_bypass_21_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_1_data_15 <= io_in_r_bypass_21_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_1_load_store_15 <= io_in_r_bypass_21_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_1_df_is_ws_15 <= io_in_r_bypass_21_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_1_stall_15 <= io_in_r_bypass_21_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_2_data_15 <= io_in_r_bypass_21_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_2_load_store_15 <= io_in_r_bypass_21_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_2_df_is_ws_15 <= io_in_r_bypass_21_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_2_stall_15 <= io_in_r_bypass_21_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_3_data_15 <= io_in_r_bypass_21_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_3_load_store_15 <= io_in_r_bypass_21_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_3_df_is_ws_15 <= io_in_r_bypass_21_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_3_stall_15 <= io_in_r_bypass_21_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_0_data_15 <= io_in_r_bypass_22_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_0_load_store_15 <= io_in_r_bypass_22_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_0_df_is_ws_15 <= io_in_r_bypass_22_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_0_stall_15 <= io_in_r_bypass_22_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_1_data_15 <= io_in_r_bypass_22_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_1_load_store_15 <= io_in_r_bypass_22_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_1_df_is_ws_15 <= io_in_r_bypass_22_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_1_stall_15 <= io_in_r_bypass_22_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_2_data_15 <= io_in_r_bypass_22_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_2_load_store_15 <= io_in_r_bypass_22_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_2_df_is_ws_15 <= io_in_r_bypass_22_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_2_stall_15 <= io_in_r_bypass_22_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_3_data_15 <= io_in_r_bypass_22_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_3_load_store_15 <= io_in_r_bypass_22_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_3_df_is_ws_15 <= io_in_r_bypass_22_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_3_stall_15 <= io_in_r_bypass_22_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_0_data_15 <= io_in_r_bypass_23_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_0_load_store_15 <= io_in_r_bypass_23_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_0_df_is_ws_15 <= io_in_r_bypass_23_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_0_stall_15 <= io_in_r_bypass_23_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_1_data_15 <= io_in_r_bypass_23_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_1_load_store_15 <= io_in_r_bypass_23_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_1_df_is_ws_15 <= io_in_r_bypass_23_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_1_stall_15 <= io_in_r_bypass_23_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_2_data_15 <= io_in_r_bypass_23_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_2_load_store_15 <= io_in_r_bypass_23_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_2_df_is_ws_15 <= io_in_r_bypass_23_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_2_stall_15 <= io_in_r_bypass_23_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_3_data_15 <= io_in_r_bypass_23_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_3_load_store_15 <= io_in_r_bypass_23_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_3_df_is_ws_15 <= io_in_r_bypass_23_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_3_stall_15 <= io_in_r_bypass_23_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_0_data_15 <= io_in_r_bypass_24_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_0_load_store_15 <= io_in_r_bypass_24_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_0_df_is_ws_15 <= io_in_r_bypass_24_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_0_stall_15 <= io_in_r_bypass_24_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_1_data_15 <= io_in_r_bypass_24_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_1_load_store_15 <= io_in_r_bypass_24_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_1_df_is_ws_15 <= io_in_r_bypass_24_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_1_stall_15 <= io_in_r_bypass_24_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_2_data_15 <= io_in_r_bypass_24_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_2_load_store_15 <= io_in_r_bypass_24_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_2_df_is_ws_15 <= io_in_r_bypass_24_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_2_stall_15 <= io_in_r_bypass_24_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_3_data_15 <= io_in_r_bypass_24_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_3_load_store_15 <= io_in_r_bypass_24_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_3_df_is_ws_15 <= io_in_r_bypass_24_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_3_stall_15 <= io_in_r_bypass_24_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_0_data_15 <= io_in_r_bypass_25_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_0_load_store_15 <= io_in_r_bypass_25_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_0_df_is_ws_15 <= io_in_r_bypass_25_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_0_stall_15 <= io_in_r_bypass_25_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_1_data_15 <= io_in_r_bypass_25_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_1_load_store_15 <= io_in_r_bypass_25_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_1_df_is_ws_15 <= io_in_r_bypass_25_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_1_stall_15 <= io_in_r_bypass_25_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_2_data_15 <= io_in_r_bypass_25_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_2_load_store_15 <= io_in_r_bypass_25_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_2_df_is_ws_15 <= io_in_r_bypass_25_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_2_stall_15 <= io_in_r_bypass_25_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_3_data_15 <= io_in_r_bypass_25_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_3_load_store_15 <= io_in_r_bypass_25_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_3_df_is_ws_15 <= io_in_r_bypass_25_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_3_stall_15 <= io_in_r_bypass_25_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_0_data_15 <= io_in_r_bypass_26_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_0_load_store_15 <= io_in_r_bypass_26_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_0_df_is_ws_15 <= io_in_r_bypass_26_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_0_stall_15 <= io_in_r_bypass_26_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_1_data_15 <= io_in_r_bypass_26_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_1_load_store_15 <= io_in_r_bypass_26_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_1_df_is_ws_15 <= io_in_r_bypass_26_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_1_stall_15 <= io_in_r_bypass_26_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_2_data_15 <= io_in_r_bypass_26_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_2_load_store_15 <= io_in_r_bypass_26_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_2_df_is_ws_15 <= io_in_r_bypass_26_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_2_stall_15 <= io_in_r_bypass_26_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_3_data_15 <= io_in_r_bypass_26_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_3_load_store_15 <= io_in_r_bypass_26_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_3_df_is_ws_15 <= io_in_r_bypass_26_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_3_stall_15 <= io_in_r_bypass_26_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_0_data_15 <= io_in_r_bypass_27_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_0_load_store_15 <= io_in_r_bypass_27_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_0_df_is_ws_15 <= io_in_r_bypass_27_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_0_stall_15 <= io_in_r_bypass_27_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_1_data_15 <= io_in_r_bypass_27_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_1_load_store_15 <= io_in_r_bypass_27_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_1_df_is_ws_15 <= io_in_r_bypass_27_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_1_stall_15 <= io_in_r_bypass_27_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_2_data_15 <= io_in_r_bypass_27_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_2_load_store_15 <= io_in_r_bypass_27_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_2_df_is_ws_15 <= io_in_r_bypass_27_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_2_stall_15 <= io_in_r_bypass_27_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_3_data_15 <= io_in_r_bypass_27_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_3_load_store_15 <= io_in_r_bypass_27_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_3_df_is_ws_15 <= io_in_r_bypass_27_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_3_stall_15 <= io_in_r_bypass_27_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_0_data_15 <= io_in_r_bypass_28_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_0_load_store_15 <= io_in_r_bypass_28_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_0_df_is_ws_15 <= io_in_r_bypass_28_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_0_stall_15 <= io_in_r_bypass_28_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_1_data_15 <= io_in_r_bypass_28_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_1_load_store_15 <= io_in_r_bypass_28_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_1_df_is_ws_15 <= io_in_r_bypass_28_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_1_stall_15 <= io_in_r_bypass_28_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_2_data_15 <= io_in_r_bypass_28_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_2_load_store_15 <= io_in_r_bypass_28_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_2_df_is_ws_15 <= io_in_r_bypass_28_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_2_stall_15 <= io_in_r_bypass_28_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_3_data_15 <= io_in_r_bypass_28_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_3_load_store_15 <= io_in_r_bypass_28_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_3_df_is_ws_15 <= io_in_r_bypass_28_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_3_stall_15 <= io_in_r_bypass_28_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_0_data_15 <= io_in_r_bypass_29_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_0_load_store_15 <= io_in_r_bypass_29_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_0_df_is_ws_15 <= io_in_r_bypass_29_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_0_stall_15 <= io_in_r_bypass_29_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_1_data_15 <= io_in_r_bypass_29_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_1_load_store_15 <= io_in_r_bypass_29_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_1_df_is_ws_15 <= io_in_r_bypass_29_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_1_stall_15 <= io_in_r_bypass_29_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_2_data_15 <= io_in_r_bypass_29_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_2_load_store_15 <= io_in_r_bypass_29_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_2_df_is_ws_15 <= io_in_r_bypass_29_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_2_stall_15 <= io_in_r_bypass_29_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_3_data_15 <= io_in_r_bypass_29_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_3_load_store_15 <= io_in_r_bypass_29_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_3_df_is_ws_15 <= io_in_r_bypass_29_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_3_stall_15 <= io_in_r_bypass_29_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_0_data_15 <= io_in_r_bypass_30_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_0_load_store_15 <= io_in_r_bypass_30_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_0_df_is_ws_15 <= io_in_r_bypass_30_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_0_stall_15 <= io_in_r_bypass_30_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_1_data_15 <= io_in_r_bypass_30_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_1_load_store_15 <= io_in_r_bypass_30_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_1_df_is_ws_15 <= io_in_r_bypass_30_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_1_stall_15 <= io_in_r_bypass_30_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_2_data_15 <= io_in_r_bypass_30_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_2_load_store_15 <= io_in_r_bypass_30_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_2_df_is_ws_15 <= io_in_r_bypass_30_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_2_stall_15 <= io_in_r_bypass_30_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_3_data_15 <= io_in_r_bypass_30_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_3_load_store_15 <= io_in_r_bypass_30_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_3_df_is_ws_15 <= io_in_r_bypass_30_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_3_stall_15 <= io_in_r_bypass_30_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_0_data_15 <= io_in_r_bypass_31_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_0_load_store_15 <= io_in_r_bypass_31_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_0_df_is_ws_15 <= io_in_r_bypass_31_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_0_stall_15 <= io_in_r_bypass_31_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_1_data_15 <= io_in_r_bypass_31_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_1_load_store_15 <= io_in_r_bypass_31_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_1_df_is_ws_15 <= io_in_r_bypass_31_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_1_stall_15 <= io_in_r_bypass_31_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_2_data_15 <= io_in_r_bypass_31_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_2_load_store_15 <= io_in_r_bypass_31_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_2_df_is_ws_15 <= io_in_r_bypass_31_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_2_stall_15 <= io_in_r_bypass_31_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_3_data_15 <= io_in_r_bypass_31_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_3_load_store_15 <= io_in_r_bypass_31_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_3_df_is_ws_15 <= io_in_r_bypass_31_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_3_stall_15 <= io_in_r_bypass_31_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_0_data_16 <= io_in_r_bypass_0_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_0_load_store_16 <= io_in_r_bypass_0_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_0_df_is_ws_16 <= io_in_r_bypass_0_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_0_stall_16 <= io_in_r_bypass_0_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_1_data_16 <= io_in_r_bypass_0_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_1_load_store_16 <= io_in_r_bypass_0_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_1_df_is_ws_16 <= io_in_r_bypass_0_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_1_stall_16 <= io_in_r_bypass_0_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_2_data_16 <= io_in_r_bypass_0_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_2_load_store_16 <= io_in_r_bypass_0_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_2_df_is_ws_16 <= io_in_r_bypass_0_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_2_stall_16 <= io_in_r_bypass_0_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_3_data_16 <= io_in_r_bypass_0_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_3_load_store_16 <= io_in_r_bypass_0_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_3_df_is_ws_16 <= io_in_r_bypass_0_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_3_stall_16 <= io_in_r_bypass_0_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_0_data_16 <= io_in_r_bypass_1_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_0_load_store_16 <= io_in_r_bypass_1_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_0_df_is_ws_16 <= io_in_r_bypass_1_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_0_stall_16 <= io_in_r_bypass_1_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_1_data_16 <= io_in_r_bypass_1_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_1_load_store_16 <= io_in_r_bypass_1_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_1_df_is_ws_16 <= io_in_r_bypass_1_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_1_stall_16 <= io_in_r_bypass_1_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_2_data_16 <= io_in_r_bypass_1_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_2_load_store_16 <= io_in_r_bypass_1_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_2_df_is_ws_16 <= io_in_r_bypass_1_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_2_stall_16 <= io_in_r_bypass_1_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_3_data_16 <= io_in_r_bypass_1_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_3_load_store_16 <= io_in_r_bypass_1_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_3_df_is_ws_16 <= io_in_r_bypass_1_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_3_stall_16 <= io_in_r_bypass_1_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_0_data_16 <= io_in_r_bypass_2_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_0_load_store_16 <= io_in_r_bypass_2_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_0_df_is_ws_16 <= io_in_r_bypass_2_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_0_stall_16 <= io_in_r_bypass_2_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_1_data_16 <= io_in_r_bypass_2_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_1_load_store_16 <= io_in_r_bypass_2_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_1_df_is_ws_16 <= io_in_r_bypass_2_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_1_stall_16 <= io_in_r_bypass_2_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_2_data_16 <= io_in_r_bypass_2_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_2_load_store_16 <= io_in_r_bypass_2_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_2_df_is_ws_16 <= io_in_r_bypass_2_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_2_stall_16 <= io_in_r_bypass_2_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_3_data_16 <= io_in_r_bypass_2_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_3_load_store_16 <= io_in_r_bypass_2_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_3_df_is_ws_16 <= io_in_r_bypass_2_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_3_stall_16 <= io_in_r_bypass_2_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_0_data_16 <= io_in_r_bypass_3_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_0_load_store_16 <= io_in_r_bypass_3_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_0_df_is_ws_16 <= io_in_r_bypass_3_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_0_stall_16 <= io_in_r_bypass_3_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_1_data_16 <= io_in_r_bypass_3_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_1_load_store_16 <= io_in_r_bypass_3_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_1_df_is_ws_16 <= io_in_r_bypass_3_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_1_stall_16 <= io_in_r_bypass_3_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_2_data_16 <= io_in_r_bypass_3_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_2_load_store_16 <= io_in_r_bypass_3_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_2_df_is_ws_16 <= io_in_r_bypass_3_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_2_stall_16 <= io_in_r_bypass_3_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_3_data_16 <= io_in_r_bypass_3_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_3_load_store_16 <= io_in_r_bypass_3_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_3_df_is_ws_16 <= io_in_r_bypass_3_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_3_stall_16 <= io_in_r_bypass_3_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_0_data_16 <= io_in_r_bypass_4_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_0_load_store_16 <= io_in_r_bypass_4_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_0_df_is_ws_16 <= io_in_r_bypass_4_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_0_stall_16 <= io_in_r_bypass_4_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_1_data_16 <= io_in_r_bypass_4_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_1_load_store_16 <= io_in_r_bypass_4_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_1_df_is_ws_16 <= io_in_r_bypass_4_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_1_stall_16 <= io_in_r_bypass_4_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_2_data_16 <= io_in_r_bypass_4_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_2_load_store_16 <= io_in_r_bypass_4_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_2_df_is_ws_16 <= io_in_r_bypass_4_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_2_stall_16 <= io_in_r_bypass_4_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_3_data_16 <= io_in_r_bypass_4_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_3_load_store_16 <= io_in_r_bypass_4_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_3_df_is_ws_16 <= io_in_r_bypass_4_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_3_stall_16 <= io_in_r_bypass_4_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_0_data_16 <= io_in_r_bypass_5_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_0_load_store_16 <= io_in_r_bypass_5_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_0_df_is_ws_16 <= io_in_r_bypass_5_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_0_stall_16 <= io_in_r_bypass_5_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_1_data_16 <= io_in_r_bypass_5_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_1_load_store_16 <= io_in_r_bypass_5_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_1_df_is_ws_16 <= io_in_r_bypass_5_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_1_stall_16 <= io_in_r_bypass_5_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_2_data_16 <= io_in_r_bypass_5_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_2_load_store_16 <= io_in_r_bypass_5_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_2_df_is_ws_16 <= io_in_r_bypass_5_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_2_stall_16 <= io_in_r_bypass_5_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_3_data_16 <= io_in_r_bypass_5_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_3_load_store_16 <= io_in_r_bypass_5_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_3_df_is_ws_16 <= io_in_r_bypass_5_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_3_stall_16 <= io_in_r_bypass_5_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_0_data_16 <= io_in_r_bypass_6_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_0_load_store_16 <= io_in_r_bypass_6_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_0_df_is_ws_16 <= io_in_r_bypass_6_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_0_stall_16 <= io_in_r_bypass_6_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_1_data_16 <= io_in_r_bypass_6_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_1_load_store_16 <= io_in_r_bypass_6_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_1_df_is_ws_16 <= io_in_r_bypass_6_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_1_stall_16 <= io_in_r_bypass_6_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_2_data_16 <= io_in_r_bypass_6_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_2_load_store_16 <= io_in_r_bypass_6_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_2_df_is_ws_16 <= io_in_r_bypass_6_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_2_stall_16 <= io_in_r_bypass_6_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_3_data_16 <= io_in_r_bypass_6_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_3_load_store_16 <= io_in_r_bypass_6_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_3_df_is_ws_16 <= io_in_r_bypass_6_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_3_stall_16 <= io_in_r_bypass_6_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_0_data_16 <= io_in_r_bypass_7_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_0_load_store_16 <= io_in_r_bypass_7_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_0_df_is_ws_16 <= io_in_r_bypass_7_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_0_stall_16 <= io_in_r_bypass_7_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_1_data_16 <= io_in_r_bypass_7_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_1_load_store_16 <= io_in_r_bypass_7_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_1_df_is_ws_16 <= io_in_r_bypass_7_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_1_stall_16 <= io_in_r_bypass_7_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_2_data_16 <= io_in_r_bypass_7_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_2_load_store_16 <= io_in_r_bypass_7_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_2_df_is_ws_16 <= io_in_r_bypass_7_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_2_stall_16 <= io_in_r_bypass_7_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_3_data_16 <= io_in_r_bypass_7_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_3_load_store_16 <= io_in_r_bypass_7_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_3_df_is_ws_16 <= io_in_r_bypass_7_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_3_stall_16 <= io_in_r_bypass_7_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_0_data_16 <= io_in_r_bypass_8_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_0_load_store_16 <= io_in_r_bypass_8_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_0_df_is_ws_16 <= io_in_r_bypass_8_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_0_stall_16 <= io_in_r_bypass_8_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_1_data_16 <= io_in_r_bypass_8_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_1_load_store_16 <= io_in_r_bypass_8_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_1_df_is_ws_16 <= io_in_r_bypass_8_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_1_stall_16 <= io_in_r_bypass_8_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_2_data_16 <= io_in_r_bypass_8_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_2_load_store_16 <= io_in_r_bypass_8_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_2_df_is_ws_16 <= io_in_r_bypass_8_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_2_stall_16 <= io_in_r_bypass_8_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_3_data_16 <= io_in_r_bypass_8_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_3_load_store_16 <= io_in_r_bypass_8_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_3_df_is_ws_16 <= io_in_r_bypass_8_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_3_stall_16 <= io_in_r_bypass_8_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_0_data_16 <= io_in_r_bypass_9_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_0_load_store_16 <= io_in_r_bypass_9_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_0_df_is_ws_16 <= io_in_r_bypass_9_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_0_stall_16 <= io_in_r_bypass_9_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_1_data_16 <= io_in_r_bypass_9_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_1_load_store_16 <= io_in_r_bypass_9_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_1_df_is_ws_16 <= io_in_r_bypass_9_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_1_stall_16 <= io_in_r_bypass_9_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_2_data_16 <= io_in_r_bypass_9_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_2_load_store_16 <= io_in_r_bypass_9_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_2_df_is_ws_16 <= io_in_r_bypass_9_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_2_stall_16 <= io_in_r_bypass_9_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_3_data_16 <= io_in_r_bypass_9_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_3_load_store_16 <= io_in_r_bypass_9_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_3_df_is_ws_16 <= io_in_r_bypass_9_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_3_stall_16 <= io_in_r_bypass_9_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_0_data_16 <= io_in_r_bypass_10_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_0_load_store_16 <= io_in_r_bypass_10_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_0_df_is_ws_16 <= io_in_r_bypass_10_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_0_stall_16 <= io_in_r_bypass_10_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_1_data_16 <= io_in_r_bypass_10_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_1_load_store_16 <= io_in_r_bypass_10_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_1_df_is_ws_16 <= io_in_r_bypass_10_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_1_stall_16 <= io_in_r_bypass_10_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_2_data_16 <= io_in_r_bypass_10_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_2_load_store_16 <= io_in_r_bypass_10_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_2_df_is_ws_16 <= io_in_r_bypass_10_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_2_stall_16 <= io_in_r_bypass_10_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_3_data_16 <= io_in_r_bypass_10_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_3_load_store_16 <= io_in_r_bypass_10_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_3_df_is_ws_16 <= io_in_r_bypass_10_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_3_stall_16 <= io_in_r_bypass_10_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_0_data_16 <= io_in_r_bypass_11_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_0_load_store_16 <= io_in_r_bypass_11_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_0_df_is_ws_16 <= io_in_r_bypass_11_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_0_stall_16 <= io_in_r_bypass_11_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_1_data_16 <= io_in_r_bypass_11_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_1_load_store_16 <= io_in_r_bypass_11_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_1_df_is_ws_16 <= io_in_r_bypass_11_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_1_stall_16 <= io_in_r_bypass_11_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_2_data_16 <= io_in_r_bypass_11_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_2_load_store_16 <= io_in_r_bypass_11_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_2_df_is_ws_16 <= io_in_r_bypass_11_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_2_stall_16 <= io_in_r_bypass_11_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_3_data_16 <= io_in_r_bypass_11_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_3_load_store_16 <= io_in_r_bypass_11_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_3_df_is_ws_16 <= io_in_r_bypass_11_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_3_stall_16 <= io_in_r_bypass_11_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_0_data_16 <= io_in_r_bypass_12_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_0_load_store_16 <= io_in_r_bypass_12_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_0_df_is_ws_16 <= io_in_r_bypass_12_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_0_stall_16 <= io_in_r_bypass_12_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_1_data_16 <= io_in_r_bypass_12_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_1_load_store_16 <= io_in_r_bypass_12_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_1_df_is_ws_16 <= io_in_r_bypass_12_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_1_stall_16 <= io_in_r_bypass_12_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_2_data_16 <= io_in_r_bypass_12_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_2_load_store_16 <= io_in_r_bypass_12_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_2_df_is_ws_16 <= io_in_r_bypass_12_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_2_stall_16 <= io_in_r_bypass_12_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_3_data_16 <= io_in_r_bypass_12_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_3_load_store_16 <= io_in_r_bypass_12_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_3_df_is_ws_16 <= io_in_r_bypass_12_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_3_stall_16 <= io_in_r_bypass_12_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_0_data_16 <= io_in_r_bypass_13_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_0_load_store_16 <= io_in_r_bypass_13_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_0_df_is_ws_16 <= io_in_r_bypass_13_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_0_stall_16 <= io_in_r_bypass_13_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_1_data_16 <= io_in_r_bypass_13_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_1_load_store_16 <= io_in_r_bypass_13_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_1_df_is_ws_16 <= io_in_r_bypass_13_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_1_stall_16 <= io_in_r_bypass_13_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_2_data_16 <= io_in_r_bypass_13_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_2_load_store_16 <= io_in_r_bypass_13_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_2_df_is_ws_16 <= io_in_r_bypass_13_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_2_stall_16 <= io_in_r_bypass_13_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_3_data_16 <= io_in_r_bypass_13_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_3_load_store_16 <= io_in_r_bypass_13_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_3_df_is_ws_16 <= io_in_r_bypass_13_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_3_stall_16 <= io_in_r_bypass_13_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_0_data_16 <= io_in_r_bypass_14_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_0_load_store_16 <= io_in_r_bypass_14_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_0_df_is_ws_16 <= io_in_r_bypass_14_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_0_stall_16 <= io_in_r_bypass_14_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_1_data_16 <= io_in_r_bypass_14_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_1_load_store_16 <= io_in_r_bypass_14_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_1_df_is_ws_16 <= io_in_r_bypass_14_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_1_stall_16 <= io_in_r_bypass_14_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_2_data_16 <= io_in_r_bypass_14_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_2_load_store_16 <= io_in_r_bypass_14_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_2_df_is_ws_16 <= io_in_r_bypass_14_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_2_stall_16 <= io_in_r_bypass_14_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_3_data_16 <= io_in_r_bypass_14_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_3_load_store_16 <= io_in_r_bypass_14_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_3_df_is_ws_16 <= io_in_r_bypass_14_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_3_stall_16 <= io_in_r_bypass_14_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_0_data_16 <= io_in_r_bypass_15_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_0_load_store_16 <= io_in_r_bypass_15_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_0_df_is_ws_16 <= io_in_r_bypass_15_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_0_stall_16 <= io_in_r_bypass_15_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_1_data_16 <= io_in_r_bypass_15_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_1_load_store_16 <= io_in_r_bypass_15_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_1_df_is_ws_16 <= io_in_r_bypass_15_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_1_stall_16 <= io_in_r_bypass_15_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_2_data_16 <= io_in_r_bypass_15_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_2_load_store_16 <= io_in_r_bypass_15_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_2_df_is_ws_16 <= io_in_r_bypass_15_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_2_stall_16 <= io_in_r_bypass_15_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_3_data_16 <= io_in_r_bypass_15_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_3_load_store_16 <= io_in_r_bypass_15_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_3_df_is_ws_16 <= io_in_r_bypass_15_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_3_stall_16 <= io_in_r_bypass_15_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_0_data_16 <= io_in_r_bypass_16_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_0_load_store_16 <= io_in_r_bypass_16_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_0_df_is_ws_16 <= io_in_r_bypass_16_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_0_stall_16 <= io_in_r_bypass_16_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_1_data_16 <= io_in_r_bypass_16_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_1_load_store_16 <= io_in_r_bypass_16_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_1_df_is_ws_16 <= io_in_r_bypass_16_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_1_stall_16 <= io_in_r_bypass_16_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_2_data_16 <= io_in_r_bypass_16_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_2_load_store_16 <= io_in_r_bypass_16_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_2_df_is_ws_16 <= io_in_r_bypass_16_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_2_stall_16 <= io_in_r_bypass_16_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_3_data_16 <= io_in_r_bypass_16_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_3_load_store_16 <= io_in_r_bypass_16_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_3_df_is_ws_16 <= io_in_r_bypass_16_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_3_stall_16 <= io_in_r_bypass_16_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_0_data_16 <= io_in_r_bypass_17_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_0_load_store_16 <= io_in_r_bypass_17_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_0_df_is_ws_16 <= io_in_r_bypass_17_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_0_stall_16 <= io_in_r_bypass_17_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_1_data_16 <= io_in_r_bypass_17_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_1_load_store_16 <= io_in_r_bypass_17_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_1_df_is_ws_16 <= io_in_r_bypass_17_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_1_stall_16 <= io_in_r_bypass_17_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_2_data_16 <= io_in_r_bypass_17_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_2_load_store_16 <= io_in_r_bypass_17_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_2_df_is_ws_16 <= io_in_r_bypass_17_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_2_stall_16 <= io_in_r_bypass_17_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_3_data_16 <= io_in_r_bypass_17_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_3_load_store_16 <= io_in_r_bypass_17_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_3_df_is_ws_16 <= io_in_r_bypass_17_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_3_stall_16 <= io_in_r_bypass_17_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_0_data_16 <= io_in_r_bypass_18_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_0_load_store_16 <= io_in_r_bypass_18_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_0_df_is_ws_16 <= io_in_r_bypass_18_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_0_stall_16 <= io_in_r_bypass_18_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_1_data_16 <= io_in_r_bypass_18_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_1_load_store_16 <= io_in_r_bypass_18_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_1_df_is_ws_16 <= io_in_r_bypass_18_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_1_stall_16 <= io_in_r_bypass_18_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_2_data_16 <= io_in_r_bypass_18_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_2_load_store_16 <= io_in_r_bypass_18_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_2_df_is_ws_16 <= io_in_r_bypass_18_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_2_stall_16 <= io_in_r_bypass_18_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_3_data_16 <= io_in_r_bypass_18_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_3_load_store_16 <= io_in_r_bypass_18_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_3_df_is_ws_16 <= io_in_r_bypass_18_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_3_stall_16 <= io_in_r_bypass_18_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_0_data_16 <= io_in_r_bypass_19_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_0_load_store_16 <= io_in_r_bypass_19_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_0_df_is_ws_16 <= io_in_r_bypass_19_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_0_stall_16 <= io_in_r_bypass_19_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_1_data_16 <= io_in_r_bypass_19_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_1_load_store_16 <= io_in_r_bypass_19_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_1_df_is_ws_16 <= io_in_r_bypass_19_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_1_stall_16 <= io_in_r_bypass_19_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_2_data_16 <= io_in_r_bypass_19_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_2_load_store_16 <= io_in_r_bypass_19_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_2_df_is_ws_16 <= io_in_r_bypass_19_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_2_stall_16 <= io_in_r_bypass_19_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_3_data_16 <= io_in_r_bypass_19_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_3_load_store_16 <= io_in_r_bypass_19_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_3_df_is_ws_16 <= io_in_r_bypass_19_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_3_stall_16 <= io_in_r_bypass_19_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_0_data_16 <= io_in_r_bypass_20_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_0_load_store_16 <= io_in_r_bypass_20_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_0_df_is_ws_16 <= io_in_r_bypass_20_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_0_stall_16 <= io_in_r_bypass_20_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_1_data_16 <= io_in_r_bypass_20_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_1_load_store_16 <= io_in_r_bypass_20_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_1_df_is_ws_16 <= io_in_r_bypass_20_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_1_stall_16 <= io_in_r_bypass_20_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_2_data_16 <= io_in_r_bypass_20_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_2_load_store_16 <= io_in_r_bypass_20_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_2_df_is_ws_16 <= io_in_r_bypass_20_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_2_stall_16 <= io_in_r_bypass_20_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_3_data_16 <= io_in_r_bypass_20_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_3_load_store_16 <= io_in_r_bypass_20_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_3_df_is_ws_16 <= io_in_r_bypass_20_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_3_stall_16 <= io_in_r_bypass_20_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_0_data_16 <= io_in_r_bypass_21_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_0_load_store_16 <= io_in_r_bypass_21_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_0_df_is_ws_16 <= io_in_r_bypass_21_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_0_stall_16 <= io_in_r_bypass_21_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_1_data_16 <= io_in_r_bypass_21_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_1_load_store_16 <= io_in_r_bypass_21_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_1_df_is_ws_16 <= io_in_r_bypass_21_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_1_stall_16 <= io_in_r_bypass_21_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_2_data_16 <= io_in_r_bypass_21_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_2_load_store_16 <= io_in_r_bypass_21_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_2_df_is_ws_16 <= io_in_r_bypass_21_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_2_stall_16 <= io_in_r_bypass_21_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_3_data_16 <= io_in_r_bypass_21_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_3_load_store_16 <= io_in_r_bypass_21_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_3_df_is_ws_16 <= io_in_r_bypass_21_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_3_stall_16 <= io_in_r_bypass_21_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_0_data_16 <= io_in_r_bypass_22_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_0_load_store_16 <= io_in_r_bypass_22_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_0_df_is_ws_16 <= io_in_r_bypass_22_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_0_stall_16 <= io_in_r_bypass_22_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_1_data_16 <= io_in_r_bypass_22_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_1_load_store_16 <= io_in_r_bypass_22_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_1_df_is_ws_16 <= io_in_r_bypass_22_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_1_stall_16 <= io_in_r_bypass_22_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_2_data_16 <= io_in_r_bypass_22_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_2_load_store_16 <= io_in_r_bypass_22_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_2_df_is_ws_16 <= io_in_r_bypass_22_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_2_stall_16 <= io_in_r_bypass_22_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_3_data_16 <= io_in_r_bypass_22_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_3_load_store_16 <= io_in_r_bypass_22_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_3_df_is_ws_16 <= io_in_r_bypass_22_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_3_stall_16 <= io_in_r_bypass_22_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_0_data_16 <= io_in_r_bypass_23_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_0_load_store_16 <= io_in_r_bypass_23_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_0_df_is_ws_16 <= io_in_r_bypass_23_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_0_stall_16 <= io_in_r_bypass_23_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_1_data_16 <= io_in_r_bypass_23_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_1_load_store_16 <= io_in_r_bypass_23_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_1_df_is_ws_16 <= io_in_r_bypass_23_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_1_stall_16 <= io_in_r_bypass_23_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_2_data_16 <= io_in_r_bypass_23_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_2_load_store_16 <= io_in_r_bypass_23_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_2_df_is_ws_16 <= io_in_r_bypass_23_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_2_stall_16 <= io_in_r_bypass_23_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_3_data_16 <= io_in_r_bypass_23_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_3_load_store_16 <= io_in_r_bypass_23_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_3_df_is_ws_16 <= io_in_r_bypass_23_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_3_stall_16 <= io_in_r_bypass_23_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_0_data_16 <= io_in_r_bypass_24_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_0_load_store_16 <= io_in_r_bypass_24_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_0_df_is_ws_16 <= io_in_r_bypass_24_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_0_stall_16 <= io_in_r_bypass_24_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_1_data_16 <= io_in_r_bypass_24_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_1_load_store_16 <= io_in_r_bypass_24_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_1_df_is_ws_16 <= io_in_r_bypass_24_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_1_stall_16 <= io_in_r_bypass_24_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_2_data_16 <= io_in_r_bypass_24_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_2_load_store_16 <= io_in_r_bypass_24_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_2_df_is_ws_16 <= io_in_r_bypass_24_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_2_stall_16 <= io_in_r_bypass_24_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_3_data_16 <= io_in_r_bypass_24_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_3_load_store_16 <= io_in_r_bypass_24_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_3_df_is_ws_16 <= io_in_r_bypass_24_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_3_stall_16 <= io_in_r_bypass_24_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_0_data_16 <= io_in_r_bypass_25_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_0_load_store_16 <= io_in_r_bypass_25_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_0_df_is_ws_16 <= io_in_r_bypass_25_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_0_stall_16 <= io_in_r_bypass_25_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_1_data_16 <= io_in_r_bypass_25_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_1_load_store_16 <= io_in_r_bypass_25_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_1_df_is_ws_16 <= io_in_r_bypass_25_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_1_stall_16 <= io_in_r_bypass_25_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_2_data_16 <= io_in_r_bypass_25_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_2_load_store_16 <= io_in_r_bypass_25_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_2_df_is_ws_16 <= io_in_r_bypass_25_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_2_stall_16 <= io_in_r_bypass_25_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_3_data_16 <= io_in_r_bypass_25_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_3_load_store_16 <= io_in_r_bypass_25_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_3_df_is_ws_16 <= io_in_r_bypass_25_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_3_stall_16 <= io_in_r_bypass_25_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_0_data_16 <= io_in_r_bypass_26_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_0_load_store_16 <= io_in_r_bypass_26_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_0_df_is_ws_16 <= io_in_r_bypass_26_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_0_stall_16 <= io_in_r_bypass_26_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_1_data_16 <= io_in_r_bypass_26_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_1_load_store_16 <= io_in_r_bypass_26_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_1_df_is_ws_16 <= io_in_r_bypass_26_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_1_stall_16 <= io_in_r_bypass_26_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_2_data_16 <= io_in_r_bypass_26_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_2_load_store_16 <= io_in_r_bypass_26_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_2_df_is_ws_16 <= io_in_r_bypass_26_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_2_stall_16 <= io_in_r_bypass_26_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_3_data_16 <= io_in_r_bypass_26_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_3_load_store_16 <= io_in_r_bypass_26_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_3_df_is_ws_16 <= io_in_r_bypass_26_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_3_stall_16 <= io_in_r_bypass_26_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_0_data_16 <= io_in_r_bypass_27_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_0_load_store_16 <= io_in_r_bypass_27_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_0_df_is_ws_16 <= io_in_r_bypass_27_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_0_stall_16 <= io_in_r_bypass_27_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_1_data_16 <= io_in_r_bypass_27_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_1_load_store_16 <= io_in_r_bypass_27_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_1_df_is_ws_16 <= io_in_r_bypass_27_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_1_stall_16 <= io_in_r_bypass_27_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_2_data_16 <= io_in_r_bypass_27_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_2_load_store_16 <= io_in_r_bypass_27_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_2_df_is_ws_16 <= io_in_r_bypass_27_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_2_stall_16 <= io_in_r_bypass_27_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_3_data_16 <= io_in_r_bypass_27_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_3_load_store_16 <= io_in_r_bypass_27_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_3_df_is_ws_16 <= io_in_r_bypass_27_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_3_stall_16 <= io_in_r_bypass_27_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_0_data_16 <= io_in_r_bypass_28_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_0_load_store_16 <= io_in_r_bypass_28_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_0_df_is_ws_16 <= io_in_r_bypass_28_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_0_stall_16 <= io_in_r_bypass_28_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_1_data_16 <= io_in_r_bypass_28_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_1_load_store_16 <= io_in_r_bypass_28_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_1_df_is_ws_16 <= io_in_r_bypass_28_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_1_stall_16 <= io_in_r_bypass_28_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_2_data_16 <= io_in_r_bypass_28_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_2_load_store_16 <= io_in_r_bypass_28_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_2_df_is_ws_16 <= io_in_r_bypass_28_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_2_stall_16 <= io_in_r_bypass_28_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_3_data_16 <= io_in_r_bypass_28_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_3_load_store_16 <= io_in_r_bypass_28_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_3_df_is_ws_16 <= io_in_r_bypass_28_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_3_stall_16 <= io_in_r_bypass_28_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_0_data_16 <= io_in_r_bypass_29_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_0_load_store_16 <= io_in_r_bypass_29_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_0_df_is_ws_16 <= io_in_r_bypass_29_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_0_stall_16 <= io_in_r_bypass_29_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_1_data_16 <= io_in_r_bypass_29_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_1_load_store_16 <= io_in_r_bypass_29_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_1_df_is_ws_16 <= io_in_r_bypass_29_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_1_stall_16 <= io_in_r_bypass_29_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_2_data_16 <= io_in_r_bypass_29_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_2_load_store_16 <= io_in_r_bypass_29_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_2_df_is_ws_16 <= io_in_r_bypass_29_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_2_stall_16 <= io_in_r_bypass_29_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_3_data_16 <= io_in_r_bypass_29_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_3_load_store_16 <= io_in_r_bypass_29_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_3_df_is_ws_16 <= io_in_r_bypass_29_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_3_stall_16 <= io_in_r_bypass_29_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_0_data_16 <= io_in_r_bypass_30_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_0_load_store_16 <= io_in_r_bypass_30_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_0_df_is_ws_16 <= io_in_r_bypass_30_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_0_stall_16 <= io_in_r_bypass_30_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_1_data_16 <= io_in_r_bypass_30_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_1_load_store_16 <= io_in_r_bypass_30_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_1_df_is_ws_16 <= io_in_r_bypass_30_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_1_stall_16 <= io_in_r_bypass_30_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_2_data_16 <= io_in_r_bypass_30_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_2_load_store_16 <= io_in_r_bypass_30_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_2_df_is_ws_16 <= io_in_r_bypass_30_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_2_stall_16 <= io_in_r_bypass_30_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_3_data_16 <= io_in_r_bypass_30_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_3_load_store_16 <= io_in_r_bypass_30_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_3_df_is_ws_16 <= io_in_r_bypass_30_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_3_stall_16 <= io_in_r_bypass_30_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_0_data_16 <= io_in_r_bypass_31_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_0_load_store_16 <= io_in_r_bypass_31_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_0_df_is_ws_16 <= io_in_r_bypass_31_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_0_stall_16 <= io_in_r_bypass_31_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_1_data_16 <= io_in_r_bypass_31_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_1_load_store_16 <= io_in_r_bypass_31_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_1_df_is_ws_16 <= io_in_r_bypass_31_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_1_stall_16 <= io_in_r_bypass_31_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_2_data_16 <= io_in_r_bypass_31_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_2_load_store_16 <= io_in_r_bypass_31_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_2_df_is_ws_16 <= io_in_r_bypass_31_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_2_stall_16 <= io_in_r_bypass_31_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_3_data_16 <= io_in_r_bypass_31_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_3_load_store_16 <= io_in_r_bypass_31_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_3_df_is_ws_16 <= io_in_r_bypass_31_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_3_stall_16 <= io_in_r_bypass_31_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_0_data_17 <= io_in_r_bypass_0_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_0_load_store_17 <= io_in_r_bypass_0_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_0_df_is_ws_17 <= io_in_r_bypass_0_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_0_stall_17 <= io_in_r_bypass_0_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_1_data_17 <= io_in_r_bypass_0_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_1_load_store_17 <= io_in_r_bypass_0_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_1_df_is_ws_17 <= io_in_r_bypass_0_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_1_stall_17 <= io_in_r_bypass_0_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_2_data_17 <= io_in_r_bypass_0_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_2_load_store_17 <= io_in_r_bypass_0_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_2_df_is_ws_17 <= io_in_r_bypass_0_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_2_stall_17 <= io_in_r_bypass_0_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_3_data_17 <= io_in_r_bypass_0_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_3_load_store_17 <= io_in_r_bypass_0_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_3_df_is_ws_17 <= io_in_r_bypass_0_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_3_stall_17 <= io_in_r_bypass_0_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_0_data_17 <= io_in_r_bypass_1_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_0_load_store_17 <= io_in_r_bypass_1_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_0_df_is_ws_17 <= io_in_r_bypass_1_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_0_stall_17 <= io_in_r_bypass_1_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_1_data_17 <= io_in_r_bypass_1_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_1_load_store_17 <= io_in_r_bypass_1_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_1_df_is_ws_17 <= io_in_r_bypass_1_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_1_stall_17 <= io_in_r_bypass_1_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_2_data_17 <= io_in_r_bypass_1_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_2_load_store_17 <= io_in_r_bypass_1_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_2_df_is_ws_17 <= io_in_r_bypass_1_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_2_stall_17 <= io_in_r_bypass_1_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_3_data_17 <= io_in_r_bypass_1_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_3_load_store_17 <= io_in_r_bypass_1_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_3_df_is_ws_17 <= io_in_r_bypass_1_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_3_stall_17 <= io_in_r_bypass_1_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_0_data_17 <= io_in_r_bypass_2_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_0_load_store_17 <= io_in_r_bypass_2_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_0_df_is_ws_17 <= io_in_r_bypass_2_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_0_stall_17 <= io_in_r_bypass_2_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_1_data_17 <= io_in_r_bypass_2_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_1_load_store_17 <= io_in_r_bypass_2_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_1_df_is_ws_17 <= io_in_r_bypass_2_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_1_stall_17 <= io_in_r_bypass_2_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_2_data_17 <= io_in_r_bypass_2_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_2_load_store_17 <= io_in_r_bypass_2_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_2_df_is_ws_17 <= io_in_r_bypass_2_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_2_stall_17 <= io_in_r_bypass_2_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_3_data_17 <= io_in_r_bypass_2_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_3_load_store_17 <= io_in_r_bypass_2_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_3_df_is_ws_17 <= io_in_r_bypass_2_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_3_stall_17 <= io_in_r_bypass_2_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_0_data_17 <= io_in_r_bypass_3_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_0_load_store_17 <= io_in_r_bypass_3_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_0_df_is_ws_17 <= io_in_r_bypass_3_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_0_stall_17 <= io_in_r_bypass_3_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_1_data_17 <= io_in_r_bypass_3_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_1_load_store_17 <= io_in_r_bypass_3_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_1_df_is_ws_17 <= io_in_r_bypass_3_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_1_stall_17 <= io_in_r_bypass_3_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_2_data_17 <= io_in_r_bypass_3_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_2_load_store_17 <= io_in_r_bypass_3_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_2_df_is_ws_17 <= io_in_r_bypass_3_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_2_stall_17 <= io_in_r_bypass_3_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_3_data_17 <= io_in_r_bypass_3_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_3_load_store_17 <= io_in_r_bypass_3_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_3_df_is_ws_17 <= io_in_r_bypass_3_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_3_stall_17 <= io_in_r_bypass_3_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_0_data_17 <= io_in_r_bypass_4_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_0_load_store_17 <= io_in_r_bypass_4_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_0_df_is_ws_17 <= io_in_r_bypass_4_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_0_stall_17 <= io_in_r_bypass_4_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_1_data_17 <= io_in_r_bypass_4_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_1_load_store_17 <= io_in_r_bypass_4_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_1_df_is_ws_17 <= io_in_r_bypass_4_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_1_stall_17 <= io_in_r_bypass_4_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_2_data_17 <= io_in_r_bypass_4_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_2_load_store_17 <= io_in_r_bypass_4_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_2_df_is_ws_17 <= io_in_r_bypass_4_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_2_stall_17 <= io_in_r_bypass_4_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_3_data_17 <= io_in_r_bypass_4_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_3_load_store_17 <= io_in_r_bypass_4_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_3_df_is_ws_17 <= io_in_r_bypass_4_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_3_stall_17 <= io_in_r_bypass_4_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_0_data_17 <= io_in_r_bypass_5_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_0_load_store_17 <= io_in_r_bypass_5_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_0_df_is_ws_17 <= io_in_r_bypass_5_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_0_stall_17 <= io_in_r_bypass_5_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_1_data_17 <= io_in_r_bypass_5_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_1_load_store_17 <= io_in_r_bypass_5_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_1_df_is_ws_17 <= io_in_r_bypass_5_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_1_stall_17 <= io_in_r_bypass_5_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_2_data_17 <= io_in_r_bypass_5_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_2_load_store_17 <= io_in_r_bypass_5_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_2_df_is_ws_17 <= io_in_r_bypass_5_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_2_stall_17 <= io_in_r_bypass_5_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_3_data_17 <= io_in_r_bypass_5_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_3_load_store_17 <= io_in_r_bypass_5_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_3_df_is_ws_17 <= io_in_r_bypass_5_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_3_stall_17 <= io_in_r_bypass_5_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_0_data_17 <= io_in_r_bypass_6_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_0_load_store_17 <= io_in_r_bypass_6_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_0_df_is_ws_17 <= io_in_r_bypass_6_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_0_stall_17 <= io_in_r_bypass_6_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_1_data_17 <= io_in_r_bypass_6_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_1_load_store_17 <= io_in_r_bypass_6_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_1_df_is_ws_17 <= io_in_r_bypass_6_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_1_stall_17 <= io_in_r_bypass_6_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_2_data_17 <= io_in_r_bypass_6_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_2_load_store_17 <= io_in_r_bypass_6_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_2_df_is_ws_17 <= io_in_r_bypass_6_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_2_stall_17 <= io_in_r_bypass_6_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_3_data_17 <= io_in_r_bypass_6_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_3_load_store_17 <= io_in_r_bypass_6_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_3_df_is_ws_17 <= io_in_r_bypass_6_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_3_stall_17 <= io_in_r_bypass_6_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_0_data_17 <= io_in_r_bypass_7_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_0_load_store_17 <= io_in_r_bypass_7_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_0_df_is_ws_17 <= io_in_r_bypass_7_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_0_stall_17 <= io_in_r_bypass_7_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_1_data_17 <= io_in_r_bypass_7_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_1_load_store_17 <= io_in_r_bypass_7_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_1_df_is_ws_17 <= io_in_r_bypass_7_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_1_stall_17 <= io_in_r_bypass_7_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_2_data_17 <= io_in_r_bypass_7_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_2_load_store_17 <= io_in_r_bypass_7_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_2_df_is_ws_17 <= io_in_r_bypass_7_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_2_stall_17 <= io_in_r_bypass_7_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_3_data_17 <= io_in_r_bypass_7_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_3_load_store_17 <= io_in_r_bypass_7_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_3_df_is_ws_17 <= io_in_r_bypass_7_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_3_stall_17 <= io_in_r_bypass_7_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_0_data_17 <= io_in_r_bypass_8_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_0_load_store_17 <= io_in_r_bypass_8_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_0_df_is_ws_17 <= io_in_r_bypass_8_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_0_stall_17 <= io_in_r_bypass_8_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_1_data_17 <= io_in_r_bypass_8_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_1_load_store_17 <= io_in_r_bypass_8_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_1_df_is_ws_17 <= io_in_r_bypass_8_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_1_stall_17 <= io_in_r_bypass_8_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_2_data_17 <= io_in_r_bypass_8_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_2_load_store_17 <= io_in_r_bypass_8_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_2_df_is_ws_17 <= io_in_r_bypass_8_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_2_stall_17 <= io_in_r_bypass_8_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_3_data_17 <= io_in_r_bypass_8_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_3_load_store_17 <= io_in_r_bypass_8_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_3_df_is_ws_17 <= io_in_r_bypass_8_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_3_stall_17 <= io_in_r_bypass_8_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_0_data_17 <= io_in_r_bypass_9_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_0_load_store_17 <= io_in_r_bypass_9_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_0_df_is_ws_17 <= io_in_r_bypass_9_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_0_stall_17 <= io_in_r_bypass_9_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_1_data_17 <= io_in_r_bypass_9_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_1_load_store_17 <= io_in_r_bypass_9_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_1_df_is_ws_17 <= io_in_r_bypass_9_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_1_stall_17 <= io_in_r_bypass_9_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_2_data_17 <= io_in_r_bypass_9_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_2_load_store_17 <= io_in_r_bypass_9_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_2_df_is_ws_17 <= io_in_r_bypass_9_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_2_stall_17 <= io_in_r_bypass_9_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_3_data_17 <= io_in_r_bypass_9_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_3_load_store_17 <= io_in_r_bypass_9_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_3_df_is_ws_17 <= io_in_r_bypass_9_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_3_stall_17 <= io_in_r_bypass_9_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_0_data_17 <= io_in_r_bypass_10_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_0_load_store_17 <= io_in_r_bypass_10_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_0_df_is_ws_17 <= io_in_r_bypass_10_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_0_stall_17 <= io_in_r_bypass_10_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_1_data_17 <= io_in_r_bypass_10_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_1_load_store_17 <= io_in_r_bypass_10_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_1_df_is_ws_17 <= io_in_r_bypass_10_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_1_stall_17 <= io_in_r_bypass_10_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_2_data_17 <= io_in_r_bypass_10_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_2_load_store_17 <= io_in_r_bypass_10_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_2_df_is_ws_17 <= io_in_r_bypass_10_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_2_stall_17 <= io_in_r_bypass_10_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_3_data_17 <= io_in_r_bypass_10_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_3_load_store_17 <= io_in_r_bypass_10_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_3_df_is_ws_17 <= io_in_r_bypass_10_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_3_stall_17 <= io_in_r_bypass_10_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_0_data_17 <= io_in_r_bypass_11_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_0_load_store_17 <= io_in_r_bypass_11_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_0_df_is_ws_17 <= io_in_r_bypass_11_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_0_stall_17 <= io_in_r_bypass_11_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_1_data_17 <= io_in_r_bypass_11_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_1_load_store_17 <= io_in_r_bypass_11_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_1_df_is_ws_17 <= io_in_r_bypass_11_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_1_stall_17 <= io_in_r_bypass_11_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_2_data_17 <= io_in_r_bypass_11_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_2_load_store_17 <= io_in_r_bypass_11_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_2_df_is_ws_17 <= io_in_r_bypass_11_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_2_stall_17 <= io_in_r_bypass_11_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_3_data_17 <= io_in_r_bypass_11_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_3_load_store_17 <= io_in_r_bypass_11_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_3_df_is_ws_17 <= io_in_r_bypass_11_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_3_stall_17 <= io_in_r_bypass_11_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_0_data_17 <= io_in_r_bypass_12_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_0_load_store_17 <= io_in_r_bypass_12_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_0_df_is_ws_17 <= io_in_r_bypass_12_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_0_stall_17 <= io_in_r_bypass_12_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_1_data_17 <= io_in_r_bypass_12_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_1_load_store_17 <= io_in_r_bypass_12_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_1_df_is_ws_17 <= io_in_r_bypass_12_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_1_stall_17 <= io_in_r_bypass_12_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_2_data_17 <= io_in_r_bypass_12_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_2_load_store_17 <= io_in_r_bypass_12_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_2_df_is_ws_17 <= io_in_r_bypass_12_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_2_stall_17 <= io_in_r_bypass_12_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_3_data_17 <= io_in_r_bypass_12_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_3_load_store_17 <= io_in_r_bypass_12_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_3_df_is_ws_17 <= io_in_r_bypass_12_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_3_stall_17 <= io_in_r_bypass_12_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_0_data_17 <= io_in_r_bypass_13_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_0_load_store_17 <= io_in_r_bypass_13_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_0_df_is_ws_17 <= io_in_r_bypass_13_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_0_stall_17 <= io_in_r_bypass_13_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_1_data_17 <= io_in_r_bypass_13_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_1_load_store_17 <= io_in_r_bypass_13_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_1_df_is_ws_17 <= io_in_r_bypass_13_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_1_stall_17 <= io_in_r_bypass_13_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_2_data_17 <= io_in_r_bypass_13_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_2_load_store_17 <= io_in_r_bypass_13_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_2_df_is_ws_17 <= io_in_r_bypass_13_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_2_stall_17 <= io_in_r_bypass_13_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_3_data_17 <= io_in_r_bypass_13_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_3_load_store_17 <= io_in_r_bypass_13_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_3_df_is_ws_17 <= io_in_r_bypass_13_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_3_stall_17 <= io_in_r_bypass_13_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_0_data_17 <= io_in_r_bypass_14_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_0_load_store_17 <= io_in_r_bypass_14_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_0_df_is_ws_17 <= io_in_r_bypass_14_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_0_stall_17 <= io_in_r_bypass_14_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_1_data_17 <= io_in_r_bypass_14_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_1_load_store_17 <= io_in_r_bypass_14_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_1_df_is_ws_17 <= io_in_r_bypass_14_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_1_stall_17 <= io_in_r_bypass_14_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_2_data_17 <= io_in_r_bypass_14_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_2_load_store_17 <= io_in_r_bypass_14_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_2_df_is_ws_17 <= io_in_r_bypass_14_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_2_stall_17 <= io_in_r_bypass_14_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_3_data_17 <= io_in_r_bypass_14_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_3_load_store_17 <= io_in_r_bypass_14_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_3_df_is_ws_17 <= io_in_r_bypass_14_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_3_stall_17 <= io_in_r_bypass_14_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_0_data_17 <= io_in_r_bypass_15_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_0_load_store_17 <= io_in_r_bypass_15_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_0_df_is_ws_17 <= io_in_r_bypass_15_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_0_stall_17 <= io_in_r_bypass_15_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_1_data_17 <= io_in_r_bypass_15_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_1_load_store_17 <= io_in_r_bypass_15_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_1_df_is_ws_17 <= io_in_r_bypass_15_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_1_stall_17 <= io_in_r_bypass_15_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_2_data_17 <= io_in_r_bypass_15_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_2_load_store_17 <= io_in_r_bypass_15_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_2_df_is_ws_17 <= io_in_r_bypass_15_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_2_stall_17 <= io_in_r_bypass_15_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_3_data_17 <= io_in_r_bypass_15_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_3_load_store_17 <= io_in_r_bypass_15_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_3_df_is_ws_17 <= io_in_r_bypass_15_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_3_stall_17 <= io_in_r_bypass_15_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_0_data_17 <= io_in_r_bypass_16_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_0_load_store_17 <= io_in_r_bypass_16_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_0_df_is_ws_17 <= io_in_r_bypass_16_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_0_stall_17 <= io_in_r_bypass_16_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_1_data_17 <= io_in_r_bypass_16_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_1_load_store_17 <= io_in_r_bypass_16_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_1_df_is_ws_17 <= io_in_r_bypass_16_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_1_stall_17 <= io_in_r_bypass_16_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_2_data_17 <= io_in_r_bypass_16_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_2_load_store_17 <= io_in_r_bypass_16_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_2_df_is_ws_17 <= io_in_r_bypass_16_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_2_stall_17 <= io_in_r_bypass_16_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_3_data_17 <= io_in_r_bypass_16_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_3_load_store_17 <= io_in_r_bypass_16_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_3_df_is_ws_17 <= io_in_r_bypass_16_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_3_stall_17 <= io_in_r_bypass_16_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_0_data_17 <= io_in_r_bypass_17_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_0_load_store_17 <= io_in_r_bypass_17_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_0_df_is_ws_17 <= io_in_r_bypass_17_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_0_stall_17 <= io_in_r_bypass_17_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_1_data_17 <= io_in_r_bypass_17_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_1_load_store_17 <= io_in_r_bypass_17_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_1_df_is_ws_17 <= io_in_r_bypass_17_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_1_stall_17 <= io_in_r_bypass_17_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_2_data_17 <= io_in_r_bypass_17_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_2_load_store_17 <= io_in_r_bypass_17_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_2_df_is_ws_17 <= io_in_r_bypass_17_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_2_stall_17 <= io_in_r_bypass_17_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_3_data_17 <= io_in_r_bypass_17_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_3_load_store_17 <= io_in_r_bypass_17_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_3_df_is_ws_17 <= io_in_r_bypass_17_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_3_stall_17 <= io_in_r_bypass_17_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_0_data_17 <= io_in_r_bypass_18_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_0_load_store_17 <= io_in_r_bypass_18_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_0_df_is_ws_17 <= io_in_r_bypass_18_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_0_stall_17 <= io_in_r_bypass_18_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_1_data_17 <= io_in_r_bypass_18_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_1_load_store_17 <= io_in_r_bypass_18_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_1_df_is_ws_17 <= io_in_r_bypass_18_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_1_stall_17 <= io_in_r_bypass_18_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_2_data_17 <= io_in_r_bypass_18_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_2_load_store_17 <= io_in_r_bypass_18_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_2_df_is_ws_17 <= io_in_r_bypass_18_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_2_stall_17 <= io_in_r_bypass_18_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_3_data_17 <= io_in_r_bypass_18_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_3_load_store_17 <= io_in_r_bypass_18_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_3_df_is_ws_17 <= io_in_r_bypass_18_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_3_stall_17 <= io_in_r_bypass_18_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_0_data_17 <= io_in_r_bypass_19_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_0_load_store_17 <= io_in_r_bypass_19_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_0_df_is_ws_17 <= io_in_r_bypass_19_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_0_stall_17 <= io_in_r_bypass_19_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_1_data_17 <= io_in_r_bypass_19_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_1_load_store_17 <= io_in_r_bypass_19_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_1_df_is_ws_17 <= io_in_r_bypass_19_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_1_stall_17 <= io_in_r_bypass_19_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_2_data_17 <= io_in_r_bypass_19_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_2_load_store_17 <= io_in_r_bypass_19_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_2_df_is_ws_17 <= io_in_r_bypass_19_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_2_stall_17 <= io_in_r_bypass_19_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_3_data_17 <= io_in_r_bypass_19_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_3_load_store_17 <= io_in_r_bypass_19_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_3_df_is_ws_17 <= io_in_r_bypass_19_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_3_stall_17 <= io_in_r_bypass_19_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_0_data_17 <= io_in_r_bypass_20_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_0_load_store_17 <= io_in_r_bypass_20_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_0_df_is_ws_17 <= io_in_r_bypass_20_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_0_stall_17 <= io_in_r_bypass_20_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_1_data_17 <= io_in_r_bypass_20_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_1_load_store_17 <= io_in_r_bypass_20_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_1_df_is_ws_17 <= io_in_r_bypass_20_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_1_stall_17 <= io_in_r_bypass_20_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_2_data_17 <= io_in_r_bypass_20_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_2_load_store_17 <= io_in_r_bypass_20_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_2_df_is_ws_17 <= io_in_r_bypass_20_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_2_stall_17 <= io_in_r_bypass_20_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_3_data_17 <= io_in_r_bypass_20_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_3_load_store_17 <= io_in_r_bypass_20_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_3_df_is_ws_17 <= io_in_r_bypass_20_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_3_stall_17 <= io_in_r_bypass_20_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_0_data_17 <= io_in_r_bypass_21_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_0_load_store_17 <= io_in_r_bypass_21_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_0_df_is_ws_17 <= io_in_r_bypass_21_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_0_stall_17 <= io_in_r_bypass_21_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_1_data_17 <= io_in_r_bypass_21_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_1_load_store_17 <= io_in_r_bypass_21_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_1_df_is_ws_17 <= io_in_r_bypass_21_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_1_stall_17 <= io_in_r_bypass_21_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_2_data_17 <= io_in_r_bypass_21_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_2_load_store_17 <= io_in_r_bypass_21_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_2_df_is_ws_17 <= io_in_r_bypass_21_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_2_stall_17 <= io_in_r_bypass_21_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_3_data_17 <= io_in_r_bypass_21_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_3_load_store_17 <= io_in_r_bypass_21_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_3_df_is_ws_17 <= io_in_r_bypass_21_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_3_stall_17 <= io_in_r_bypass_21_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_0_data_17 <= io_in_r_bypass_22_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_0_load_store_17 <= io_in_r_bypass_22_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_0_df_is_ws_17 <= io_in_r_bypass_22_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_0_stall_17 <= io_in_r_bypass_22_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_1_data_17 <= io_in_r_bypass_22_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_1_load_store_17 <= io_in_r_bypass_22_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_1_df_is_ws_17 <= io_in_r_bypass_22_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_1_stall_17 <= io_in_r_bypass_22_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_2_data_17 <= io_in_r_bypass_22_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_2_load_store_17 <= io_in_r_bypass_22_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_2_df_is_ws_17 <= io_in_r_bypass_22_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_2_stall_17 <= io_in_r_bypass_22_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_3_data_17 <= io_in_r_bypass_22_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_3_load_store_17 <= io_in_r_bypass_22_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_3_df_is_ws_17 <= io_in_r_bypass_22_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_3_stall_17 <= io_in_r_bypass_22_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_0_data_17 <= io_in_r_bypass_23_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_0_load_store_17 <= io_in_r_bypass_23_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_0_df_is_ws_17 <= io_in_r_bypass_23_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_0_stall_17 <= io_in_r_bypass_23_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_1_data_17 <= io_in_r_bypass_23_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_1_load_store_17 <= io_in_r_bypass_23_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_1_df_is_ws_17 <= io_in_r_bypass_23_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_1_stall_17 <= io_in_r_bypass_23_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_2_data_17 <= io_in_r_bypass_23_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_2_load_store_17 <= io_in_r_bypass_23_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_2_df_is_ws_17 <= io_in_r_bypass_23_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_2_stall_17 <= io_in_r_bypass_23_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_3_data_17 <= io_in_r_bypass_23_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_3_load_store_17 <= io_in_r_bypass_23_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_3_df_is_ws_17 <= io_in_r_bypass_23_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_3_stall_17 <= io_in_r_bypass_23_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_0_data_17 <= io_in_r_bypass_24_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_0_load_store_17 <= io_in_r_bypass_24_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_0_df_is_ws_17 <= io_in_r_bypass_24_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_0_stall_17 <= io_in_r_bypass_24_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_1_data_17 <= io_in_r_bypass_24_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_1_load_store_17 <= io_in_r_bypass_24_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_1_df_is_ws_17 <= io_in_r_bypass_24_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_1_stall_17 <= io_in_r_bypass_24_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_2_data_17 <= io_in_r_bypass_24_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_2_load_store_17 <= io_in_r_bypass_24_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_2_df_is_ws_17 <= io_in_r_bypass_24_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_2_stall_17 <= io_in_r_bypass_24_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_3_data_17 <= io_in_r_bypass_24_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_3_load_store_17 <= io_in_r_bypass_24_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_3_df_is_ws_17 <= io_in_r_bypass_24_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_3_stall_17 <= io_in_r_bypass_24_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_0_data_17 <= io_in_r_bypass_25_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_0_load_store_17 <= io_in_r_bypass_25_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_0_df_is_ws_17 <= io_in_r_bypass_25_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_0_stall_17 <= io_in_r_bypass_25_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_1_data_17 <= io_in_r_bypass_25_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_1_load_store_17 <= io_in_r_bypass_25_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_1_df_is_ws_17 <= io_in_r_bypass_25_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_1_stall_17 <= io_in_r_bypass_25_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_2_data_17 <= io_in_r_bypass_25_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_2_load_store_17 <= io_in_r_bypass_25_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_2_df_is_ws_17 <= io_in_r_bypass_25_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_2_stall_17 <= io_in_r_bypass_25_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_3_data_17 <= io_in_r_bypass_25_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_3_load_store_17 <= io_in_r_bypass_25_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_3_df_is_ws_17 <= io_in_r_bypass_25_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_3_stall_17 <= io_in_r_bypass_25_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_0_data_17 <= io_in_r_bypass_26_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_0_load_store_17 <= io_in_r_bypass_26_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_0_df_is_ws_17 <= io_in_r_bypass_26_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_0_stall_17 <= io_in_r_bypass_26_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_1_data_17 <= io_in_r_bypass_26_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_1_load_store_17 <= io_in_r_bypass_26_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_1_df_is_ws_17 <= io_in_r_bypass_26_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_1_stall_17 <= io_in_r_bypass_26_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_2_data_17 <= io_in_r_bypass_26_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_2_load_store_17 <= io_in_r_bypass_26_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_2_df_is_ws_17 <= io_in_r_bypass_26_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_2_stall_17 <= io_in_r_bypass_26_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_3_data_17 <= io_in_r_bypass_26_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_3_load_store_17 <= io_in_r_bypass_26_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_3_df_is_ws_17 <= io_in_r_bypass_26_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_3_stall_17 <= io_in_r_bypass_26_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_0_data_17 <= io_in_r_bypass_27_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_0_load_store_17 <= io_in_r_bypass_27_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_0_df_is_ws_17 <= io_in_r_bypass_27_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_0_stall_17 <= io_in_r_bypass_27_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_1_data_17 <= io_in_r_bypass_27_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_1_load_store_17 <= io_in_r_bypass_27_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_1_df_is_ws_17 <= io_in_r_bypass_27_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_1_stall_17 <= io_in_r_bypass_27_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_2_data_17 <= io_in_r_bypass_27_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_2_load_store_17 <= io_in_r_bypass_27_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_2_df_is_ws_17 <= io_in_r_bypass_27_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_2_stall_17 <= io_in_r_bypass_27_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_3_data_17 <= io_in_r_bypass_27_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_3_load_store_17 <= io_in_r_bypass_27_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_3_df_is_ws_17 <= io_in_r_bypass_27_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_3_stall_17 <= io_in_r_bypass_27_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_0_data_17 <= io_in_r_bypass_28_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_0_load_store_17 <= io_in_r_bypass_28_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_0_df_is_ws_17 <= io_in_r_bypass_28_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_0_stall_17 <= io_in_r_bypass_28_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_1_data_17 <= io_in_r_bypass_28_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_1_load_store_17 <= io_in_r_bypass_28_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_1_df_is_ws_17 <= io_in_r_bypass_28_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_1_stall_17 <= io_in_r_bypass_28_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_2_data_17 <= io_in_r_bypass_28_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_2_load_store_17 <= io_in_r_bypass_28_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_2_df_is_ws_17 <= io_in_r_bypass_28_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_2_stall_17 <= io_in_r_bypass_28_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_3_data_17 <= io_in_r_bypass_28_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_3_load_store_17 <= io_in_r_bypass_28_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_3_df_is_ws_17 <= io_in_r_bypass_28_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_3_stall_17 <= io_in_r_bypass_28_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_0_data_17 <= io_in_r_bypass_29_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_0_load_store_17 <= io_in_r_bypass_29_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_0_df_is_ws_17 <= io_in_r_bypass_29_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_0_stall_17 <= io_in_r_bypass_29_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_1_data_17 <= io_in_r_bypass_29_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_1_load_store_17 <= io_in_r_bypass_29_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_1_df_is_ws_17 <= io_in_r_bypass_29_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_1_stall_17 <= io_in_r_bypass_29_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_2_data_17 <= io_in_r_bypass_29_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_2_load_store_17 <= io_in_r_bypass_29_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_2_df_is_ws_17 <= io_in_r_bypass_29_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_2_stall_17 <= io_in_r_bypass_29_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_3_data_17 <= io_in_r_bypass_29_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_3_load_store_17 <= io_in_r_bypass_29_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_3_df_is_ws_17 <= io_in_r_bypass_29_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_3_stall_17 <= io_in_r_bypass_29_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_0_data_17 <= io_in_r_bypass_30_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_0_load_store_17 <= io_in_r_bypass_30_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_0_df_is_ws_17 <= io_in_r_bypass_30_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_0_stall_17 <= io_in_r_bypass_30_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_1_data_17 <= io_in_r_bypass_30_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_1_load_store_17 <= io_in_r_bypass_30_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_1_df_is_ws_17 <= io_in_r_bypass_30_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_1_stall_17 <= io_in_r_bypass_30_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_2_data_17 <= io_in_r_bypass_30_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_2_load_store_17 <= io_in_r_bypass_30_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_2_df_is_ws_17 <= io_in_r_bypass_30_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_2_stall_17 <= io_in_r_bypass_30_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_3_data_17 <= io_in_r_bypass_30_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_3_load_store_17 <= io_in_r_bypass_30_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_3_df_is_ws_17 <= io_in_r_bypass_30_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_3_stall_17 <= io_in_r_bypass_30_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_0_data_17 <= io_in_r_bypass_31_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_0_load_store_17 <= io_in_r_bypass_31_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_0_df_is_ws_17 <= io_in_r_bypass_31_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_0_stall_17 <= io_in_r_bypass_31_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_1_data_17 <= io_in_r_bypass_31_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_1_load_store_17 <= io_in_r_bypass_31_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_1_df_is_ws_17 <= io_in_r_bypass_31_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_1_stall_17 <= io_in_r_bypass_31_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_2_data_17 <= io_in_r_bypass_31_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_2_load_store_17 <= io_in_r_bypass_31_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_2_df_is_ws_17 <= io_in_r_bypass_31_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_2_stall_17 <= io_in_r_bypass_31_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_3_data_17 <= io_in_r_bypass_31_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_3_load_store_17 <= io_in_r_bypass_31_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_3_df_is_ws_17 <= io_in_r_bypass_31_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_3_stall_17 <= io_in_r_bypass_31_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_0_data_18 <= io_in_r_bypass_0_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_0_load_store_18 <= io_in_r_bypass_0_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_0_df_is_ws_18 <= io_in_r_bypass_0_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_0_stall_18 <= io_in_r_bypass_0_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_1_data_18 <= io_in_r_bypass_0_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_1_load_store_18 <= io_in_r_bypass_0_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_1_df_is_ws_18 <= io_in_r_bypass_0_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_1_stall_18 <= io_in_r_bypass_0_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_2_data_18 <= io_in_r_bypass_0_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_2_load_store_18 <= io_in_r_bypass_0_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_2_df_is_ws_18 <= io_in_r_bypass_0_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_2_stall_18 <= io_in_r_bypass_0_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_3_data_18 <= io_in_r_bypass_0_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_3_load_store_18 <= io_in_r_bypass_0_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_3_df_is_ws_18 <= io_in_r_bypass_0_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_3_stall_18 <= io_in_r_bypass_0_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_0_data_18 <= io_in_r_bypass_1_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_0_load_store_18 <= io_in_r_bypass_1_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_0_df_is_ws_18 <= io_in_r_bypass_1_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_0_stall_18 <= io_in_r_bypass_1_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_1_data_18 <= io_in_r_bypass_1_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_1_load_store_18 <= io_in_r_bypass_1_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_1_df_is_ws_18 <= io_in_r_bypass_1_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_1_stall_18 <= io_in_r_bypass_1_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_2_data_18 <= io_in_r_bypass_1_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_2_load_store_18 <= io_in_r_bypass_1_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_2_df_is_ws_18 <= io_in_r_bypass_1_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_2_stall_18 <= io_in_r_bypass_1_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_3_data_18 <= io_in_r_bypass_1_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_3_load_store_18 <= io_in_r_bypass_1_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_3_df_is_ws_18 <= io_in_r_bypass_1_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_3_stall_18 <= io_in_r_bypass_1_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_0_data_18 <= io_in_r_bypass_2_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_0_load_store_18 <= io_in_r_bypass_2_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_0_df_is_ws_18 <= io_in_r_bypass_2_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_0_stall_18 <= io_in_r_bypass_2_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_1_data_18 <= io_in_r_bypass_2_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_1_load_store_18 <= io_in_r_bypass_2_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_1_df_is_ws_18 <= io_in_r_bypass_2_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_1_stall_18 <= io_in_r_bypass_2_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_2_data_18 <= io_in_r_bypass_2_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_2_load_store_18 <= io_in_r_bypass_2_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_2_df_is_ws_18 <= io_in_r_bypass_2_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_2_stall_18 <= io_in_r_bypass_2_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_3_data_18 <= io_in_r_bypass_2_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_3_load_store_18 <= io_in_r_bypass_2_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_3_df_is_ws_18 <= io_in_r_bypass_2_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_3_stall_18 <= io_in_r_bypass_2_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_0_data_18 <= io_in_r_bypass_3_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_0_load_store_18 <= io_in_r_bypass_3_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_0_df_is_ws_18 <= io_in_r_bypass_3_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_0_stall_18 <= io_in_r_bypass_3_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_1_data_18 <= io_in_r_bypass_3_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_1_load_store_18 <= io_in_r_bypass_3_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_1_df_is_ws_18 <= io_in_r_bypass_3_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_1_stall_18 <= io_in_r_bypass_3_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_2_data_18 <= io_in_r_bypass_3_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_2_load_store_18 <= io_in_r_bypass_3_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_2_df_is_ws_18 <= io_in_r_bypass_3_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_2_stall_18 <= io_in_r_bypass_3_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_3_data_18 <= io_in_r_bypass_3_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_3_load_store_18 <= io_in_r_bypass_3_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_3_df_is_ws_18 <= io_in_r_bypass_3_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_3_stall_18 <= io_in_r_bypass_3_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_0_data_18 <= io_in_r_bypass_4_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_0_load_store_18 <= io_in_r_bypass_4_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_0_df_is_ws_18 <= io_in_r_bypass_4_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_0_stall_18 <= io_in_r_bypass_4_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_1_data_18 <= io_in_r_bypass_4_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_1_load_store_18 <= io_in_r_bypass_4_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_1_df_is_ws_18 <= io_in_r_bypass_4_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_1_stall_18 <= io_in_r_bypass_4_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_2_data_18 <= io_in_r_bypass_4_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_2_load_store_18 <= io_in_r_bypass_4_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_2_df_is_ws_18 <= io_in_r_bypass_4_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_2_stall_18 <= io_in_r_bypass_4_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_3_data_18 <= io_in_r_bypass_4_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_3_load_store_18 <= io_in_r_bypass_4_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_3_df_is_ws_18 <= io_in_r_bypass_4_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_3_stall_18 <= io_in_r_bypass_4_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_0_data_18 <= io_in_r_bypass_5_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_0_load_store_18 <= io_in_r_bypass_5_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_0_df_is_ws_18 <= io_in_r_bypass_5_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_0_stall_18 <= io_in_r_bypass_5_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_1_data_18 <= io_in_r_bypass_5_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_1_load_store_18 <= io_in_r_bypass_5_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_1_df_is_ws_18 <= io_in_r_bypass_5_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_1_stall_18 <= io_in_r_bypass_5_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_2_data_18 <= io_in_r_bypass_5_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_2_load_store_18 <= io_in_r_bypass_5_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_2_df_is_ws_18 <= io_in_r_bypass_5_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_2_stall_18 <= io_in_r_bypass_5_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_3_data_18 <= io_in_r_bypass_5_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_3_load_store_18 <= io_in_r_bypass_5_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_3_df_is_ws_18 <= io_in_r_bypass_5_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_3_stall_18 <= io_in_r_bypass_5_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_0_data_18 <= io_in_r_bypass_6_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_0_load_store_18 <= io_in_r_bypass_6_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_0_df_is_ws_18 <= io_in_r_bypass_6_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_0_stall_18 <= io_in_r_bypass_6_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_1_data_18 <= io_in_r_bypass_6_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_1_load_store_18 <= io_in_r_bypass_6_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_1_df_is_ws_18 <= io_in_r_bypass_6_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_1_stall_18 <= io_in_r_bypass_6_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_2_data_18 <= io_in_r_bypass_6_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_2_load_store_18 <= io_in_r_bypass_6_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_2_df_is_ws_18 <= io_in_r_bypass_6_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_2_stall_18 <= io_in_r_bypass_6_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_3_data_18 <= io_in_r_bypass_6_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_3_load_store_18 <= io_in_r_bypass_6_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_3_df_is_ws_18 <= io_in_r_bypass_6_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_3_stall_18 <= io_in_r_bypass_6_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_0_data_18 <= io_in_r_bypass_7_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_0_load_store_18 <= io_in_r_bypass_7_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_0_df_is_ws_18 <= io_in_r_bypass_7_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_0_stall_18 <= io_in_r_bypass_7_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_1_data_18 <= io_in_r_bypass_7_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_1_load_store_18 <= io_in_r_bypass_7_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_1_df_is_ws_18 <= io_in_r_bypass_7_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_1_stall_18 <= io_in_r_bypass_7_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_2_data_18 <= io_in_r_bypass_7_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_2_load_store_18 <= io_in_r_bypass_7_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_2_df_is_ws_18 <= io_in_r_bypass_7_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_2_stall_18 <= io_in_r_bypass_7_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_3_data_18 <= io_in_r_bypass_7_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_3_load_store_18 <= io_in_r_bypass_7_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_3_df_is_ws_18 <= io_in_r_bypass_7_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_3_stall_18 <= io_in_r_bypass_7_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_0_data_18 <= io_in_r_bypass_8_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_0_load_store_18 <= io_in_r_bypass_8_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_0_df_is_ws_18 <= io_in_r_bypass_8_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_0_stall_18 <= io_in_r_bypass_8_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_1_data_18 <= io_in_r_bypass_8_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_1_load_store_18 <= io_in_r_bypass_8_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_1_df_is_ws_18 <= io_in_r_bypass_8_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_1_stall_18 <= io_in_r_bypass_8_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_2_data_18 <= io_in_r_bypass_8_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_2_load_store_18 <= io_in_r_bypass_8_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_2_df_is_ws_18 <= io_in_r_bypass_8_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_2_stall_18 <= io_in_r_bypass_8_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_3_data_18 <= io_in_r_bypass_8_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_3_load_store_18 <= io_in_r_bypass_8_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_3_df_is_ws_18 <= io_in_r_bypass_8_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_3_stall_18 <= io_in_r_bypass_8_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_0_data_18 <= io_in_r_bypass_9_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_0_load_store_18 <= io_in_r_bypass_9_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_0_df_is_ws_18 <= io_in_r_bypass_9_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_0_stall_18 <= io_in_r_bypass_9_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_1_data_18 <= io_in_r_bypass_9_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_1_load_store_18 <= io_in_r_bypass_9_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_1_df_is_ws_18 <= io_in_r_bypass_9_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_1_stall_18 <= io_in_r_bypass_9_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_2_data_18 <= io_in_r_bypass_9_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_2_load_store_18 <= io_in_r_bypass_9_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_2_df_is_ws_18 <= io_in_r_bypass_9_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_2_stall_18 <= io_in_r_bypass_9_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_3_data_18 <= io_in_r_bypass_9_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_3_load_store_18 <= io_in_r_bypass_9_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_3_df_is_ws_18 <= io_in_r_bypass_9_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_3_stall_18 <= io_in_r_bypass_9_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_0_data_18 <= io_in_r_bypass_10_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_0_load_store_18 <= io_in_r_bypass_10_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_0_df_is_ws_18 <= io_in_r_bypass_10_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_0_stall_18 <= io_in_r_bypass_10_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_1_data_18 <= io_in_r_bypass_10_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_1_load_store_18 <= io_in_r_bypass_10_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_1_df_is_ws_18 <= io_in_r_bypass_10_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_1_stall_18 <= io_in_r_bypass_10_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_2_data_18 <= io_in_r_bypass_10_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_2_load_store_18 <= io_in_r_bypass_10_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_2_df_is_ws_18 <= io_in_r_bypass_10_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_2_stall_18 <= io_in_r_bypass_10_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_3_data_18 <= io_in_r_bypass_10_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_3_load_store_18 <= io_in_r_bypass_10_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_3_df_is_ws_18 <= io_in_r_bypass_10_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_3_stall_18 <= io_in_r_bypass_10_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_0_data_18 <= io_in_r_bypass_11_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_0_load_store_18 <= io_in_r_bypass_11_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_0_df_is_ws_18 <= io_in_r_bypass_11_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_0_stall_18 <= io_in_r_bypass_11_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_1_data_18 <= io_in_r_bypass_11_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_1_load_store_18 <= io_in_r_bypass_11_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_1_df_is_ws_18 <= io_in_r_bypass_11_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_1_stall_18 <= io_in_r_bypass_11_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_2_data_18 <= io_in_r_bypass_11_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_2_load_store_18 <= io_in_r_bypass_11_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_2_df_is_ws_18 <= io_in_r_bypass_11_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_2_stall_18 <= io_in_r_bypass_11_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_3_data_18 <= io_in_r_bypass_11_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_3_load_store_18 <= io_in_r_bypass_11_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_3_df_is_ws_18 <= io_in_r_bypass_11_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_3_stall_18 <= io_in_r_bypass_11_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_0_data_18 <= io_in_r_bypass_12_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_0_load_store_18 <= io_in_r_bypass_12_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_0_df_is_ws_18 <= io_in_r_bypass_12_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_0_stall_18 <= io_in_r_bypass_12_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_1_data_18 <= io_in_r_bypass_12_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_1_load_store_18 <= io_in_r_bypass_12_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_1_df_is_ws_18 <= io_in_r_bypass_12_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_1_stall_18 <= io_in_r_bypass_12_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_2_data_18 <= io_in_r_bypass_12_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_2_load_store_18 <= io_in_r_bypass_12_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_2_df_is_ws_18 <= io_in_r_bypass_12_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_2_stall_18 <= io_in_r_bypass_12_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_3_data_18 <= io_in_r_bypass_12_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_3_load_store_18 <= io_in_r_bypass_12_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_3_df_is_ws_18 <= io_in_r_bypass_12_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_3_stall_18 <= io_in_r_bypass_12_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_0_data_18 <= io_in_r_bypass_13_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_0_load_store_18 <= io_in_r_bypass_13_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_0_df_is_ws_18 <= io_in_r_bypass_13_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_0_stall_18 <= io_in_r_bypass_13_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_1_data_18 <= io_in_r_bypass_13_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_1_load_store_18 <= io_in_r_bypass_13_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_1_df_is_ws_18 <= io_in_r_bypass_13_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_1_stall_18 <= io_in_r_bypass_13_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_2_data_18 <= io_in_r_bypass_13_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_2_load_store_18 <= io_in_r_bypass_13_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_2_df_is_ws_18 <= io_in_r_bypass_13_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_2_stall_18 <= io_in_r_bypass_13_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_3_data_18 <= io_in_r_bypass_13_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_3_load_store_18 <= io_in_r_bypass_13_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_3_df_is_ws_18 <= io_in_r_bypass_13_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_3_stall_18 <= io_in_r_bypass_13_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_0_data_18 <= io_in_r_bypass_14_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_0_load_store_18 <= io_in_r_bypass_14_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_0_df_is_ws_18 <= io_in_r_bypass_14_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_0_stall_18 <= io_in_r_bypass_14_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_1_data_18 <= io_in_r_bypass_14_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_1_load_store_18 <= io_in_r_bypass_14_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_1_df_is_ws_18 <= io_in_r_bypass_14_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_1_stall_18 <= io_in_r_bypass_14_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_2_data_18 <= io_in_r_bypass_14_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_2_load_store_18 <= io_in_r_bypass_14_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_2_df_is_ws_18 <= io_in_r_bypass_14_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_2_stall_18 <= io_in_r_bypass_14_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_3_data_18 <= io_in_r_bypass_14_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_3_load_store_18 <= io_in_r_bypass_14_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_3_df_is_ws_18 <= io_in_r_bypass_14_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_3_stall_18 <= io_in_r_bypass_14_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_0_data_18 <= io_in_r_bypass_15_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_0_load_store_18 <= io_in_r_bypass_15_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_0_df_is_ws_18 <= io_in_r_bypass_15_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_0_stall_18 <= io_in_r_bypass_15_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_1_data_18 <= io_in_r_bypass_15_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_1_load_store_18 <= io_in_r_bypass_15_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_1_df_is_ws_18 <= io_in_r_bypass_15_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_1_stall_18 <= io_in_r_bypass_15_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_2_data_18 <= io_in_r_bypass_15_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_2_load_store_18 <= io_in_r_bypass_15_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_2_df_is_ws_18 <= io_in_r_bypass_15_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_2_stall_18 <= io_in_r_bypass_15_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_3_data_18 <= io_in_r_bypass_15_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_3_load_store_18 <= io_in_r_bypass_15_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_3_df_is_ws_18 <= io_in_r_bypass_15_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_3_stall_18 <= io_in_r_bypass_15_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_0_data_18 <= io_in_r_bypass_16_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_0_load_store_18 <= io_in_r_bypass_16_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_0_df_is_ws_18 <= io_in_r_bypass_16_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_0_stall_18 <= io_in_r_bypass_16_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_1_data_18 <= io_in_r_bypass_16_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_1_load_store_18 <= io_in_r_bypass_16_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_1_df_is_ws_18 <= io_in_r_bypass_16_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_1_stall_18 <= io_in_r_bypass_16_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_2_data_18 <= io_in_r_bypass_16_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_2_load_store_18 <= io_in_r_bypass_16_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_2_df_is_ws_18 <= io_in_r_bypass_16_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_2_stall_18 <= io_in_r_bypass_16_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_3_data_18 <= io_in_r_bypass_16_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_3_load_store_18 <= io_in_r_bypass_16_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_3_df_is_ws_18 <= io_in_r_bypass_16_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_3_stall_18 <= io_in_r_bypass_16_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_0_data_18 <= io_in_r_bypass_17_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_0_load_store_18 <= io_in_r_bypass_17_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_0_df_is_ws_18 <= io_in_r_bypass_17_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_0_stall_18 <= io_in_r_bypass_17_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_1_data_18 <= io_in_r_bypass_17_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_1_load_store_18 <= io_in_r_bypass_17_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_1_df_is_ws_18 <= io_in_r_bypass_17_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_1_stall_18 <= io_in_r_bypass_17_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_2_data_18 <= io_in_r_bypass_17_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_2_load_store_18 <= io_in_r_bypass_17_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_2_df_is_ws_18 <= io_in_r_bypass_17_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_2_stall_18 <= io_in_r_bypass_17_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_3_data_18 <= io_in_r_bypass_17_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_3_load_store_18 <= io_in_r_bypass_17_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_3_df_is_ws_18 <= io_in_r_bypass_17_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_3_stall_18 <= io_in_r_bypass_17_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_0_data_18 <= io_in_r_bypass_18_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_0_load_store_18 <= io_in_r_bypass_18_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_0_df_is_ws_18 <= io_in_r_bypass_18_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_0_stall_18 <= io_in_r_bypass_18_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_1_data_18 <= io_in_r_bypass_18_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_1_load_store_18 <= io_in_r_bypass_18_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_1_df_is_ws_18 <= io_in_r_bypass_18_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_1_stall_18 <= io_in_r_bypass_18_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_2_data_18 <= io_in_r_bypass_18_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_2_load_store_18 <= io_in_r_bypass_18_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_2_df_is_ws_18 <= io_in_r_bypass_18_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_2_stall_18 <= io_in_r_bypass_18_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_3_data_18 <= io_in_r_bypass_18_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_3_load_store_18 <= io_in_r_bypass_18_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_3_df_is_ws_18 <= io_in_r_bypass_18_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_3_stall_18 <= io_in_r_bypass_18_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_0_data_18 <= io_in_r_bypass_19_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_0_load_store_18 <= io_in_r_bypass_19_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_0_df_is_ws_18 <= io_in_r_bypass_19_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_0_stall_18 <= io_in_r_bypass_19_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_1_data_18 <= io_in_r_bypass_19_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_1_load_store_18 <= io_in_r_bypass_19_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_1_df_is_ws_18 <= io_in_r_bypass_19_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_1_stall_18 <= io_in_r_bypass_19_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_2_data_18 <= io_in_r_bypass_19_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_2_load_store_18 <= io_in_r_bypass_19_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_2_df_is_ws_18 <= io_in_r_bypass_19_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_2_stall_18 <= io_in_r_bypass_19_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_3_data_18 <= io_in_r_bypass_19_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_3_load_store_18 <= io_in_r_bypass_19_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_3_df_is_ws_18 <= io_in_r_bypass_19_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_3_stall_18 <= io_in_r_bypass_19_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_0_data_18 <= io_in_r_bypass_20_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_0_load_store_18 <= io_in_r_bypass_20_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_0_df_is_ws_18 <= io_in_r_bypass_20_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_0_stall_18 <= io_in_r_bypass_20_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_1_data_18 <= io_in_r_bypass_20_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_1_load_store_18 <= io_in_r_bypass_20_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_1_df_is_ws_18 <= io_in_r_bypass_20_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_1_stall_18 <= io_in_r_bypass_20_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_2_data_18 <= io_in_r_bypass_20_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_2_load_store_18 <= io_in_r_bypass_20_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_2_df_is_ws_18 <= io_in_r_bypass_20_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_2_stall_18 <= io_in_r_bypass_20_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_3_data_18 <= io_in_r_bypass_20_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_3_load_store_18 <= io_in_r_bypass_20_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_3_df_is_ws_18 <= io_in_r_bypass_20_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_3_stall_18 <= io_in_r_bypass_20_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_0_data_18 <= io_in_r_bypass_21_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_0_load_store_18 <= io_in_r_bypass_21_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_0_df_is_ws_18 <= io_in_r_bypass_21_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_0_stall_18 <= io_in_r_bypass_21_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_1_data_18 <= io_in_r_bypass_21_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_1_load_store_18 <= io_in_r_bypass_21_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_1_df_is_ws_18 <= io_in_r_bypass_21_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_1_stall_18 <= io_in_r_bypass_21_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_2_data_18 <= io_in_r_bypass_21_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_2_load_store_18 <= io_in_r_bypass_21_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_2_df_is_ws_18 <= io_in_r_bypass_21_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_2_stall_18 <= io_in_r_bypass_21_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_3_data_18 <= io_in_r_bypass_21_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_3_load_store_18 <= io_in_r_bypass_21_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_3_df_is_ws_18 <= io_in_r_bypass_21_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_3_stall_18 <= io_in_r_bypass_21_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_0_data_18 <= io_in_r_bypass_22_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_0_load_store_18 <= io_in_r_bypass_22_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_0_df_is_ws_18 <= io_in_r_bypass_22_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_0_stall_18 <= io_in_r_bypass_22_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_1_data_18 <= io_in_r_bypass_22_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_1_load_store_18 <= io_in_r_bypass_22_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_1_df_is_ws_18 <= io_in_r_bypass_22_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_1_stall_18 <= io_in_r_bypass_22_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_2_data_18 <= io_in_r_bypass_22_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_2_load_store_18 <= io_in_r_bypass_22_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_2_df_is_ws_18 <= io_in_r_bypass_22_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_2_stall_18 <= io_in_r_bypass_22_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_3_data_18 <= io_in_r_bypass_22_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_3_load_store_18 <= io_in_r_bypass_22_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_3_df_is_ws_18 <= io_in_r_bypass_22_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_3_stall_18 <= io_in_r_bypass_22_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_0_data_18 <= io_in_r_bypass_23_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_0_load_store_18 <= io_in_r_bypass_23_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_0_df_is_ws_18 <= io_in_r_bypass_23_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_0_stall_18 <= io_in_r_bypass_23_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_1_data_18 <= io_in_r_bypass_23_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_1_load_store_18 <= io_in_r_bypass_23_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_1_df_is_ws_18 <= io_in_r_bypass_23_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_1_stall_18 <= io_in_r_bypass_23_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_2_data_18 <= io_in_r_bypass_23_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_2_load_store_18 <= io_in_r_bypass_23_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_2_df_is_ws_18 <= io_in_r_bypass_23_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_2_stall_18 <= io_in_r_bypass_23_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_3_data_18 <= io_in_r_bypass_23_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_3_load_store_18 <= io_in_r_bypass_23_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_3_df_is_ws_18 <= io_in_r_bypass_23_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_3_stall_18 <= io_in_r_bypass_23_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_0_data_18 <= io_in_r_bypass_24_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_0_load_store_18 <= io_in_r_bypass_24_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_0_df_is_ws_18 <= io_in_r_bypass_24_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_0_stall_18 <= io_in_r_bypass_24_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_1_data_18 <= io_in_r_bypass_24_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_1_load_store_18 <= io_in_r_bypass_24_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_1_df_is_ws_18 <= io_in_r_bypass_24_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_1_stall_18 <= io_in_r_bypass_24_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_2_data_18 <= io_in_r_bypass_24_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_2_load_store_18 <= io_in_r_bypass_24_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_2_df_is_ws_18 <= io_in_r_bypass_24_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_2_stall_18 <= io_in_r_bypass_24_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_3_data_18 <= io_in_r_bypass_24_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_3_load_store_18 <= io_in_r_bypass_24_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_3_df_is_ws_18 <= io_in_r_bypass_24_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_3_stall_18 <= io_in_r_bypass_24_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_0_data_18 <= io_in_r_bypass_25_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_0_load_store_18 <= io_in_r_bypass_25_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_0_df_is_ws_18 <= io_in_r_bypass_25_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_0_stall_18 <= io_in_r_bypass_25_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_1_data_18 <= io_in_r_bypass_25_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_1_load_store_18 <= io_in_r_bypass_25_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_1_df_is_ws_18 <= io_in_r_bypass_25_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_1_stall_18 <= io_in_r_bypass_25_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_2_data_18 <= io_in_r_bypass_25_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_2_load_store_18 <= io_in_r_bypass_25_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_2_df_is_ws_18 <= io_in_r_bypass_25_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_2_stall_18 <= io_in_r_bypass_25_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_3_data_18 <= io_in_r_bypass_25_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_3_load_store_18 <= io_in_r_bypass_25_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_3_df_is_ws_18 <= io_in_r_bypass_25_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_3_stall_18 <= io_in_r_bypass_25_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_0_data_18 <= io_in_r_bypass_26_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_0_load_store_18 <= io_in_r_bypass_26_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_0_df_is_ws_18 <= io_in_r_bypass_26_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_0_stall_18 <= io_in_r_bypass_26_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_1_data_18 <= io_in_r_bypass_26_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_1_load_store_18 <= io_in_r_bypass_26_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_1_df_is_ws_18 <= io_in_r_bypass_26_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_1_stall_18 <= io_in_r_bypass_26_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_2_data_18 <= io_in_r_bypass_26_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_2_load_store_18 <= io_in_r_bypass_26_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_2_df_is_ws_18 <= io_in_r_bypass_26_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_2_stall_18 <= io_in_r_bypass_26_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_3_data_18 <= io_in_r_bypass_26_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_3_load_store_18 <= io_in_r_bypass_26_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_3_df_is_ws_18 <= io_in_r_bypass_26_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_3_stall_18 <= io_in_r_bypass_26_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_0_data_18 <= io_in_r_bypass_27_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_0_load_store_18 <= io_in_r_bypass_27_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_0_df_is_ws_18 <= io_in_r_bypass_27_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_0_stall_18 <= io_in_r_bypass_27_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_1_data_18 <= io_in_r_bypass_27_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_1_load_store_18 <= io_in_r_bypass_27_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_1_df_is_ws_18 <= io_in_r_bypass_27_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_1_stall_18 <= io_in_r_bypass_27_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_2_data_18 <= io_in_r_bypass_27_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_2_load_store_18 <= io_in_r_bypass_27_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_2_df_is_ws_18 <= io_in_r_bypass_27_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_2_stall_18 <= io_in_r_bypass_27_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_3_data_18 <= io_in_r_bypass_27_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_3_load_store_18 <= io_in_r_bypass_27_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_3_df_is_ws_18 <= io_in_r_bypass_27_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_3_stall_18 <= io_in_r_bypass_27_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_0_data_18 <= io_in_r_bypass_28_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_0_load_store_18 <= io_in_r_bypass_28_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_0_df_is_ws_18 <= io_in_r_bypass_28_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_0_stall_18 <= io_in_r_bypass_28_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_1_data_18 <= io_in_r_bypass_28_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_1_load_store_18 <= io_in_r_bypass_28_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_1_df_is_ws_18 <= io_in_r_bypass_28_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_1_stall_18 <= io_in_r_bypass_28_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_2_data_18 <= io_in_r_bypass_28_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_2_load_store_18 <= io_in_r_bypass_28_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_2_df_is_ws_18 <= io_in_r_bypass_28_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_2_stall_18 <= io_in_r_bypass_28_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_3_data_18 <= io_in_r_bypass_28_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_3_load_store_18 <= io_in_r_bypass_28_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_3_df_is_ws_18 <= io_in_r_bypass_28_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_3_stall_18 <= io_in_r_bypass_28_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_0_data_18 <= io_in_r_bypass_29_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_0_load_store_18 <= io_in_r_bypass_29_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_0_df_is_ws_18 <= io_in_r_bypass_29_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_0_stall_18 <= io_in_r_bypass_29_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_1_data_18 <= io_in_r_bypass_29_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_1_load_store_18 <= io_in_r_bypass_29_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_1_df_is_ws_18 <= io_in_r_bypass_29_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_1_stall_18 <= io_in_r_bypass_29_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_2_data_18 <= io_in_r_bypass_29_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_2_load_store_18 <= io_in_r_bypass_29_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_2_df_is_ws_18 <= io_in_r_bypass_29_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_2_stall_18 <= io_in_r_bypass_29_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_3_data_18 <= io_in_r_bypass_29_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_3_load_store_18 <= io_in_r_bypass_29_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_3_df_is_ws_18 <= io_in_r_bypass_29_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_3_stall_18 <= io_in_r_bypass_29_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_0_data_18 <= io_in_r_bypass_30_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_0_load_store_18 <= io_in_r_bypass_30_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_0_df_is_ws_18 <= io_in_r_bypass_30_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_0_stall_18 <= io_in_r_bypass_30_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_1_data_18 <= io_in_r_bypass_30_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_1_load_store_18 <= io_in_r_bypass_30_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_1_df_is_ws_18 <= io_in_r_bypass_30_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_1_stall_18 <= io_in_r_bypass_30_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_2_data_18 <= io_in_r_bypass_30_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_2_load_store_18 <= io_in_r_bypass_30_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_2_df_is_ws_18 <= io_in_r_bypass_30_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_2_stall_18 <= io_in_r_bypass_30_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_3_data_18 <= io_in_r_bypass_30_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_3_load_store_18 <= io_in_r_bypass_30_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_3_df_is_ws_18 <= io_in_r_bypass_30_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_3_stall_18 <= io_in_r_bypass_30_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_0_data_18 <= io_in_r_bypass_31_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_0_load_store_18 <= io_in_r_bypass_31_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_0_df_is_ws_18 <= io_in_r_bypass_31_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_0_stall_18 <= io_in_r_bypass_31_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_1_data_18 <= io_in_r_bypass_31_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_1_load_store_18 <= io_in_r_bypass_31_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_1_df_is_ws_18 <= io_in_r_bypass_31_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_1_stall_18 <= io_in_r_bypass_31_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_2_data_18 <= io_in_r_bypass_31_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_2_load_store_18 <= io_in_r_bypass_31_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_2_df_is_ws_18 <= io_in_r_bypass_31_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_2_stall_18 <= io_in_r_bypass_31_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_3_data_18 <= io_in_r_bypass_31_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_3_load_store_18 <= io_in_r_bypass_31_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_3_df_is_ws_18 <= io_in_r_bypass_31_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_3_stall_18 <= io_in_r_bypass_31_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_0_data_19 <= io_in_r_bypass_0_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_0_load_store_19 <= io_in_r_bypass_0_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_0_df_is_ws_19 <= io_in_r_bypass_0_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_0_stall_19 <= io_in_r_bypass_0_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_1_data_19 <= io_in_r_bypass_0_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_1_load_store_19 <= io_in_r_bypass_0_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_1_df_is_ws_19 <= io_in_r_bypass_0_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_1_stall_19 <= io_in_r_bypass_0_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_2_data_19 <= io_in_r_bypass_0_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_2_load_store_19 <= io_in_r_bypass_0_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_2_df_is_ws_19 <= io_in_r_bypass_0_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_2_stall_19 <= io_in_r_bypass_0_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_3_data_19 <= io_in_r_bypass_0_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_3_load_store_19 <= io_in_r_bypass_0_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_3_df_is_ws_19 <= io_in_r_bypass_0_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_3_stall_19 <= io_in_r_bypass_0_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_0_data_19 <= io_in_r_bypass_1_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_0_load_store_19 <= io_in_r_bypass_1_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_0_df_is_ws_19 <= io_in_r_bypass_1_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_0_stall_19 <= io_in_r_bypass_1_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_1_data_19 <= io_in_r_bypass_1_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_1_load_store_19 <= io_in_r_bypass_1_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_1_df_is_ws_19 <= io_in_r_bypass_1_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_1_stall_19 <= io_in_r_bypass_1_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_2_data_19 <= io_in_r_bypass_1_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_2_load_store_19 <= io_in_r_bypass_1_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_2_df_is_ws_19 <= io_in_r_bypass_1_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_2_stall_19 <= io_in_r_bypass_1_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_3_data_19 <= io_in_r_bypass_1_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_3_load_store_19 <= io_in_r_bypass_1_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_3_df_is_ws_19 <= io_in_r_bypass_1_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_3_stall_19 <= io_in_r_bypass_1_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_0_data_19 <= io_in_r_bypass_2_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_0_load_store_19 <= io_in_r_bypass_2_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_0_df_is_ws_19 <= io_in_r_bypass_2_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_0_stall_19 <= io_in_r_bypass_2_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_1_data_19 <= io_in_r_bypass_2_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_1_load_store_19 <= io_in_r_bypass_2_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_1_df_is_ws_19 <= io_in_r_bypass_2_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_1_stall_19 <= io_in_r_bypass_2_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_2_data_19 <= io_in_r_bypass_2_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_2_load_store_19 <= io_in_r_bypass_2_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_2_df_is_ws_19 <= io_in_r_bypass_2_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_2_stall_19 <= io_in_r_bypass_2_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_3_data_19 <= io_in_r_bypass_2_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_3_load_store_19 <= io_in_r_bypass_2_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_3_df_is_ws_19 <= io_in_r_bypass_2_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_3_stall_19 <= io_in_r_bypass_2_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_0_data_19 <= io_in_r_bypass_3_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_0_load_store_19 <= io_in_r_bypass_3_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_0_df_is_ws_19 <= io_in_r_bypass_3_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_0_stall_19 <= io_in_r_bypass_3_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_1_data_19 <= io_in_r_bypass_3_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_1_load_store_19 <= io_in_r_bypass_3_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_1_df_is_ws_19 <= io_in_r_bypass_3_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_1_stall_19 <= io_in_r_bypass_3_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_2_data_19 <= io_in_r_bypass_3_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_2_load_store_19 <= io_in_r_bypass_3_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_2_df_is_ws_19 <= io_in_r_bypass_3_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_2_stall_19 <= io_in_r_bypass_3_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_3_data_19 <= io_in_r_bypass_3_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_3_load_store_19 <= io_in_r_bypass_3_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_3_df_is_ws_19 <= io_in_r_bypass_3_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_3_stall_19 <= io_in_r_bypass_3_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_0_data_19 <= io_in_r_bypass_4_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_0_load_store_19 <= io_in_r_bypass_4_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_0_df_is_ws_19 <= io_in_r_bypass_4_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_0_stall_19 <= io_in_r_bypass_4_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_1_data_19 <= io_in_r_bypass_4_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_1_load_store_19 <= io_in_r_bypass_4_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_1_df_is_ws_19 <= io_in_r_bypass_4_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_1_stall_19 <= io_in_r_bypass_4_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_2_data_19 <= io_in_r_bypass_4_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_2_load_store_19 <= io_in_r_bypass_4_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_2_df_is_ws_19 <= io_in_r_bypass_4_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_2_stall_19 <= io_in_r_bypass_4_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_3_data_19 <= io_in_r_bypass_4_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_3_load_store_19 <= io_in_r_bypass_4_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_3_df_is_ws_19 <= io_in_r_bypass_4_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_3_stall_19 <= io_in_r_bypass_4_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_0_data_19 <= io_in_r_bypass_5_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_0_load_store_19 <= io_in_r_bypass_5_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_0_df_is_ws_19 <= io_in_r_bypass_5_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_0_stall_19 <= io_in_r_bypass_5_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_1_data_19 <= io_in_r_bypass_5_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_1_load_store_19 <= io_in_r_bypass_5_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_1_df_is_ws_19 <= io_in_r_bypass_5_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_1_stall_19 <= io_in_r_bypass_5_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_2_data_19 <= io_in_r_bypass_5_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_2_load_store_19 <= io_in_r_bypass_5_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_2_df_is_ws_19 <= io_in_r_bypass_5_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_2_stall_19 <= io_in_r_bypass_5_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_3_data_19 <= io_in_r_bypass_5_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_3_load_store_19 <= io_in_r_bypass_5_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_3_df_is_ws_19 <= io_in_r_bypass_5_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_3_stall_19 <= io_in_r_bypass_5_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_0_data_19 <= io_in_r_bypass_6_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_0_load_store_19 <= io_in_r_bypass_6_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_0_df_is_ws_19 <= io_in_r_bypass_6_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_0_stall_19 <= io_in_r_bypass_6_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_1_data_19 <= io_in_r_bypass_6_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_1_load_store_19 <= io_in_r_bypass_6_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_1_df_is_ws_19 <= io_in_r_bypass_6_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_1_stall_19 <= io_in_r_bypass_6_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_2_data_19 <= io_in_r_bypass_6_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_2_load_store_19 <= io_in_r_bypass_6_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_2_df_is_ws_19 <= io_in_r_bypass_6_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_2_stall_19 <= io_in_r_bypass_6_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_3_data_19 <= io_in_r_bypass_6_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_3_load_store_19 <= io_in_r_bypass_6_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_3_df_is_ws_19 <= io_in_r_bypass_6_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_3_stall_19 <= io_in_r_bypass_6_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_0_data_19 <= io_in_r_bypass_7_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_0_load_store_19 <= io_in_r_bypass_7_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_0_df_is_ws_19 <= io_in_r_bypass_7_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_0_stall_19 <= io_in_r_bypass_7_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_1_data_19 <= io_in_r_bypass_7_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_1_load_store_19 <= io_in_r_bypass_7_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_1_df_is_ws_19 <= io_in_r_bypass_7_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_1_stall_19 <= io_in_r_bypass_7_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_2_data_19 <= io_in_r_bypass_7_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_2_load_store_19 <= io_in_r_bypass_7_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_2_df_is_ws_19 <= io_in_r_bypass_7_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_2_stall_19 <= io_in_r_bypass_7_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_3_data_19 <= io_in_r_bypass_7_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_3_load_store_19 <= io_in_r_bypass_7_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_3_df_is_ws_19 <= io_in_r_bypass_7_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_3_stall_19 <= io_in_r_bypass_7_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_0_data_19 <= io_in_r_bypass_8_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_0_load_store_19 <= io_in_r_bypass_8_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_0_df_is_ws_19 <= io_in_r_bypass_8_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_0_stall_19 <= io_in_r_bypass_8_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_1_data_19 <= io_in_r_bypass_8_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_1_load_store_19 <= io_in_r_bypass_8_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_1_df_is_ws_19 <= io_in_r_bypass_8_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_1_stall_19 <= io_in_r_bypass_8_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_2_data_19 <= io_in_r_bypass_8_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_2_load_store_19 <= io_in_r_bypass_8_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_2_df_is_ws_19 <= io_in_r_bypass_8_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_2_stall_19 <= io_in_r_bypass_8_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_3_data_19 <= io_in_r_bypass_8_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_3_load_store_19 <= io_in_r_bypass_8_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_3_df_is_ws_19 <= io_in_r_bypass_8_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_3_stall_19 <= io_in_r_bypass_8_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_0_data_19 <= io_in_r_bypass_9_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_0_load_store_19 <= io_in_r_bypass_9_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_0_df_is_ws_19 <= io_in_r_bypass_9_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_0_stall_19 <= io_in_r_bypass_9_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_1_data_19 <= io_in_r_bypass_9_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_1_load_store_19 <= io_in_r_bypass_9_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_1_df_is_ws_19 <= io_in_r_bypass_9_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_1_stall_19 <= io_in_r_bypass_9_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_2_data_19 <= io_in_r_bypass_9_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_2_load_store_19 <= io_in_r_bypass_9_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_2_df_is_ws_19 <= io_in_r_bypass_9_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_2_stall_19 <= io_in_r_bypass_9_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_3_data_19 <= io_in_r_bypass_9_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_3_load_store_19 <= io_in_r_bypass_9_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_3_df_is_ws_19 <= io_in_r_bypass_9_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_3_stall_19 <= io_in_r_bypass_9_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_0_data_19 <= io_in_r_bypass_10_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_0_load_store_19 <= io_in_r_bypass_10_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_0_df_is_ws_19 <= io_in_r_bypass_10_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_0_stall_19 <= io_in_r_bypass_10_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_1_data_19 <= io_in_r_bypass_10_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_1_load_store_19 <= io_in_r_bypass_10_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_1_df_is_ws_19 <= io_in_r_bypass_10_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_1_stall_19 <= io_in_r_bypass_10_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_2_data_19 <= io_in_r_bypass_10_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_2_load_store_19 <= io_in_r_bypass_10_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_2_df_is_ws_19 <= io_in_r_bypass_10_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_2_stall_19 <= io_in_r_bypass_10_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_3_data_19 <= io_in_r_bypass_10_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_3_load_store_19 <= io_in_r_bypass_10_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_3_df_is_ws_19 <= io_in_r_bypass_10_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_3_stall_19 <= io_in_r_bypass_10_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_0_data_19 <= io_in_r_bypass_11_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_0_load_store_19 <= io_in_r_bypass_11_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_0_df_is_ws_19 <= io_in_r_bypass_11_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_0_stall_19 <= io_in_r_bypass_11_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_1_data_19 <= io_in_r_bypass_11_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_1_load_store_19 <= io_in_r_bypass_11_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_1_df_is_ws_19 <= io_in_r_bypass_11_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_1_stall_19 <= io_in_r_bypass_11_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_2_data_19 <= io_in_r_bypass_11_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_2_load_store_19 <= io_in_r_bypass_11_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_2_df_is_ws_19 <= io_in_r_bypass_11_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_2_stall_19 <= io_in_r_bypass_11_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_3_data_19 <= io_in_r_bypass_11_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_3_load_store_19 <= io_in_r_bypass_11_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_3_df_is_ws_19 <= io_in_r_bypass_11_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_3_stall_19 <= io_in_r_bypass_11_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_0_data_19 <= io_in_r_bypass_12_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_0_load_store_19 <= io_in_r_bypass_12_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_0_df_is_ws_19 <= io_in_r_bypass_12_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_0_stall_19 <= io_in_r_bypass_12_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_1_data_19 <= io_in_r_bypass_12_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_1_load_store_19 <= io_in_r_bypass_12_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_1_df_is_ws_19 <= io_in_r_bypass_12_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_1_stall_19 <= io_in_r_bypass_12_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_2_data_19 <= io_in_r_bypass_12_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_2_load_store_19 <= io_in_r_bypass_12_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_2_df_is_ws_19 <= io_in_r_bypass_12_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_2_stall_19 <= io_in_r_bypass_12_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_3_data_19 <= io_in_r_bypass_12_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_3_load_store_19 <= io_in_r_bypass_12_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_3_df_is_ws_19 <= io_in_r_bypass_12_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_3_stall_19 <= io_in_r_bypass_12_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_0_data_19 <= io_in_r_bypass_13_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_0_load_store_19 <= io_in_r_bypass_13_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_0_df_is_ws_19 <= io_in_r_bypass_13_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_0_stall_19 <= io_in_r_bypass_13_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_1_data_19 <= io_in_r_bypass_13_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_1_load_store_19 <= io_in_r_bypass_13_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_1_df_is_ws_19 <= io_in_r_bypass_13_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_1_stall_19 <= io_in_r_bypass_13_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_2_data_19 <= io_in_r_bypass_13_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_2_load_store_19 <= io_in_r_bypass_13_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_2_df_is_ws_19 <= io_in_r_bypass_13_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_2_stall_19 <= io_in_r_bypass_13_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_3_data_19 <= io_in_r_bypass_13_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_3_load_store_19 <= io_in_r_bypass_13_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_3_df_is_ws_19 <= io_in_r_bypass_13_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_3_stall_19 <= io_in_r_bypass_13_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_0_data_19 <= io_in_r_bypass_14_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_0_load_store_19 <= io_in_r_bypass_14_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_0_df_is_ws_19 <= io_in_r_bypass_14_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_0_stall_19 <= io_in_r_bypass_14_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_1_data_19 <= io_in_r_bypass_14_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_1_load_store_19 <= io_in_r_bypass_14_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_1_df_is_ws_19 <= io_in_r_bypass_14_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_1_stall_19 <= io_in_r_bypass_14_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_2_data_19 <= io_in_r_bypass_14_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_2_load_store_19 <= io_in_r_bypass_14_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_2_df_is_ws_19 <= io_in_r_bypass_14_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_2_stall_19 <= io_in_r_bypass_14_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_3_data_19 <= io_in_r_bypass_14_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_3_load_store_19 <= io_in_r_bypass_14_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_3_df_is_ws_19 <= io_in_r_bypass_14_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_3_stall_19 <= io_in_r_bypass_14_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_0_data_19 <= io_in_r_bypass_15_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_0_load_store_19 <= io_in_r_bypass_15_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_0_df_is_ws_19 <= io_in_r_bypass_15_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_0_stall_19 <= io_in_r_bypass_15_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_1_data_19 <= io_in_r_bypass_15_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_1_load_store_19 <= io_in_r_bypass_15_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_1_df_is_ws_19 <= io_in_r_bypass_15_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_1_stall_19 <= io_in_r_bypass_15_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_2_data_19 <= io_in_r_bypass_15_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_2_load_store_19 <= io_in_r_bypass_15_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_2_df_is_ws_19 <= io_in_r_bypass_15_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_2_stall_19 <= io_in_r_bypass_15_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_3_data_19 <= io_in_r_bypass_15_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_3_load_store_19 <= io_in_r_bypass_15_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_3_df_is_ws_19 <= io_in_r_bypass_15_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_3_stall_19 <= io_in_r_bypass_15_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_0_data_19 <= io_in_r_bypass_16_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_0_load_store_19 <= io_in_r_bypass_16_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_0_df_is_ws_19 <= io_in_r_bypass_16_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_0_stall_19 <= io_in_r_bypass_16_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_1_data_19 <= io_in_r_bypass_16_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_1_load_store_19 <= io_in_r_bypass_16_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_1_df_is_ws_19 <= io_in_r_bypass_16_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_1_stall_19 <= io_in_r_bypass_16_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_2_data_19 <= io_in_r_bypass_16_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_2_load_store_19 <= io_in_r_bypass_16_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_2_df_is_ws_19 <= io_in_r_bypass_16_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_2_stall_19 <= io_in_r_bypass_16_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_3_data_19 <= io_in_r_bypass_16_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_3_load_store_19 <= io_in_r_bypass_16_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_3_df_is_ws_19 <= io_in_r_bypass_16_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_3_stall_19 <= io_in_r_bypass_16_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_0_data_19 <= io_in_r_bypass_17_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_0_load_store_19 <= io_in_r_bypass_17_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_0_df_is_ws_19 <= io_in_r_bypass_17_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_0_stall_19 <= io_in_r_bypass_17_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_1_data_19 <= io_in_r_bypass_17_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_1_load_store_19 <= io_in_r_bypass_17_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_1_df_is_ws_19 <= io_in_r_bypass_17_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_1_stall_19 <= io_in_r_bypass_17_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_2_data_19 <= io_in_r_bypass_17_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_2_load_store_19 <= io_in_r_bypass_17_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_2_df_is_ws_19 <= io_in_r_bypass_17_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_2_stall_19 <= io_in_r_bypass_17_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_3_data_19 <= io_in_r_bypass_17_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_3_load_store_19 <= io_in_r_bypass_17_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_3_df_is_ws_19 <= io_in_r_bypass_17_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_3_stall_19 <= io_in_r_bypass_17_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_0_data_19 <= io_in_r_bypass_18_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_0_load_store_19 <= io_in_r_bypass_18_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_0_df_is_ws_19 <= io_in_r_bypass_18_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_0_stall_19 <= io_in_r_bypass_18_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_1_data_19 <= io_in_r_bypass_18_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_1_load_store_19 <= io_in_r_bypass_18_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_1_df_is_ws_19 <= io_in_r_bypass_18_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_1_stall_19 <= io_in_r_bypass_18_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_2_data_19 <= io_in_r_bypass_18_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_2_load_store_19 <= io_in_r_bypass_18_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_2_df_is_ws_19 <= io_in_r_bypass_18_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_2_stall_19 <= io_in_r_bypass_18_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_3_data_19 <= io_in_r_bypass_18_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_3_load_store_19 <= io_in_r_bypass_18_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_3_df_is_ws_19 <= io_in_r_bypass_18_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_3_stall_19 <= io_in_r_bypass_18_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_0_data_19 <= io_in_r_bypass_19_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_0_load_store_19 <= io_in_r_bypass_19_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_0_df_is_ws_19 <= io_in_r_bypass_19_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_0_stall_19 <= io_in_r_bypass_19_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_1_data_19 <= io_in_r_bypass_19_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_1_load_store_19 <= io_in_r_bypass_19_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_1_df_is_ws_19 <= io_in_r_bypass_19_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_1_stall_19 <= io_in_r_bypass_19_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_2_data_19 <= io_in_r_bypass_19_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_2_load_store_19 <= io_in_r_bypass_19_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_2_df_is_ws_19 <= io_in_r_bypass_19_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_2_stall_19 <= io_in_r_bypass_19_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_3_data_19 <= io_in_r_bypass_19_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_3_load_store_19 <= io_in_r_bypass_19_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_3_df_is_ws_19 <= io_in_r_bypass_19_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_3_stall_19 <= io_in_r_bypass_19_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_0_data_19 <= io_in_r_bypass_20_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_0_load_store_19 <= io_in_r_bypass_20_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_0_df_is_ws_19 <= io_in_r_bypass_20_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_0_stall_19 <= io_in_r_bypass_20_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_1_data_19 <= io_in_r_bypass_20_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_1_load_store_19 <= io_in_r_bypass_20_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_1_df_is_ws_19 <= io_in_r_bypass_20_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_1_stall_19 <= io_in_r_bypass_20_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_2_data_19 <= io_in_r_bypass_20_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_2_load_store_19 <= io_in_r_bypass_20_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_2_df_is_ws_19 <= io_in_r_bypass_20_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_2_stall_19 <= io_in_r_bypass_20_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_3_data_19 <= io_in_r_bypass_20_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_3_load_store_19 <= io_in_r_bypass_20_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_3_df_is_ws_19 <= io_in_r_bypass_20_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_3_stall_19 <= io_in_r_bypass_20_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_0_data_19 <= io_in_r_bypass_21_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_0_load_store_19 <= io_in_r_bypass_21_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_0_df_is_ws_19 <= io_in_r_bypass_21_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_0_stall_19 <= io_in_r_bypass_21_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_1_data_19 <= io_in_r_bypass_21_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_1_load_store_19 <= io_in_r_bypass_21_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_1_df_is_ws_19 <= io_in_r_bypass_21_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_1_stall_19 <= io_in_r_bypass_21_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_2_data_19 <= io_in_r_bypass_21_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_2_load_store_19 <= io_in_r_bypass_21_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_2_df_is_ws_19 <= io_in_r_bypass_21_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_2_stall_19 <= io_in_r_bypass_21_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_3_data_19 <= io_in_r_bypass_21_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_3_load_store_19 <= io_in_r_bypass_21_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_3_df_is_ws_19 <= io_in_r_bypass_21_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_3_stall_19 <= io_in_r_bypass_21_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_0_data_19 <= io_in_r_bypass_22_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_0_load_store_19 <= io_in_r_bypass_22_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_0_df_is_ws_19 <= io_in_r_bypass_22_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_0_stall_19 <= io_in_r_bypass_22_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_1_data_19 <= io_in_r_bypass_22_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_1_load_store_19 <= io_in_r_bypass_22_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_1_df_is_ws_19 <= io_in_r_bypass_22_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_1_stall_19 <= io_in_r_bypass_22_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_2_data_19 <= io_in_r_bypass_22_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_2_load_store_19 <= io_in_r_bypass_22_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_2_df_is_ws_19 <= io_in_r_bypass_22_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_2_stall_19 <= io_in_r_bypass_22_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_3_data_19 <= io_in_r_bypass_22_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_3_load_store_19 <= io_in_r_bypass_22_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_3_df_is_ws_19 <= io_in_r_bypass_22_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_3_stall_19 <= io_in_r_bypass_22_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_0_data_19 <= io_in_r_bypass_23_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_0_load_store_19 <= io_in_r_bypass_23_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_0_df_is_ws_19 <= io_in_r_bypass_23_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_0_stall_19 <= io_in_r_bypass_23_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_1_data_19 <= io_in_r_bypass_23_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_1_load_store_19 <= io_in_r_bypass_23_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_1_df_is_ws_19 <= io_in_r_bypass_23_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_1_stall_19 <= io_in_r_bypass_23_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_2_data_19 <= io_in_r_bypass_23_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_2_load_store_19 <= io_in_r_bypass_23_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_2_df_is_ws_19 <= io_in_r_bypass_23_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_2_stall_19 <= io_in_r_bypass_23_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_3_data_19 <= io_in_r_bypass_23_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_3_load_store_19 <= io_in_r_bypass_23_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_3_df_is_ws_19 <= io_in_r_bypass_23_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_3_stall_19 <= io_in_r_bypass_23_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_0_data_19 <= io_in_r_bypass_24_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_0_load_store_19 <= io_in_r_bypass_24_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_0_df_is_ws_19 <= io_in_r_bypass_24_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_0_stall_19 <= io_in_r_bypass_24_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_1_data_19 <= io_in_r_bypass_24_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_1_load_store_19 <= io_in_r_bypass_24_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_1_df_is_ws_19 <= io_in_r_bypass_24_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_1_stall_19 <= io_in_r_bypass_24_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_2_data_19 <= io_in_r_bypass_24_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_2_load_store_19 <= io_in_r_bypass_24_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_2_df_is_ws_19 <= io_in_r_bypass_24_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_2_stall_19 <= io_in_r_bypass_24_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_3_data_19 <= io_in_r_bypass_24_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_3_load_store_19 <= io_in_r_bypass_24_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_3_df_is_ws_19 <= io_in_r_bypass_24_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_3_stall_19 <= io_in_r_bypass_24_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_0_data_19 <= io_in_r_bypass_25_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_0_load_store_19 <= io_in_r_bypass_25_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_0_df_is_ws_19 <= io_in_r_bypass_25_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_0_stall_19 <= io_in_r_bypass_25_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_1_data_19 <= io_in_r_bypass_25_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_1_load_store_19 <= io_in_r_bypass_25_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_1_df_is_ws_19 <= io_in_r_bypass_25_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_1_stall_19 <= io_in_r_bypass_25_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_2_data_19 <= io_in_r_bypass_25_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_2_load_store_19 <= io_in_r_bypass_25_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_2_df_is_ws_19 <= io_in_r_bypass_25_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_2_stall_19 <= io_in_r_bypass_25_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_3_data_19 <= io_in_r_bypass_25_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_3_load_store_19 <= io_in_r_bypass_25_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_3_df_is_ws_19 <= io_in_r_bypass_25_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_3_stall_19 <= io_in_r_bypass_25_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_0_data_19 <= io_in_r_bypass_26_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_0_load_store_19 <= io_in_r_bypass_26_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_0_df_is_ws_19 <= io_in_r_bypass_26_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_0_stall_19 <= io_in_r_bypass_26_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_1_data_19 <= io_in_r_bypass_26_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_1_load_store_19 <= io_in_r_bypass_26_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_1_df_is_ws_19 <= io_in_r_bypass_26_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_1_stall_19 <= io_in_r_bypass_26_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_2_data_19 <= io_in_r_bypass_26_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_2_load_store_19 <= io_in_r_bypass_26_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_2_df_is_ws_19 <= io_in_r_bypass_26_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_2_stall_19 <= io_in_r_bypass_26_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_3_data_19 <= io_in_r_bypass_26_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_3_load_store_19 <= io_in_r_bypass_26_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_3_df_is_ws_19 <= io_in_r_bypass_26_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_3_stall_19 <= io_in_r_bypass_26_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_0_data_19 <= io_in_r_bypass_27_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_0_load_store_19 <= io_in_r_bypass_27_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_0_df_is_ws_19 <= io_in_r_bypass_27_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_0_stall_19 <= io_in_r_bypass_27_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_1_data_19 <= io_in_r_bypass_27_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_1_load_store_19 <= io_in_r_bypass_27_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_1_df_is_ws_19 <= io_in_r_bypass_27_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_1_stall_19 <= io_in_r_bypass_27_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_2_data_19 <= io_in_r_bypass_27_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_2_load_store_19 <= io_in_r_bypass_27_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_2_df_is_ws_19 <= io_in_r_bypass_27_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_2_stall_19 <= io_in_r_bypass_27_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_3_data_19 <= io_in_r_bypass_27_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_3_load_store_19 <= io_in_r_bypass_27_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_3_df_is_ws_19 <= io_in_r_bypass_27_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_3_stall_19 <= io_in_r_bypass_27_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_0_data_19 <= io_in_r_bypass_28_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_0_load_store_19 <= io_in_r_bypass_28_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_0_df_is_ws_19 <= io_in_r_bypass_28_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_0_stall_19 <= io_in_r_bypass_28_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_1_data_19 <= io_in_r_bypass_28_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_1_load_store_19 <= io_in_r_bypass_28_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_1_df_is_ws_19 <= io_in_r_bypass_28_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_1_stall_19 <= io_in_r_bypass_28_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_2_data_19 <= io_in_r_bypass_28_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_2_load_store_19 <= io_in_r_bypass_28_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_2_df_is_ws_19 <= io_in_r_bypass_28_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_2_stall_19 <= io_in_r_bypass_28_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_3_data_19 <= io_in_r_bypass_28_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_3_load_store_19 <= io_in_r_bypass_28_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_3_df_is_ws_19 <= io_in_r_bypass_28_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_3_stall_19 <= io_in_r_bypass_28_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_0_data_19 <= io_in_r_bypass_29_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_0_load_store_19 <= io_in_r_bypass_29_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_0_df_is_ws_19 <= io_in_r_bypass_29_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_0_stall_19 <= io_in_r_bypass_29_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_1_data_19 <= io_in_r_bypass_29_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_1_load_store_19 <= io_in_r_bypass_29_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_1_df_is_ws_19 <= io_in_r_bypass_29_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_1_stall_19 <= io_in_r_bypass_29_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_2_data_19 <= io_in_r_bypass_29_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_2_load_store_19 <= io_in_r_bypass_29_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_2_df_is_ws_19 <= io_in_r_bypass_29_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_2_stall_19 <= io_in_r_bypass_29_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_3_data_19 <= io_in_r_bypass_29_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_3_load_store_19 <= io_in_r_bypass_29_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_3_df_is_ws_19 <= io_in_r_bypass_29_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_3_stall_19 <= io_in_r_bypass_29_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_0_data_19 <= io_in_r_bypass_30_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_0_load_store_19 <= io_in_r_bypass_30_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_0_df_is_ws_19 <= io_in_r_bypass_30_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_0_stall_19 <= io_in_r_bypass_30_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_1_data_19 <= io_in_r_bypass_30_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_1_load_store_19 <= io_in_r_bypass_30_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_1_df_is_ws_19 <= io_in_r_bypass_30_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_1_stall_19 <= io_in_r_bypass_30_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_2_data_19 <= io_in_r_bypass_30_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_2_load_store_19 <= io_in_r_bypass_30_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_2_df_is_ws_19 <= io_in_r_bypass_30_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_2_stall_19 <= io_in_r_bypass_30_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_3_data_19 <= io_in_r_bypass_30_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_3_load_store_19 <= io_in_r_bypass_30_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_3_df_is_ws_19 <= io_in_r_bypass_30_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_3_stall_19 <= io_in_r_bypass_30_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_0_data_19 <= io_in_r_bypass_31_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_0_load_store_19 <= io_in_r_bypass_31_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_0_df_is_ws_19 <= io_in_r_bypass_31_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_0_stall_19 <= io_in_r_bypass_31_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_1_data_19 <= io_in_r_bypass_31_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_1_load_store_19 <= io_in_r_bypass_31_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_1_df_is_ws_19 <= io_in_r_bypass_31_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_1_stall_19 <= io_in_r_bypass_31_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_2_data_19 <= io_in_r_bypass_31_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_2_load_store_19 <= io_in_r_bypass_31_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_2_df_is_ws_19 <= io_in_r_bypass_31_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_2_stall_19 <= io_in_r_bypass_31_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_3_data_19 <= io_in_r_bypass_31_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_3_load_store_19 <= io_in_r_bypass_31_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_3_df_is_ws_19 <= io_in_r_bypass_31_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_3_stall_19 <= io_in_r_bypass_31_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_0_data_20 <= io_in_r_bypass_0_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_0_load_store_20 <= io_in_r_bypass_0_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_0_df_is_ws_20 <= io_in_r_bypass_0_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_0_stall_20 <= io_in_r_bypass_0_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_1_data_20 <= io_in_r_bypass_0_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_1_load_store_20 <= io_in_r_bypass_0_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_1_df_is_ws_20 <= io_in_r_bypass_0_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_1_stall_20 <= io_in_r_bypass_0_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_2_data_20 <= io_in_r_bypass_0_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_2_load_store_20 <= io_in_r_bypass_0_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_2_df_is_ws_20 <= io_in_r_bypass_0_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_2_stall_20 <= io_in_r_bypass_0_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_3_data_20 <= io_in_r_bypass_0_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_3_load_store_20 <= io_in_r_bypass_0_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_3_df_is_ws_20 <= io_in_r_bypass_0_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_3_stall_20 <= io_in_r_bypass_0_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_0_data_20 <= io_in_r_bypass_1_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_0_load_store_20 <= io_in_r_bypass_1_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_0_df_is_ws_20 <= io_in_r_bypass_1_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_0_stall_20 <= io_in_r_bypass_1_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_1_data_20 <= io_in_r_bypass_1_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_1_load_store_20 <= io_in_r_bypass_1_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_1_df_is_ws_20 <= io_in_r_bypass_1_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_1_stall_20 <= io_in_r_bypass_1_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_2_data_20 <= io_in_r_bypass_1_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_2_load_store_20 <= io_in_r_bypass_1_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_2_df_is_ws_20 <= io_in_r_bypass_1_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_2_stall_20 <= io_in_r_bypass_1_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_3_data_20 <= io_in_r_bypass_1_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_3_load_store_20 <= io_in_r_bypass_1_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_3_df_is_ws_20 <= io_in_r_bypass_1_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_3_stall_20 <= io_in_r_bypass_1_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_0_data_20 <= io_in_r_bypass_2_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_0_load_store_20 <= io_in_r_bypass_2_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_0_df_is_ws_20 <= io_in_r_bypass_2_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_0_stall_20 <= io_in_r_bypass_2_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_1_data_20 <= io_in_r_bypass_2_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_1_load_store_20 <= io_in_r_bypass_2_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_1_df_is_ws_20 <= io_in_r_bypass_2_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_1_stall_20 <= io_in_r_bypass_2_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_2_data_20 <= io_in_r_bypass_2_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_2_load_store_20 <= io_in_r_bypass_2_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_2_df_is_ws_20 <= io_in_r_bypass_2_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_2_stall_20 <= io_in_r_bypass_2_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_3_data_20 <= io_in_r_bypass_2_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_3_load_store_20 <= io_in_r_bypass_2_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_3_df_is_ws_20 <= io_in_r_bypass_2_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_3_stall_20 <= io_in_r_bypass_2_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_0_data_20 <= io_in_r_bypass_3_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_0_load_store_20 <= io_in_r_bypass_3_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_0_df_is_ws_20 <= io_in_r_bypass_3_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_0_stall_20 <= io_in_r_bypass_3_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_1_data_20 <= io_in_r_bypass_3_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_1_load_store_20 <= io_in_r_bypass_3_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_1_df_is_ws_20 <= io_in_r_bypass_3_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_1_stall_20 <= io_in_r_bypass_3_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_2_data_20 <= io_in_r_bypass_3_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_2_load_store_20 <= io_in_r_bypass_3_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_2_df_is_ws_20 <= io_in_r_bypass_3_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_2_stall_20 <= io_in_r_bypass_3_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_3_data_20 <= io_in_r_bypass_3_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_3_load_store_20 <= io_in_r_bypass_3_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_3_df_is_ws_20 <= io_in_r_bypass_3_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_3_stall_20 <= io_in_r_bypass_3_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_0_data_20 <= io_in_r_bypass_4_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_0_load_store_20 <= io_in_r_bypass_4_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_0_df_is_ws_20 <= io_in_r_bypass_4_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_0_stall_20 <= io_in_r_bypass_4_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_1_data_20 <= io_in_r_bypass_4_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_1_load_store_20 <= io_in_r_bypass_4_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_1_df_is_ws_20 <= io_in_r_bypass_4_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_1_stall_20 <= io_in_r_bypass_4_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_2_data_20 <= io_in_r_bypass_4_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_2_load_store_20 <= io_in_r_bypass_4_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_2_df_is_ws_20 <= io_in_r_bypass_4_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_2_stall_20 <= io_in_r_bypass_4_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_3_data_20 <= io_in_r_bypass_4_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_3_load_store_20 <= io_in_r_bypass_4_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_3_df_is_ws_20 <= io_in_r_bypass_4_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_3_stall_20 <= io_in_r_bypass_4_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_0_data_20 <= io_in_r_bypass_5_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_0_load_store_20 <= io_in_r_bypass_5_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_0_df_is_ws_20 <= io_in_r_bypass_5_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_0_stall_20 <= io_in_r_bypass_5_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_1_data_20 <= io_in_r_bypass_5_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_1_load_store_20 <= io_in_r_bypass_5_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_1_df_is_ws_20 <= io_in_r_bypass_5_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_1_stall_20 <= io_in_r_bypass_5_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_2_data_20 <= io_in_r_bypass_5_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_2_load_store_20 <= io_in_r_bypass_5_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_2_df_is_ws_20 <= io_in_r_bypass_5_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_2_stall_20 <= io_in_r_bypass_5_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_3_data_20 <= io_in_r_bypass_5_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_3_load_store_20 <= io_in_r_bypass_5_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_3_df_is_ws_20 <= io_in_r_bypass_5_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_3_stall_20 <= io_in_r_bypass_5_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_0_data_20 <= io_in_r_bypass_6_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_0_load_store_20 <= io_in_r_bypass_6_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_0_df_is_ws_20 <= io_in_r_bypass_6_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_0_stall_20 <= io_in_r_bypass_6_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_1_data_20 <= io_in_r_bypass_6_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_1_load_store_20 <= io_in_r_bypass_6_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_1_df_is_ws_20 <= io_in_r_bypass_6_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_1_stall_20 <= io_in_r_bypass_6_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_2_data_20 <= io_in_r_bypass_6_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_2_load_store_20 <= io_in_r_bypass_6_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_2_df_is_ws_20 <= io_in_r_bypass_6_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_2_stall_20 <= io_in_r_bypass_6_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_3_data_20 <= io_in_r_bypass_6_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_3_load_store_20 <= io_in_r_bypass_6_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_3_df_is_ws_20 <= io_in_r_bypass_6_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_3_stall_20 <= io_in_r_bypass_6_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_0_data_20 <= io_in_r_bypass_7_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_0_load_store_20 <= io_in_r_bypass_7_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_0_df_is_ws_20 <= io_in_r_bypass_7_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_0_stall_20 <= io_in_r_bypass_7_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_1_data_20 <= io_in_r_bypass_7_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_1_load_store_20 <= io_in_r_bypass_7_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_1_df_is_ws_20 <= io_in_r_bypass_7_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_1_stall_20 <= io_in_r_bypass_7_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_2_data_20 <= io_in_r_bypass_7_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_2_load_store_20 <= io_in_r_bypass_7_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_2_df_is_ws_20 <= io_in_r_bypass_7_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_2_stall_20 <= io_in_r_bypass_7_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_3_data_20 <= io_in_r_bypass_7_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_3_load_store_20 <= io_in_r_bypass_7_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_3_df_is_ws_20 <= io_in_r_bypass_7_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_3_stall_20 <= io_in_r_bypass_7_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_0_data_20 <= io_in_r_bypass_8_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_0_load_store_20 <= io_in_r_bypass_8_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_0_df_is_ws_20 <= io_in_r_bypass_8_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_0_stall_20 <= io_in_r_bypass_8_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_1_data_20 <= io_in_r_bypass_8_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_1_load_store_20 <= io_in_r_bypass_8_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_1_df_is_ws_20 <= io_in_r_bypass_8_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_1_stall_20 <= io_in_r_bypass_8_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_2_data_20 <= io_in_r_bypass_8_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_2_load_store_20 <= io_in_r_bypass_8_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_2_df_is_ws_20 <= io_in_r_bypass_8_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_2_stall_20 <= io_in_r_bypass_8_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_3_data_20 <= io_in_r_bypass_8_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_3_load_store_20 <= io_in_r_bypass_8_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_3_df_is_ws_20 <= io_in_r_bypass_8_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_3_stall_20 <= io_in_r_bypass_8_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_0_data_20 <= io_in_r_bypass_9_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_0_load_store_20 <= io_in_r_bypass_9_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_0_df_is_ws_20 <= io_in_r_bypass_9_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_0_stall_20 <= io_in_r_bypass_9_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_1_data_20 <= io_in_r_bypass_9_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_1_load_store_20 <= io_in_r_bypass_9_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_1_df_is_ws_20 <= io_in_r_bypass_9_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_1_stall_20 <= io_in_r_bypass_9_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_2_data_20 <= io_in_r_bypass_9_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_2_load_store_20 <= io_in_r_bypass_9_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_2_df_is_ws_20 <= io_in_r_bypass_9_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_2_stall_20 <= io_in_r_bypass_9_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_3_data_20 <= io_in_r_bypass_9_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_3_load_store_20 <= io_in_r_bypass_9_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_3_df_is_ws_20 <= io_in_r_bypass_9_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_3_stall_20 <= io_in_r_bypass_9_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_0_data_20 <= io_in_r_bypass_10_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_0_load_store_20 <= io_in_r_bypass_10_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_0_df_is_ws_20 <= io_in_r_bypass_10_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_0_stall_20 <= io_in_r_bypass_10_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_1_data_20 <= io_in_r_bypass_10_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_1_load_store_20 <= io_in_r_bypass_10_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_1_df_is_ws_20 <= io_in_r_bypass_10_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_1_stall_20 <= io_in_r_bypass_10_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_2_data_20 <= io_in_r_bypass_10_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_2_load_store_20 <= io_in_r_bypass_10_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_2_df_is_ws_20 <= io_in_r_bypass_10_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_2_stall_20 <= io_in_r_bypass_10_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_3_data_20 <= io_in_r_bypass_10_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_3_load_store_20 <= io_in_r_bypass_10_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_3_df_is_ws_20 <= io_in_r_bypass_10_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_3_stall_20 <= io_in_r_bypass_10_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_0_data_20 <= io_in_r_bypass_11_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_0_load_store_20 <= io_in_r_bypass_11_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_0_df_is_ws_20 <= io_in_r_bypass_11_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_0_stall_20 <= io_in_r_bypass_11_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_1_data_20 <= io_in_r_bypass_11_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_1_load_store_20 <= io_in_r_bypass_11_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_1_df_is_ws_20 <= io_in_r_bypass_11_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_1_stall_20 <= io_in_r_bypass_11_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_2_data_20 <= io_in_r_bypass_11_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_2_load_store_20 <= io_in_r_bypass_11_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_2_df_is_ws_20 <= io_in_r_bypass_11_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_2_stall_20 <= io_in_r_bypass_11_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_3_data_20 <= io_in_r_bypass_11_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_3_load_store_20 <= io_in_r_bypass_11_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_3_df_is_ws_20 <= io_in_r_bypass_11_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_3_stall_20 <= io_in_r_bypass_11_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_0_data_20 <= io_in_r_bypass_12_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_0_load_store_20 <= io_in_r_bypass_12_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_0_df_is_ws_20 <= io_in_r_bypass_12_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_0_stall_20 <= io_in_r_bypass_12_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_1_data_20 <= io_in_r_bypass_12_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_1_load_store_20 <= io_in_r_bypass_12_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_1_df_is_ws_20 <= io_in_r_bypass_12_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_1_stall_20 <= io_in_r_bypass_12_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_2_data_20 <= io_in_r_bypass_12_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_2_load_store_20 <= io_in_r_bypass_12_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_2_df_is_ws_20 <= io_in_r_bypass_12_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_2_stall_20 <= io_in_r_bypass_12_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_3_data_20 <= io_in_r_bypass_12_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_3_load_store_20 <= io_in_r_bypass_12_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_3_df_is_ws_20 <= io_in_r_bypass_12_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_3_stall_20 <= io_in_r_bypass_12_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_0_data_20 <= io_in_r_bypass_13_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_0_load_store_20 <= io_in_r_bypass_13_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_0_df_is_ws_20 <= io_in_r_bypass_13_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_0_stall_20 <= io_in_r_bypass_13_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_1_data_20 <= io_in_r_bypass_13_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_1_load_store_20 <= io_in_r_bypass_13_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_1_df_is_ws_20 <= io_in_r_bypass_13_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_1_stall_20 <= io_in_r_bypass_13_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_2_data_20 <= io_in_r_bypass_13_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_2_load_store_20 <= io_in_r_bypass_13_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_2_df_is_ws_20 <= io_in_r_bypass_13_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_2_stall_20 <= io_in_r_bypass_13_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_3_data_20 <= io_in_r_bypass_13_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_3_load_store_20 <= io_in_r_bypass_13_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_3_df_is_ws_20 <= io_in_r_bypass_13_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_3_stall_20 <= io_in_r_bypass_13_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_0_data_20 <= io_in_r_bypass_14_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_0_load_store_20 <= io_in_r_bypass_14_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_0_df_is_ws_20 <= io_in_r_bypass_14_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_0_stall_20 <= io_in_r_bypass_14_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_1_data_20 <= io_in_r_bypass_14_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_1_load_store_20 <= io_in_r_bypass_14_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_1_df_is_ws_20 <= io_in_r_bypass_14_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_1_stall_20 <= io_in_r_bypass_14_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_2_data_20 <= io_in_r_bypass_14_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_2_load_store_20 <= io_in_r_bypass_14_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_2_df_is_ws_20 <= io_in_r_bypass_14_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_2_stall_20 <= io_in_r_bypass_14_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_3_data_20 <= io_in_r_bypass_14_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_3_load_store_20 <= io_in_r_bypass_14_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_3_df_is_ws_20 <= io_in_r_bypass_14_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_3_stall_20 <= io_in_r_bypass_14_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_0_data_20 <= io_in_r_bypass_15_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_0_load_store_20 <= io_in_r_bypass_15_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_0_df_is_ws_20 <= io_in_r_bypass_15_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_0_stall_20 <= io_in_r_bypass_15_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_1_data_20 <= io_in_r_bypass_15_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_1_load_store_20 <= io_in_r_bypass_15_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_1_df_is_ws_20 <= io_in_r_bypass_15_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_1_stall_20 <= io_in_r_bypass_15_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_2_data_20 <= io_in_r_bypass_15_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_2_load_store_20 <= io_in_r_bypass_15_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_2_df_is_ws_20 <= io_in_r_bypass_15_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_2_stall_20 <= io_in_r_bypass_15_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_3_data_20 <= io_in_r_bypass_15_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_3_load_store_20 <= io_in_r_bypass_15_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_3_df_is_ws_20 <= io_in_r_bypass_15_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_3_stall_20 <= io_in_r_bypass_15_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_0_data_20 <= io_in_r_bypass_16_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_0_load_store_20 <= io_in_r_bypass_16_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_0_df_is_ws_20 <= io_in_r_bypass_16_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_0_stall_20 <= io_in_r_bypass_16_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_1_data_20 <= io_in_r_bypass_16_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_1_load_store_20 <= io_in_r_bypass_16_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_1_df_is_ws_20 <= io_in_r_bypass_16_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_1_stall_20 <= io_in_r_bypass_16_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_2_data_20 <= io_in_r_bypass_16_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_2_load_store_20 <= io_in_r_bypass_16_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_2_df_is_ws_20 <= io_in_r_bypass_16_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_2_stall_20 <= io_in_r_bypass_16_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_3_data_20 <= io_in_r_bypass_16_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_3_load_store_20 <= io_in_r_bypass_16_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_3_df_is_ws_20 <= io_in_r_bypass_16_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_3_stall_20 <= io_in_r_bypass_16_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_0_data_20 <= io_in_r_bypass_17_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_0_load_store_20 <= io_in_r_bypass_17_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_0_df_is_ws_20 <= io_in_r_bypass_17_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_0_stall_20 <= io_in_r_bypass_17_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_1_data_20 <= io_in_r_bypass_17_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_1_load_store_20 <= io_in_r_bypass_17_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_1_df_is_ws_20 <= io_in_r_bypass_17_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_1_stall_20 <= io_in_r_bypass_17_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_2_data_20 <= io_in_r_bypass_17_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_2_load_store_20 <= io_in_r_bypass_17_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_2_df_is_ws_20 <= io_in_r_bypass_17_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_2_stall_20 <= io_in_r_bypass_17_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_3_data_20 <= io_in_r_bypass_17_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_3_load_store_20 <= io_in_r_bypass_17_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_3_df_is_ws_20 <= io_in_r_bypass_17_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_3_stall_20 <= io_in_r_bypass_17_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_0_data_20 <= io_in_r_bypass_18_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_0_load_store_20 <= io_in_r_bypass_18_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_0_df_is_ws_20 <= io_in_r_bypass_18_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_0_stall_20 <= io_in_r_bypass_18_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_1_data_20 <= io_in_r_bypass_18_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_1_load_store_20 <= io_in_r_bypass_18_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_1_df_is_ws_20 <= io_in_r_bypass_18_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_1_stall_20 <= io_in_r_bypass_18_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_2_data_20 <= io_in_r_bypass_18_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_2_load_store_20 <= io_in_r_bypass_18_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_2_df_is_ws_20 <= io_in_r_bypass_18_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_2_stall_20 <= io_in_r_bypass_18_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_3_data_20 <= io_in_r_bypass_18_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_3_load_store_20 <= io_in_r_bypass_18_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_3_df_is_ws_20 <= io_in_r_bypass_18_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_3_stall_20 <= io_in_r_bypass_18_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_0_data_20 <= io_in_r_bypass_19_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_0_load_store_20 <= io_in_r_bypass_19_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_0_df_is_ws_20 <= io_in_r_bypass_19_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_0_stall_20 <= io_in_r_bypass_19_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_1_data_20 <= io_in_r_bypass_19_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_1_load_store_20 <= io_in_r_bypass_19_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_1_df_is_ws_20 <= io_in_r_bypass_19_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_1_stall_20 <= io_in_r_bypass_19_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_2_data_20 <= io_in_r_bypass_19_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_2_load_store_20 <= io_in_r_bypass_19_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_2_df_is_ws_20 <= io_in_r_bypass_19_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_2_stall_20 <= io_in_r_bypass_19_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_3_data_20 <= io_in_r_bypass_19_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_3_load_store_20 <= io_in_r_bypass_19_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_3_df_is_ws_20 <= io_in_r_bypass_19_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_3_stall_20 <= io_in_r_bypass_19_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_0_data_20 <= io_in_r_bypass_20_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_0_load_store_20 <= io_in_r_bypass_20_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_0_df_is_ws_20 <= io_in_r_bypass_20_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_0_stall_20 <= io_in_r_bypass_20_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_1_data_20 <= io_in_r_bypass_20_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_1_load_store_20 <= io_in_r_bypass_20_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_1_df_is_ws_20 <= io_in_r_bypass_20_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_1_stall_20 <= io_in_r_bypass_20_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_2_data_20 <= io_in_r_bypass_20_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_2_load_store_20 <= io_in_r_bypass_20_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_2_df_is_ws_20 <= io_in_r_bypass_20_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_2_stall_20 <= io_in_r_bypass_20_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_3_data_20 <= io_in_r_bypass_20_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_3_load_store_20 <= io_in_r_bypass_20_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_3_df_is_ws_20 <= io_in_r_bypass_20_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_3_stall_20 <= io_in_r_bypass_20_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_0_data_20 <= io_in_r_bypass_21_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_0_load_store_20 <= io_in_r_bypass_21_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_0_df_is_ws_20 <= io_in_r_bypass_21_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_0_stall_20 <= io_in_r_bypass_21_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_1_data_20 <= io_in_r_bypass_21_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_1_load_store_20 <= io_in_r_bypass_21_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_1_df_is_ws_20 <= io_in_r_bypass_21_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_1_stall_20 <= io_in_r_bypass_21_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_2_data_20 <= io_in_r_bypass_21_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_2_load_store_20 <= io_in_r_bypass_21_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_2_df_is_ws_20 <= io_in_r_bypass_21_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_2_stall_20 <= io_in_r_bypass_21_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_3_data_20 <= io_in_r_bypass_21_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_3_load_store_20 <= io_in_r_bypass_21_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_3_df_is_ws_20 <= io_in_r_bypass_21_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_3_stall_20 <= io_in_r_bypass_21_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_0_data_20 <= io_in_r_bypass_22_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_0_load_store_20 <= io_in_r_bypass_22_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_0_df_is_ws_20 <= io_in_r_bypass_22_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_0_stall_20 <= io_in_r_bypass_22_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_1_data_20 <= io_in_r_bypass_22_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_1_load_store_20 <= io_in_r_bypass_22_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_1_df_is_ws_20 <= io_in_r_bypass_22_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_1_stall_20 <= io_in_r_bypass_22_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_2_data_20 <= io_in_r_bypass_22_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_2_load_store_20 <= io_in_r_bypass_22_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_2_df_is_ws_20 <= io_in_r_bypass_22_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_2_stall_20 <= io_in_r_bypass_22_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_3_data_20 <= io_in_r_bypass_22_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_3_load_store_20 <= io_in_r_bypass_22_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_3_df_is_ws_20 <= io_in_r_bypass_22_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_3_stall_20 <= io_in_r_bypass_22_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_0_data_20 <= io_in_r_bypass_23_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_0_load_store_20 <= io_in_r_bypass_23_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_0_df_is_ws_20 <= io_in_r_bypass_23_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_0_stall_20 <= io_in_r_bypass_23_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_1_data_20 <= io_in_r_bypass_23_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_1_load_store_20 <= io_in_r_bypass_23_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_1_df_is_ws_20 <= io_in_r_bypass_23_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_1_stall_20 <= io_in_r_bypass_23_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_2_data_20 <= io_in_r_bypass_23_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_2_load_store_20 <= io_in_r_bypass_23_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_2_df_is_ws_20 <= io_in_r_bypass_23_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_2_stall_20 <= io_in_r_bypass_23_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_3_data_20 <= io_in_r_bypass_23_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_3_load_store_20 <= io_in_r_bypass_23_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_3_df_is_ws_20 <= io_in_r_bypass_23_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_3_stall_20 <= io_in_r_bypass_23_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_0_data_20 <= io_in_r_bypass_24_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_0_load_store_20 <= io_in_r_bypass_24_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_0_df_is_ws_20 <= io_in_r_bypass_24_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_0_stall_20 <= io_in_r_bypass_24_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_1_data_20 <= io_in_r_bypass_24_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_1_load_store_20 <= io_in_r_bypass_24_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_1_df_is_ws_20 <= io_in_r_bypass_24_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_1_stall_20 <= io_in_r_bypass_24_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_2_data_20 <= io_in_r_bypass_24_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_2_load_store_20 <= io_in_r_bypass_24_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_2_df_is_ws_20 <= io_in_r_bypass_24_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_2_stall_20 <= io_in_r_bypass_24_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_3_data_20 <= io_in_r_bypass_24_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_3_load_store_20 <= io_in_r_bypass_24_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_3_df_is_ws_20 <= io_in_r_bypass_24_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_3_stall_20 <= io_in_r_bypass_24_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_0_data_20 <= io_in_r_bypass_25_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_0_load_store_20 <= io_in_r_bypass_25_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_0_df_is_ws_20 <= io_in_r_bypass_25_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_0_stall_20 <= io_in_r_bypass_25_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_1_data_20 <= io_in_r_bypass_25_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_1_load_store_20 <= io_in_r_bypass_25_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_1_df_is_ws_20 <= io_in_r_bypass_25_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_1_stall_20 <= io_in_r_bypass_25_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_2_data_20 <= io_in_r_bypass_25_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_2_load_store_20 <= io_in_r_bypass_25_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_2_df_is_ws_20 <= io_in_r_bypass_25_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_2_stall_20 <= io_in_r_bypass_25_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_3_data_20 <= io_in_r_bypass_25_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_3_load_store_20 <= io_in_r_bypass_25_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_3_df_is_ws_20 <= io_in_r_bypass_25_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_3_stall_20 <= io_in_r_bypass_25_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_0_data_20 <= io_in_r_bypass_26_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_0_load_store_20 <= io_in_r_bypass_26_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_0_df_is_ws_20 <= io_in_r_bypass_26_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_0_stall_20 <= io_in_r_bypass_26_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_1_data_20 <= io_in_r_bypass_26_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_1_load_store_20 <= io_in_r_bypass_26_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_1_df_is_ws_20 <= io_in_r_bypass_26_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_1_stall_20 <= io_in_r_bypass_26_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_2_data_20 <= io_in_r_bypass_26_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_2_load_store_20 <= io_in_r_bypass_26_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_2_df_is_ws_20 <= io_in_r_bypass_26_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_2_stall_20 <= io_in_r_bypass_26_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_3_data_20 <= io_in_r_bypass_26_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_3_load_store_20 <= io_in_r_bypass_26_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_3_df_is_ws_20 <= io_in_r_bypass_26_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_3_stall_20 <= io_in_r_bypass_26_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_0_data_20 <= io_in_r_bypass_27_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_0_load_store_20 <= io_in_r_bypass_27_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_0_df_is_ws_20 <= io_in_r_bypass_27_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_0_stall_20 <= io_in_r_bypass_27_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_1_data_20 <= io_in_r_bypass_27_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_1_load_store_20 <= io_in_r_bypass_27_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_1_df_is_ws_20 <= io_in_r_bypass_27_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_1_stall_20 <= io_in_r_bypass_27_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_2_data_20 <= io_in_r_bypass_27_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_2_load_store_20 <= io_in_r_bypass_27_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_2_df_is_ws_20 <= io_in_r_bypass_27_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_2_stall_20 <= io_in_r_bypass_27_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_3_data_20 <= io_in_r_bypass_27_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_3_load_store_20 <= io_in_r_bypass_27_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_3_df_is_ws_20 <= io_in_r_bypass_27_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_3_stall_20 <= io_in_r_bypass_27_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_0_data_20 <= io_in_r_bypass_28_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_0_load_store_20 <= io_in_r_bypass_28_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_0_df_is_ws_20 <= io_in_r_bypass_28_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_0_stall_20 <= io_in_r_bypass_28_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_1_data_20 <= io_in_r_bypass_28_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_1_load_store_20 <= io_in_r_bypass_28_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_1_df_is_ws_20 <= io_in_r_bypass_28_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_1_stall_20 <= io_in_r_bypass_28_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_2_data_20 <= io_in_r_bypass_28_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_2_load_store_20 <= io_in_r_bypass_28_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_2_df_is_ws_20 <= io_in_r_bypass_28_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_2_stall_20 <= io_in_r_bypass_28_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_3_data_20 <= io_in_r_bypass_28_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_3_load_store_20 <= io_in_r_bypass_28_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_3_df_is_ws_20 <= io_in_r_bypass_28_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_3_stall_20 <= io_in_r_bypass_28_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_0_data_20 <= io_in_r_bypass_29_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_0_load_store_20 <= io_in_r_bypass_29_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_0_df_is_ws_20 <= io_in_r_bypass_29_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_0_stall_20 <= io_in_r_bypass_29_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_1_data_20 <= io_in_r_bypass_29_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_1_load_store_20 <= io_in_r_bypass_29_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_1_df_is_ws_20 <= io_in_r_bypass_29_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_1_stall_20 <= io_in_r_bypass_29_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_2_data_20 <= io_in_r_bypass_29_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_2_load_store_20 <= io_in_r_bypass_29_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_2_df_is_ws_20 <= io_in_r_bypass_29_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_2_stall_20 <= io_in_r_bypass_29_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_3_data_20 <= io_in_r_bypass_29_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_3_load_store_20 <= io_in_r_bypass_29_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_3_df_is_ws_20 <= io_in_r_bypass_29_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_3_stall_20 <= io_in_r_bypass_29_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_0_data_20 <= io_in_r_bypass_30_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_0_load_store_20 <= io_in_r_bypass_30_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_0_df_is_ws_20 <= io_in_r_bypass_30_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_0_stall_20 <= io_in_r_bypass_30_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_1_data_20 <= io_in_r_bypass_30_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_1_load_store_20 <= io_in_r_bypass_30_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_1_df_is_ws_20 <= io_in_r_bypass_30_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_1_stall_20 <= io_in_r_bypass_30_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_2_data_20 <= io_in_r_bypass_30_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_2_load_store_20 <= io_in_r_bypass_30_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_2_df_is_ws_20 <= io_in_r_bypass_30_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_2_stall_20 <= io_in_r_bypass_30_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_3_data_20 <= io_in_r_bypass_30_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_3_load_store_20 <= io_in_r_bypass_30_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_3_df_is_ws_20 <= io_in_r_bypass_30_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_3_stall_20 <= io_in_r_bypass_30_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_0_data_20 <= io_in_r_bypass_31_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_0_load_store_20 <= io_in_r_bypass_31_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_0_df_is_ws_20 <= io_in_r_bypass_31_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_0_stall_20 <= io_in_r_bypass_31_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_1_data_20 <= io_in_r_bypass_31_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_1_load_store_20 <= io_in_r_bypass_31_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_1_df_is_ws_20 <= io_in_r_bypass_31_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_1_stall_20 <= io_in_r_bypass_31_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_2_data_20 <= io_in_r_bypass_31_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_2_load_store_20 <= io_in_r_bypass_31_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_2_df_is_ws_20 <= io_in_r_bypass_31_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_2_stall_20 <= io_in_r_bypass_31_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_3_data_20 <= io_in_r_bypass_31_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_3_load_store_20 <= io_in_r_bypass_31_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_3_df_is_ws_20 <= io_in_r_bypass_31_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_3_stall_20 <= io_in_r_bypass_31_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_0_data_21 <= io_in_r_bypass_0_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_0_load_store_21 <= io_in_r_bypass_0_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_0_df_is_ws_21 <= io_in_r_bypass_0_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_0_stall_21 <= io_in_r_bypass_0_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_1_data_21 <= io_in_r_bypass_0_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_1_load_store_21 <= io_in_r_bypass_0_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_1_df_is_ws_21 <= io_in_r_bypass_0_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_1_stall_21 <= io_in_r_bypass_0_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_2_data_21 <= io_in_r_bypass_0_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_2_load_store_21 <= io_in_r_bypass_0_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_2_df_is_ws_21 <= io_in_r_bypass_0_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_2_stall_21 <= io_in_r_bypass_0_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_3_data_21 <= io_in_r_bypass_0_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_3_load_store_21 <= io_in_r_bypass_0_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_3_df_is_ws_21 <= io_in_r_bypass_0_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_3_stall_21 <= io_in_r_bypass_0_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_0_data_21 <= io_in_r_bypass_1_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_0_load_store_21 <= io_in_r_bypass_1_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_0_df_is_ws_21 <= io_in_r_bypass_1_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_0_stall_21 <= io_in_r_bypass_1_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_1_data_21 <= io_in_r_bypass_1_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_1_load_store_21 <= io_in_r_bypass_1_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_1_df_is_ws_21 <= io_in_r_bypass_1_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_1_stall_21 <= io_in_r_bypass_1_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_2_data_21 <= io_in_r_bypass_1_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_2_load_store_21 <= io_in_r_bypass_1_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_2_df_is_ws_21 <= io_in_r_bypass_1_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_2_stall_21 <= io_in_r_bypass_1_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_3_data_21 <= io_in_r_bypass_1_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_3_load_store_21 <= io_in_r_bypass_1_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_3_df_is_ws_21 <= io_in_r_bypass_1_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_3_stall_21 <= io_in_r_bypass_1_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_0_data_21 <= io_in_r_bypass_2_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_0_load_store_21 <= io_in_r_bypass_2_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_0_df_is_ws_21 <= io_in_r_bypass_2_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_0_stall_21 <= io_in_r_bypass_2_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_1_data_21 <= io_in_r_bypass_2_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_1_load_store_21 <= io_in_r_bypass_2_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_1_df_is_ws_21 <= io_in_r_bypass_2_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_1_stall_21 <= io_in_r_bypass_2_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_2_data_21 <= io_in_r_bypass_2_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_2_load_store_21 <= io_in_r_bypass_2_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_2_df_is_ws_21 <= io_in_r_bypass_2_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_2_stall_21 <= io_in_r_bypass_2_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_3_data_21 <= io_in_r_bypass_2_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_3_load_store_21 <= io_in_r_bypass_2_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_3_df_is_ws_21 <= io_in_r_bypass_2_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_3_stall_21 <= io_in_r_bypass_2_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_0_data_21 <= io_in_r_bypass_3_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_0_load_store_21 <= io_in_r_bypass_3_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_0_df_is_ws_21 <= io_in_r_bypass_3_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_0_stall_21 <= io_in_r_bypass_3_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_1_data_21 <= io_in_r_bypass_3_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_1_load_store_21 <= io_in_r_bypass_3_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_1_df_is_ws_21 <= io_in_r_bypass_3_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_1_stall_21 <= io_in_r_bypass_3_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_2_data_21 <= io_in_r_bypass_3_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_2_load_store_21 <= io_in_r_bypass_3_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_2_df_is_ws_21 <= io_in_r_bypass_3_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_2_stall_21 <= io_in_r_bypass_3_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_3_data_21 <= io_in_r_bypass_3_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_3_load_store_21 <= io_in_r_bypass_3_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_3_df_is_ws_21 <= io_in_r_bypass_3_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_3_stall_21 <= io_in_r_bypass_3_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_0_data_21 <= io_in_r_bypass_4_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_0_load_store_21 <= io_in_r_bypass_4_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_0_df_is_ws_21 <= io_in_r_bypass_4_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_0_stall_21 <= io_in_r_bypass_4_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_1_data_21 <= io_in_r_bypass_4_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_1_load_store_21 <= io_in_r_bypass_4_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_1_df_is_ws_21 <= io_in_r_bypass_4_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_1_stall_21 <= io_in_r_bypass_4_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_2_data_21 <= io_in_r_bypass_4_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_2_load_store_21 <= io_in_r_bypass_4_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_2_df_is_ws_21 <= io_in_r_bypass_4_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_2_stall_21 <= io_in_r_bypass_4_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_3_data_21 <= io_in_r_bypass_4_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_3_load_store_21 <= io_in_r_bypass_4_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_3_df_is_ws_21 <= io_in_r_bypass_4_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_3_stall_21 <= io_in_r_bypass_4_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_0_data_21 <= io_in_r_bypass_5_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_0_load_store_21 <= io_in_r_bypass_5_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_0_df_is_ws_21 <= io_in_r_bypass_5_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_0_stall_21 <= io_in_r_bypass_5_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_1_data_21 <= io_in_r_bypass_5_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_1_load_store_21 <= io_in_r_bypass_5_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_1_df_is_ws_21 <= io_in_r_bypass_5_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_1_stall_21 <= io_in_r_bypass_5_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_2_data_21 <= io_in_r_bypass_5_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_2_load_store_21 <= io_in_r_bypass_5_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_2_df_is_ws_21 <= io_in_r_bypass_5_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_2_stall_21 <= io_in_r_bypass_5_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_3_data_21 <= io_in_r_bypass_5_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_3_load_store_21 <= io_in_r_bypass_5_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_3_df_is_ws_21 <= io_in_r_bypass_5_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_3_stall_21 <= io_in_r_bypass_5_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_0_data_21 <= io_in_r_bypass_6_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_0_load_store_21 <= io_in_r_bypass_6_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_0_df_is_ws_21 <= io_in_r_bypass_6_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_0_stall_21 <= io_in_r_bypass_6_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_1_data_21 <= io_in_r_bypass_6_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_1_load_store_21 <= io_in_r_bypass_6_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_1_df_is_ws_21 <= io_in_r_bypass_6_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_1_stall_21 <= io_in_r_bypass_6_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_2_data_21 <= io_in_r_bypass_6_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_2_load_store_21 <= io_in_r_bypass_6_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_2_df_is_ws_21 <= io_in_r_bypass_6_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_2_stall_21 <= io_in_r_bypass_6_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_3_data_21 <= io_in_r_bypass_6_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_3_load_store_21 <= io_in_r_bypass_6_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_3_df_is_ws_21 <= io_in_r_bypass_6_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_3_stall_21 <= io_in_r_bypass_6_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_0_data_21 <= io_in_r_bypass_7_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_0_load_store_21 <= io_in_r_bypass_7_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_0_df_is_ws_21 <= io_in_r_bypass_7_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_0_stall_21 <= io_in_r_bypass_7_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_1_data_21 <= io_in_r_bypass_7_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_1_load_store_21 <= io_in_r_bypass_7_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_1_df_is_ws_21 <= io_in_r_bypass_7_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_1_stall_21 <= io_in_r_bypass_7_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_2_data_21 <= io_in_r_bypass_7_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_2_load_store_21 <= io_in_r_bypass_7_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_2_df_is_ws_21 <= io_in_r_bypass_7_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_2_stall_21 <= io_in_r_bypass_7_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_3_data_21 <= io_in_r_bypass_7_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_3_load_store_21 <= io_in_r_bypass_7_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_3_df_is_ws_21 <= io_in_r_bypass_7_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_3_stall_21 <= io_in_r_bypass_7_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_0_data_21 <= io_in_r_bypass_8_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_0_load_store_21 <= io_in_r_bypass_8_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_0_df_is_ws_21 <= io_in_r_bypass_8_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_0_stall_21 <= io_in_r_bypass_8_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_1_data_21 <= io_in_r_bypass_8_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_1_load_store_21 <= io_in_r_bypass_8_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_1_df_is_ws_21 <= io_in_r_bypass_8_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_1_stall_21 <= io_in_r_bypass_8_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_2_data_21 <= io_in_r_bypass_8_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_2_load_store_21 <= io_in_r_bypass_8_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_2_df_is_ws_21 <= io_in_r_bypass_8_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_2_stall_21 <= io_in_r_bypass_8_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_3_data_21 <= io_in_r_bypass_8_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_3_load_store_21 <= io_in_r_bypass_8_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_3_df_is_ws_21 <= io_in_r_bypass_8_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_3_stall_21 <= io_in_r_bypass_8_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_0_data_21 <= io_in_r_bypass_9_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_0_load_store_21 <= io_in_r_bypass_9_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_0_df_is_ws_21 <= io_in_r_bypass_9_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_0_stall_21 <= io_in_r_bypass_9_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_1_data_21 <= io_in_r_bypass_9_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_1_load_store_21 <= io_in_r_bypass_9_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_1_df_is_ws_21 <= io_in_r_bypass_9_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_1_stall_21 <= io_in_r_bypass_9_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_2_data_21 <= io_in_r_bypass_9_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_2_load_store_21 <= io_in_r_bypass_9_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_2_df_is_ws_21 <= io_in_r_bypass_9_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_2_stall_21 <= io_in_r_bypass_9_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_3_data_21 <= io_in_r_bypass_9_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_3_load_store_21 <= io_in_r_bypass_9_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_3_df_is_ws_21 <= io_in_r_bypass_9_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_3_stall_21 <= io_in_r_bypass_9_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_0_data_21 <= io_in_r_bypass_10_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_0_load_store_21 <= io_in_r_bypass_10_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_0_df_is_ws_21 <= io_in_r_bypass_10_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_0_stall_21 <= io_in_r_bypass_10_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_1_data_21 <= io_in_r_bypass_10_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_1_load_store_21 <= io_in_r_bypass_10_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_1_df_is_ws_21 <= io_in_r_bypass_10_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_1_stall_21 <= io_in_r_bypass_10_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_2_data_21 <= io_in_r_bypass_10_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_2_load_store_21 <= io_in_r_bypass_10_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_2_df_is_ws_21 <= io_in_r_bypass_10_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_2_stall_21 <= io_in_r_bypass_10_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_3_data_21 <= io_in_r_bypass_10_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_3_load_store_21 <= io_in_r_bypass_10_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_3_df_is_ws_21 <= io_in_r_bypass_10_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_3_stall_21 <= io_in_r_bypass_10_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_0_data_21 <= io_in_r_bypass_11_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_0_load_store_21 <= io_in_r_bypass_11_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_0_df_is_ws_21 <= io_in_r_bypass_11_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_0_stall_21 <= io_in_r_bypass_11_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_1_data_21 <= io_in_r_bypass_11_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_1_load_store_21 <= io_in_r_bypass_11_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_1_df_is_ws_21 <= io_in_r_bypass_11_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_1_stall_21 <= io_in_r_bypass_11_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_2_data_21 <= io_in_r_bypass_11_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_2_load_store_21 <= io_in_r_bypass_11_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_2_df_is_ws_21 <= io_in_r_bypass_11_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_2_stall_21 <= io_in_r_bypass_11_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_3_data_21 <= io_in_r_bypass_11_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_3_load_store_21 <= io_in_r_bypass_11_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_3_df_is_ws_21 <= io_in_r_bypass_11_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_3_stall_21 <= io_in_r_bypass_11_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_0_data_21 <= io_in_r_bypass_12_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_0_load_store_21 <= io_in_r_bypass_12_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_0_df_is_ws_21 <= io_in_r_bypass_12_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_0_stall_21 <= io_in_r_bypass_12_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_1_data_21 <= io_in_r_bypass_12_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_1_load_store_21 <= io_in_r_bypass_12_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_1_df_is_ws_21 <= io_in_r_bypass_12_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_1_stall_21 <= io_in_r_bypass_12_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_2_data_21 <= io_in_r_bypass_12_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_2_load_store_21 <= io_in_r_bypass_12_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_2_df_is_ws_21 <= io_in_r_bypass_12_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_2_stall_21 <= io_in_r_bypass_12_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_3_data_21 <= io_in_r_bypass_12_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_3_load_store_21 <= io_in_r_bypass_12_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_3_df_is_ws_21 <= io_in_r_bypass_12_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_3_stall_21 <= io_in_r_bypass_12_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_0_data_21 <= io_in_r_bypass_13_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_0_load_store_21 <= io_in_r_bypass_13_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_0_df_is_ws_21 <= io_in_r_bypass_13_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_0_stall_21 <= io_in_r_bypass_13_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_1_data_21 <= io_in_r_bypass_13_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_1_load_store_21 <= io_in_r_bypass_13_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_1_df_is_ws_21 <= io_in_r_bypass_13_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_1_stall_21 <= io_in_r_bypass_13_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_2_data_21 <= io_in_r_bypass_13_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_2_load_store_21 <= io_in_r_bypass_13_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_2_df_is_ws_21 <= io_in_r_bypass_13_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_2_stall_21 <= io_in_r_bypass_13_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_3_data_21 <= io_in_r_bypass_13_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_3_load_store_21 <= io_in_r_bypass_13_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_3_df_is_ws_21 <= io_in_r_bypass_13_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_3_stall_21 <= io_in_r_bypass_13_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_0_data_21 <= io_in_r_bypass_14_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_0_load_store_21 <= io_in_r_bypass_14_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_0_df_is_ws_21 <= io_in_r_bypass_14_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_0_stall_21 <= io_in_r_bypass_14_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_1_data_21 <= io_in_r_bypass_14_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_1_load_store_21 <= io_in_r_bypass_14_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_1_df_is_ws_21 <= io_in_r_bypass_14_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_1_stall_21 <= io_in_r_bypass_14_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_2_data_21 <= io_in_r_bypass_14_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_2_load_store_21 <= io_in_r_bypass_14_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_2_df_is_ws_21 <= io_in_r_bypass_14_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_2_stall_21 <= io_in_r_bypass_14_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_3_data_21 <= io_in_r_bypass_14_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_3_load_store_21 <= io_in_r_bypass_14_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_3_df_is_ws_21 <= io_in_r_bypass_14_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_3_stall_21 <= io_in_r_bypass_14_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_0_data_21 <= io_in_r_bypass_15_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_0_load_store_21 <= io_in_r_bypass_15_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_0_df_is_ws_21 <= io_in_r_bypass_15_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_0_stall_21 <= io_in_r_bypass_15_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_1_data_21 <= io_in_r_bypass_15_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_1_load_store_21 <= io_in_r_bypass_15_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_1_df_is_ws_21 <= io_in_r_bypass_15_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_1_stall_21 <= io_in_r_bypass_15_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_2_data_21 <= io_in_r_bypass_15_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_2_load_store_21 <= io_in_r_bypass_15_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_2_df_is_ws_21 <= io_in_r_bypass_15_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_2_stall_21 <= io_in_r_bypass_15_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_3_data_21 <= io_in_r_bypass_15_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_3_load_store_21 <= io_in_r_bypass_15_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_3_df_is_ws_21 <= io_in_r_bypass_15_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_3_stall_21 <= io_in_r_bypass_15_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_0_data_21 <= io_in_r_bypass_16_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_0_load_store_21 <= io_in_r_bypass_16_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_0_df_is_ws_21 <= io_in_r_bypass_16_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_0_stall_21 <= io_in_r_bypass_16_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_1_data_21 <= io_in_r_bypass_16_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_1_load_store_21 <= io_in_r_bypass_16_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_1_df_is_ws_21 <= io_in_r_bypass_16_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_1_stall_21 <= io_in_r_bypass_16_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_2_data_21 <= io_in_r_bypass_16_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_2_load_store_21 <= io_in_r_bypass_16_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_2_df_is_ws_21 <= io_in_r_bypass_16_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_2_stall_21 <= io_in_r_bypass_16_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_3_data_21 <= io_in_r_bypass_16_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_3_load_store_21 <= io_in_r_bypass_16_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_3_df_is_ws_21 <= io_in_r_bypass_16_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_3_stall_21 <= io_in_r_bypass_16_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_0_data_21 <= io_in_r_bypass_17_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_0_load_store_21 <= io_in_r_bypass_17_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_0_df_is_ws_21 <= io_in_r_bypass_17_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_0_stall_21 <= io_in_r_bypass_17_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_1_data_21 <= io_in_r_bypass_17_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_1_load_store_21 <= io_in_r_bypass_17_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_1_df_is_ws_21 <= io_in_r_bypass_17_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_1_stall_21 <= io_in_r_bypass_17_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_2_data_21 <= io_in_r_bypass_17_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_2_load_store_21 <= io_in_r_bypass_17_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_2_df_is_ws_21 <= io_in_r_bypass_17_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_2_stall_21 <= io_in_r_bypass_17_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_3_data_21 <= io_in_r_bypass_17_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_3_load_store_21 <= io_in_r_bypass_17_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_3_df_is_ws_21 <= io_in_r_bypass_17_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_3_stall_21 <= io_in_r_bypass_17_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_0_data_21 <= io_in_r_bypass_18_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_0_load_store_21 <= io_in_r_bypass_18_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_0_df_is_ws_21 <= io_in_r_bypass_18_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_0_stall_21 <= io_in_r_bypass_18_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_1_data_21 <= io_in_r_bypass_18_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_1_load_store_21 <= io_in_r_bypass_18_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_1_df_is_ws_21 <= io_in_r_bypass_18_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_1_stall_21 <= io_in_r_bypass_18_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_2_data_21 <= io_in_r_bypass_18_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_2_load_store_21 <= io_in_r_bypass_18_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_2_df_is_ws_21 <= io_in_r_bypass_18_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_2_stall_21 <= io_in_r_bypass_18_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_3_data_21 <= io_in_r_bypass_18_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_3_load_store_21 <= io_in_r_bypass_18_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_3_df_is_ws_21 <= io_in_r_bypass_18_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_3_stall_21 <= io_in_r_bypass_18_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_0_data_21 <= io_in_r_bypass_19_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_0_load_store_21 <= io_in_r_bypass_19_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_0_df_is_ws_21 <= io_in_r_bypass_19_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_0_stall_21 <= io_in_r_bypass_19_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_1_data_21 <= io_in_r_bypass_19_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_1_load_store_21 <= io_in_r_bypass_19_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_1_df_is_ws_21 <= io_in_r_bypass_19_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_1_stall_21 <= io_in_r_bypass_19_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_2_data_21 <= io_in_r_bypass_19_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_2_load_store_21 <= io_in_r_bypass_19_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_2_df_is_ws_21 <= io_in_r_bypass_19_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_2_stall_21 <= io_in_r_bypass_19_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_3_data_21 <= io_in_r_bypass_19_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_3_load_store_21 <= io_in_r_bypass_19_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_3_df_is_ws_21 <= io_in_r_bypass_19_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_3_stall_21 <= io_in_r_bypass_19_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_0_data_21 <= io_in_r_bypass_20_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_0_load_store_21 <= io_in_r_bypass_20_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_0_df_is_ws_21 <= io_in_r_bypass_20_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_0_stall_21 <= io_in_r_bypass_20_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_1_data_21 <= io_in_r_bypass_20_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_1_load_store_21 <= io_in_r_bypass_20_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_1_df_is_ws_21 <= io_in_r_bypass_20_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_1_stall_21 <= io_in_r_bypass_20_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_2_data_21 <= io_in_r_bypass_20_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_2_load_store_21 <= io_in_r_bypass_20_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_2_df_is_ws_21 <= io_in_r_bypass_20_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_2_stall_21 <= io_in_r_bypass_20_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_3_data_21 <= io_in_r_bypass_20_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_3_load_store_21 <= io_in_r_bypass_20_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_3_df_is_ws_21 <= io_in_r_bypass_20_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_3_stall_21 <= io_in_r_bypass_20_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_0_data_21 <= io_in_r_bypass_21_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_0_load_store_21 <= io_in_r_bypass_21_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_0_df_is_ws_21 <= io_in_r_bypass_21_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_0_stall_21 <= io_in_r_bypass_21_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_1_data_21 <= io_in_r_bypass_21_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_1_load_store_21 <= io_in_r_bypass_21_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_1_df_is_ws_21 <= io_in_r_bypass_21_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_1_stall_21 <= io_in_r_bypass_21_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_2_data_21 <= io_in_r_bypass_21_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_2_load_store_21 <= io_in_r_bypass_21_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_2_df_is_ws_21 <= io_in_r_bypass_21_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_2_stall_21 <= io_in_r_bypass_21_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_3_data_21 <= io_in_r_bypass_21_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_3_load_store_21 <= io_in_r_bypass_21_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_3_df_is_ws_21 <= io_in_r_bypass_21_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_3_stall_21 <= io_in_r_bypass_21_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_0_data_21 <= io_in_r_bypass_22_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_0_load_store_21 <= io_in_r_bypass_22_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_0_df_is_ws_21 <= io_in_r_bypass_22_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_0_stall_21 <= io_in_r_bypass_22_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_1_data_21 <= io_in_r_bypass_22_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_1_load_store_21 <= io_in_r_bypass_22_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_1_df_is_ws_21 <= io_in_r_bypass_22_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_1_stall_21 <= io_in_r_bypass_22_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_2_data_21 <= io_in_r_bypass_22_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_2_load_store_21 <= io_in_r_bypass_22_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_2_df_is_ws_21 <= io_in_r_bypass_22_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_2_stall_21 <= io_in_r_bypass_22_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_3_data_21 <= io_in_r_bypass_22_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_3_load_store_21 <= io_in_r_bypass_22_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_3_df_is_ws_21 <= io_in_r_bypass_22_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_3_stall_21 <= io_in_r_bypass_22_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_0_data_21 <= io_in_r_bypass_23_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_0_load_store_21 <= io_in_r_bypass_23_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_0_df_is_ws_21 <= io_in_r_bypass_23_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_0_stall_21 <= io_in_r_bypass_23_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_1_data_21 <= io_in_r_bypass_23_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_1_load_store_21 <= io_in_r_bypass_23_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_1_df_is_ws_21 <= io_in_r_bypass_23_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_1_stall_21 <= io_in_r_bypass_23_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_2_data_21 <= io_in_r_bypass_23_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_2_load_store_21 <= io_in_r_bypass_23_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_2_df_is_ws_21 <= io_in_r_bypass_23_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_2_stall_21 <= io_in_r_bypass_23_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_3_data_21 <= io_in_r_bypass_23_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_3_load_store_21 <= io_in_r_bypass_23_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_3_df_is_ws_21 <= io_in_r_bypass_23_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_3_stall_21 <= io_in_r_bypass_23_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_0_data_21 <= io_in_r_bypass_24_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_0_load_store_21 <= io_in_r_bypass_24_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_0_df_is_ws_21 <= io_in_r_bypass_24_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_0_stall_21 <= io_in_r_bypass_24_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_1_data_21 <= io_in_r_bypass_24_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_1_load_store_21 <= io_in_r_bypass_24_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_1_df_is_ws_21 <= io_in_r_bypass_24_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_1_stall_21 <= io_in_r_bypass_24_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_2_data_21 <= io_in_r_bypass_24_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_2_load_store_21 <= io_in_r_bypass_24_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_2_df_is_ws_21 <= io_in_r_bypass_24_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_2_stall_21 <= io_in_r_bypass_24_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_3_data_21 <= io_in_r_bypass_24_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_3_load_store_21 <= io_in_r_bypass_24_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_3_df_is_ws_21 <= io_in_r_bypass_24_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_3_stall_21 <= io_in_r_bypass_24_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_0_data_21 <= io_in_r_bypass_25_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_0_load_store_21 <= io_in_r_bypass_25_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_0_df_is_ws_21 <= io_in_r_bypass_25_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_0_stall_21 <= io_in_r_bypass_25_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_1_data_21 <= io_in_r_bypass_25_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_1_load_store_21 <= io_in_r_bypass_25_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_1_df_is_ws_21 <= io_in_r_bypass_25_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_1_stall_21 <= io_in_r_bypass_25_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_2_data_21 <= io_in_r_bypass_25_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_2_load_store_21 <= io_in_r_bypass_25_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_2_df_is_ws_21 <= io_in_r_bypass_25_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_2_stall_21 <= io_in_r_bypass_25_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_3_data_21 <= io_in_r_bypass_25_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_3_load_store_21 <= io_in_r_bypass_25_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_3_df_is_ws_21 <= io_in_r_bypass_25_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_3_stall_21 <= io_in_r_bypass_25_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_0_data_21 <= io_in_r_bypass_26_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_0_load_store_21 <= io_in_r_bypass_26_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_0_df_is_ws_21 <= io_in_r_bypass_26_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_0_stall_21 <= io_in_r_bypass_26_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_1_data_21 <= io_in_r_bypass_26_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_1_load_store_21 <= io_in_r_bypass_26_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_1_df_is_ws_21 <= io_in_r_bypass_26_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_1_stall_21 <= io_in_r_bypass_26_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_2_data_21 <= io_in_r_bypass_26_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_2_load_store_21 <= io_in_r_bypass_26_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_2_df_is_ws_21 <= io_in_r_bypass_26_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_2_stall_21 <= io_in_r_bypass_26_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_3_data_21 <= io_in_r_bypass_26_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_3_load_store_21 <= io_in_r_bypass_26_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_3_df_is_ws_21 <= io_in_r_bypass_26_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_3_stall_21 <= io_in_r_bypass_26_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_0_data_21 <= io_in_r_bypass_27_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_0_load_store_21 <= io_in_r_bypass_27_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_0_df_is_ws_21 <= io_in_r_bypass_27_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_0_stall_21 <= io_in_r_bypass_27_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_1_data_21 <= io_in_r_bypass_27_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_1_load_store_21 <= io_in_r_bypass_27_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_1_df_is_ws_21 <= io_in_r_bypass_27_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_1_stall_21 <= io_in_r_bypass_27_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_2_data_21 <= io_in_r_bypass_27_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_2_load_store_21 <= io_in_r_bypass_27_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_2_df_is_ws_21 <= io_in_r_bypass_27_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_2_stall_21 <= io_in_r_bypass_27_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_3_data_21 <= io_in_r_bypass_27_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_3_load_store_21 <= io_in_r_bypass_27_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_3_df_is_ws_21 <= io_in_r_bypass_27_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_3_stall_21 <= io_in_r_bypass_27_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_0_data_21 <= io_in_r_bypass_28_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_0_load_store_21 <= io_in_r_bypass_28_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_0_df_is_ws_21 <= io_in_r_bypass_28_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_0_stall_21 <= io_in_r_bypass_28_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_1_data_21 <= io_in_r_bypass_28_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_1_load_store_21 <= io_in_r_bypass_28_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_1_df_is_ws_21 <= io_in_r_bypass_28_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_1_stall_21 <= io_in_r_bypass_28_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_2_data_21 <= io_in_r_bypass_28_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_2_load_store_21 <= io_in_r_bypass_28_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_2_df_is_ws_21 <= io_in_r_bypass_28_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_2_stall_21 <= io_in_r_bypass_28_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_3_data_21 <= io_in_r_bypass_28_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_3_load_store_21 <= io_in_r_bypass_28_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_3_df_is_ws_21 <= io_in_r_bypass_28_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_3_stall_21 <= io_in_r_bypass_28_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_0_data_21 <= io_in_r_bypass_29_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_0_load_store_21 <= io_in_r_bypass_29_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_0_df_is_ws_21 <= io_in_r_bypass_29_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_0_stall_21 <= io_in_r_bypass_29_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_1_data_21 <= io_in_r_bypass_29_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_1_load_store_21 <= io_in_r_bypass_29_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_1_df_is_ws_21 <= io_in_r_bypass_29_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_1_stall_21 <= io_in_r_bypass_29_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_2_data_21 <= io_in_r_bypass_29_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_2_load_store_21 <= io_in_r_bypass_29_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_2_df_is_ws_21 <= io_in_r_bypass_29_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_2_stall_21 <= io_in_r_bypass_29_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_3_data_21 <= io_in_r_bypass_29_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_3_load_store_21 <= io_in_r_bypass_29_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_3_df_is_ws_21 <= io_in_r_bypass_29_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_3_stall_21 <= io_in_r_bypass_29_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_0_data_21 <= io_in_r_bypass_30_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_0_load_store_21 <= io_in_r_bypass_30_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_0_df_is_ws_21 <= io_in_r_bypass_30_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_0_stall_21 <= io_in_r_bypass_30_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_1_data_21 <= io_in_r_bypass_30_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_1_load_store_21 <= io_in_r_bypass_30_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_1_df_is_ws_21 <= io_in_r_bypass_30_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_1_stall_21 <= io_in_r_bypass_30_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_2_data_21 <= io_in_r_bypass_30_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_2_load_store_21 <= io_in_r_bypass_30_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_2_df_is_ws_21 <= io_in_r_bypass_30_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_2_stall_21 <= io_in_r_bypass_30_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_3_data_21 <= io_in_r_bypass_30_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_3_load_store_21 <= io_in_r_bypass_30_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_3_df_is_ws_21 <= io_in_r_bypass_30_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_3_stall_21 <= io_in_r_bypass_30_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_0_data_21 <= io_in_r_bypass_31_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_0_load_store_21 <= io_in_r_bypass_31_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_0_df_is_ws_21 <= io_in_r_bypass_31_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_0_stall_21 <= io_in_r_bypass_31_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_1_data_21 <= io_in_r_bypass_31_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_1_load_store_21 <= io_in_r_bypass_31_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_1_df_is_ws_21 <= io_in_r_bypass_31_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_1_stall_21 <= io_in_r_bypass_31_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_2_data_21 <= io_in_r_bypass_31_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_2_load_store_21 <= io_in_r_bypass_31_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_2_df_is_ws_21 <= io_in_r_bypass_31_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_2_stall_21 <= io_in_r_bypass_31_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_3_data_21 <= io_in_r_bypass_31_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_3_load_store_21 <= io_in_r_bypass_31_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_3_df_is_ws_21 <= io_in_r_bypass_31_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_3_stall_21 <= io_in_r_bypass_31_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_0_data_22 <= io_in_r_bypass_0_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_0_load_store_22 <= io_in_r_bypass_0_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_0_df_is_ws_22 <= io_in_r_bypass_0_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_0_stall_22 <= io_in_r_bypass_0_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_1_data_22 <= io_in_r_bypass_0_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_1_load_store_22 <= io_in_r_bypass_0_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_1_df_is_ws_22 <= io_in_r_bypass_0_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_1_stall_22 <= io_in_r_bypass_0_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_2_data_22 <= io_in_r_bypass_0_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_2_load_store_22 <= io_in_r_bypass_0_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_2_df_is_ws_22 <= io_in_r_bypass_0_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_2_stall_22 <= io_in_r_bypass_0_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_3_data_22 <= io_in_r_bypass_0_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_3_load_store_22 <= io_in_r_bypass_0_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_3_df_is_ws_22 <= io_in_r_bypass_0_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_3_stall_22 <= io_in_r_bypass_0_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_0_data_22 <= io_in_r_bypass_1_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_0_load_store_22 <= io_in_r_bypass_1_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_0_df_is_ws_22 <= io_in_r_bypass_1_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_0_stall_22 <= io_in_r_bypass_1_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_1_data_22 <= io_in_r_bypass_1_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_1_load_store_22 <= io_in_r_bypass_1_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_1_df_is_ws_22 <= io_in_r_bypass_1_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_1_stall_22 <= io_in_r_bypass_1_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_2_data_22 <= io_in_r_bypass_1_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_2_load_store_22 <= io_in_r_bypass_1_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_2_df_is_ws_22 <= io_in_r_bypass_1_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_2_stall_22 <= io_in_r_bypass_1_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_3_data_22 <= io_in_r_bypass_1_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_3_load_store_22 <= io_in_r_bypass_1_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_3_df_is_ws_22 <= io_in_r_bypass_1_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_3_stall_22 <= io_in_r_bypass_1_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_0_data_22 <= io_in_r_bypass_2_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_0_load_store_22 <= io_in_r_bypass_2_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_0_df_is_ws_22 <= io_in_r_bypass_2_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_0_stall_22 <= io_in_r_bypass_2_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_1_data_22 <= io_in_r_bypass_2_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_1_load_store_22 <= io_in_r_bypass_2_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_1_df_is_ws_22 <= io_in_r_bypass_2_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_1_stall_22 <= io_in_r_bypass_2_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_2_data_22 <= io_in_r_bypass_2_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_2_load_store_22 <= io_in_r_bypass_2_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_2_df_is_ws_22 <= io_in_r_bypass_2_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_2_stall_22 <= io_in_r_bypass_2_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_3_data_22 <= io_in_r_bypass_2_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_3_load_store_22 <= io_in_r_bypass_2_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_3_df_is_ws_22 <= io_in_r_bypass_2_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_3_stall_22 <= io_in_r_bypass_2_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_0_data_22 <= io_in_r_bypass_3_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_0_load_store_22 <= io_in_r_bypass_3_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_0_df_is_ws_22 <= io_in_r_bypass_3_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_0_stall_22 <= io_in_r_bypass_3_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_1_data_22 <= io_in_r_bypass_3_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_1_load_store_22 <= io_in_r_bypass_3_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_1_df_is_ws_22 <= io_in_r_bypass_3_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_1_stall_22 <= io_in_r_bypass_3_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_2_data_22 <= io_in_r_bypass_3_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_2_load_store_22 <= io_in_r_bypass_3_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_2_df_is_ws_22 <= io_in_r_bypass_3_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_2_stall_22 <= io_in_r_bypass_3_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_3_data_22 <= io_in_r_bypass_3_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_3_load_store_22 <= io_in_r_bypass_3_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_3_df_is_ws_22 <= io_in_r_bypass_3_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_3_stall_22 <= io_in_r_bypass_3_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_0_data_22 <= io_in_r_bypass_4_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_0_load_store_22 <= io_in_r_bypass_4_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_0_df_is_ws_22 <= io_in_r_bypass_4_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_0_stall_22 <= io_in_r_bypass_4_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_1_data_22 <= io_in_r_bypass_4_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_1_load_store_22 <= io_in_r_bypass_4_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_1_df_is_ws_22 <= io_in_r_bypass_4_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_1_stall_22 <= io_in_r_bypass_4_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_2_data_22 <= io_in_r_bypass_4_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_2_load_store_22 <= io_in_r_bypass_4_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_2_df_is_ws_22 <= io_in_r_bypass_4_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_2_stall_22 <= io_in_r_bypass_4_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_3_data_22 <= io_in_r_bypass_4_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_3_load_store_22 <= io_in_r_bypass_4_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_3_df_is_ws_22 <= io_in_r_bypass_4_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_3_stall_22 <= io_in_r_bypass_4_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_0_data_22 <= io_in_r_bypass_5_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_0_load_store_22 <= io_in_r_bypass_5_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_0_df_is_ws_22 <= io_in_r_bypass_5_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_0_stall_22 <= io_in_r_bypass_5_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_1_data_22 <= io_in_r_bypass_5_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_1_load_store_22 <= io_in_r_bypass_5_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_1_df_is_ws_22 <= io_in_r_bypass_5_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_1_stall_22 <= io_in_r_bypass_5_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_2_data_22 <= io_in_r_bypass_5_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_2_load_store_22 <= io_in_r_bypass_5_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_2_df_is_ws_22 <= io_in_r_bypass_5_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_2_stall_22 <= io_in_r_bypass_5_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_3_data_22 <= io_in_r_bypass_5_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_3_load_store_22 <= io_in_r_bypass_5_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_3_df_is_ws_22 <= io_in_r_bypass_5_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_3_stall_22 <= io_in_r_bypass_5_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_0_data_22 <= io_in_r_bypass_6_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_0_load_store_22 <= io_in_r_bypass_6_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_0_df_is_ws_22 <= io_in_r_bypass_6_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_0_stall_22 <= io_in_r_bypass_6_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_1_data_22 <= io_in_r_bypass_6_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_1_load_store_22 <= io_in_r_bypass_6_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_1_df_is_ws_22 <= io_in_r_bypass_6_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_1_stall_22 <= io_in_r_bypass_6_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_2_data_22 <= io_in_r_bypass_6_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_2_load_store_22 <= io_in_r_bypass_6_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_2_df_is_ws_22 <= io_in_r_bypass_6_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_2_stall_22 <= io_in_r_bypass_6_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_3_data_22 <= io_in_r_bypass_6_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_3_load_store_22 <= io_in_r_bypass_6_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_3_df_is_ws_22 <= io_in_r_bypass_6_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_3_stall_22 <= io_in_r_bypass_6_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_0_data_22 <= io_in_r_bypass_7_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_0_load_store_22 <= io_in_r_bypass_7_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_0_df_is_ws_22 <= io_in_r_bypass_7_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_0_stall_22 <= io_in_r_bypass_7_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_1_data_22 <= io_in_r_bypass_7_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_1_load_store_22 <= io_in_r_bypass_7_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_1_df_is_ws_22 <= io_in_r_bypass_7_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_1_stall_22 <= io_in_r_bypass_7_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_2_data_22 <= io_in_r_bypass_7_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_2_load_store_22 <= io_in_r_bypass_7_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_2_df_is_ws_22 <= io_in_r_bypass_7_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_2_stall_22 <= io_in_r_bypass_7_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_3_data_22 <= io_in_r_bypass_7_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_3_load_store_22 <= io_in_r_bypass_7_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_3_df_is_ws_22 <= io_in_r_bypass_7_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_3_stall_22 <= io_in_r_bypass_7_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_0_data_22 <= io_in_r_bypass_8_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_0_load_store_22 <= io_in_r_bypass_8_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_0_df_is_ws_22 <= io_in_r_bypass_8_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_0_stall_22 <= io_in_r_bypass_8_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_1_data_22 <= io_in_r_bypass_8_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_1_load_store_22 <= io_in_r_bypass_8_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_1_df_is_ws_22 <= io_in_r_bypass_8_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_1_stall_22 <= io_in_r_bypass_8_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_2_data_22 <= io_in_r_bypass_8_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_2_load_store_22 <= io_in_r_bypass_8_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_2_df_is_ws_22 <= io_in_r_bypass_8_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_2_stall_22 <= io_in_r_bypass_8_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_3_data_22 <= io_in_r_bypass_8_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_3_load_store_22 <= io_in_r_bypass_8_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_3_df_is_ws_22 <= io_in_r_bypass_8_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_3_stall_22 <= io_in_r_bypass_8_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_0_data_22 <= io_in_r_bypass_9_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_0_load_store_22 <= io_in_r_bypass_9_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_0_df_is_ws_22 <= io_in_r_bypass_9_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_0_stall_22 <= io_in_r_bypass_9_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_1_data_22 <= io_in_r_bypass_9_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_1_load_store_22 <= io_in_r_bypass_9_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_1_df_is_ws_22 <= io_in_r_bypass_9_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_1_stall_22 <= io_in_r_bypass_9_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_2_data_22 <= io_in_r_bypass_9_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_2_load_store_22 <= io_in_r_bypass_9_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_2_df_is_ws_22 <= io_in_r_bypass_9_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_2_stall_22 <= io_in_r_bypass_9_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_3_data_22 <= io_in_r_bypass_9_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_3_load_store_22 <= io_in_r_bypass_9_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_3_df_is_ws_22 <= io_in_r_bypass_9_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_3_stall_22 <= io_in_r_bypass_9_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_0_data_22 <= io_in_r_bypass_10_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_0_load_store_22 <= io_in_r_bypass_10_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_0_df_is_ws_22 <= io_in_r_bypass_10_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_0_stall_22 <= io_in_r_bypass_10_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_1_data_22 <= io_in_r_bypass_10_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_1_load_store_22 <= io_in_r_bypass_10_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_1_df_is_ws_22 <= io_in_r_bypass_10_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_1_stall_22 <= io_in_r_bypass_10_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_2_data_22 <= io_in_r_bypass_10_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_2_load_store_22 <= io_in_r_bypass_10_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_2_df_is_ws_22 <= io_in_r_bypass_10_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_2_stall_22 <= io_in_r_bypass_10_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_3_data_22 <= io_in_r_bypass_10_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_3_load_store_22 <= io_in_r_bypass_10_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_3_df_is_ws_22 <= io_in_r_bypass_10_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_3_stall_22 <= io_in_r_bypass_10_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_0_data_22 <= io_in_r_bypass_11_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_0_load_store_22 <= io_in_r_bypass_11_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_0_df_is_ws_22 <= io_in_r_bypass_11_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_0_stall_22 <= io_in_r_bypass_11_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_1_data_22 <= io_in_r_bypass_11_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_1_load_store_22 <= io_in_r_bypass_11_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_1_df_is_ws_22 <= io_in_r_bypass_11_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_1_stall_22 <= io_in_r_bypass_11_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_2_data_22 <= io_in_r_bypass_11_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_2_load_store_22 <= io_in_r_bypass_11_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_2_df_is_ws_22 <= io_in_r_bypass_11_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_2_stall_22 <= io_in_r_bypass_11_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_3_data_22 <= io_in_r_bypass_11_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_3_load_store_22 <= io_in_r_bypass_11_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_3_df_is_ws_22 <= io_in_r_bypass_11_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_3_stall_22 <= io_in_r_bypass_11_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_0_data_22 <= io_in_r_bypass_12_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_0_load_store_22 <= io_in_r_bypass_12_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_0_df_is_ws_22 <= io_in_r_bypass_12_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_0_stall_22 <= io_in_r_bypass_12_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_1_data_22 <= io_in_r_bypass_12_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_1_load_store_22 <= io_in_r_bypass_12_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_1_df_is_ws_22 <= io_in_r_bypass_12_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_1_stall_22 <= io_in_r_bypass_12_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_2_data_22 <= io_in_r_bypass_12_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_2_load_store_22 <= io_in_r_bypass_12_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_2_df_is_ws_22 <= io_in_r_bypass_12_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_2_stall_22 <= io_in_r_bypass_12_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_3_data_22 <= io_in_r_bypass_12_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_3_load_store_22 <= io_in_r_bypass_12_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_3_df_is_ws_22 <= io_in_r_bypass_12_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_3_stall_22 <= io_in_r_bypass_12_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_0_data_22 <= io_in_r_bypass_13_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_0_load_store_22 <= io_in_r_bypass_13_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_0_df_is_ws_22 <= io_in_r_bypass_13_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_0_stall_22 <= io_in_r_bypass_13_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_1_data_22 <= io_in_r_bypass_13_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_1_load_store_22 <= io_in_r_bypass_13_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_1_df_is_ws_22 <= io_in_r_bypass_13_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_1_stall_22 <= io_in_r_bypass_13_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_2_data_22 <= io_in_r_bypass_13_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_2_load_store_22 <= io_in_r_bypass_13_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_2_df_is_ws_22 <= io_in_r_bypass_13_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_2_stall_22 <= io_in_r_bypass_13_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_3_data_22 <= io_in_r_bypass_13_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_3_load_store_22 <= io_in_r_bypass_13_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_3_df_is_ws_22 <= io_in_r_bypass_13_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_3_stall_22 <= io_in_r_bypass_13_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_0_data_22 <= io_in_r_bypass_14_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_0_load_store_22 <= io_in_r_bypass_14_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_0_df_is_ws_22 <= io_in_r_bypass_14_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_0_stall_22 <= io_in_r_bypass_14_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_1_data_22 <= io_in_r_bypass_14_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_1_load_store_22 <= io_in_r_bypass_14_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_1_df_is_ws_22 <= io_in_r_bypass_14_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_1_stall_22 <= io_in_r_bypass_14_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_2_data_22 <= io_in_r_bypass_14_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_2_load_store_22 <= io_in_r_bypass_14_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_2_df_is_ws_22 <= io_in_r_bypass_14_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_2_stall_22 <= io_in_r_bypass_14_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_3_data_22 <= io_in_r_bypass_14_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_3_load_store_22 <= io_in_r_bypass_14_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_3_df_is_ws_22 <= io_in_r_bypass_14_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_3_stall_22 <= io_in_r_bypass_14_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_0_data_22 <= io_in_r_bypass_15_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_0_load_store_22 <= io_in_r_bypass_15_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_0_df_is_ws_22 <= io_in_r_bypass_15_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_0_stall_22 <= io_in_r_bypass_15_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_1_data_22 <= io_in_r_bypass_15_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_1_load_store_22 <= io_in_r_bypass_15_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_1_df_is_ws_22 <= io_in_r_bypass_15_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_1_stall_22 <= io_in_r_bypass_15_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_2_data_22 <= io_in_r_bypass_15_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_2_load_store_22 <= io_in_r_bypass_15_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_2_df_is_ws_22 <= io_in_r_bypass_15_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_2_stall_22 <= io_in_r_bypass_15_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_3_data_22 <= io_in_r_bypass_15_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_3_load_store_22 <= io_in_r_bypass_15_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_3_df_is_ws_22 <= io_in_r_bypass_15_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_3_stall_22 <= io_in_r_bypass_15_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_0_data_22 <= io_in_r_bypass_16_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_0_load_store_22 <= io_in_r_bypass_16_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_0_df_is_ws_22 <= io_in_r_bypass_16_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_0_stall_22 <= io_in_r_bypass_16_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_1_data_22 <= io_in_r_bypass_16_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_1_load_store_22 <= io_in_r_bypass_16_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_1_df_is_ws_22 <= io_in_r_bypass_16_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_1_stall_22 <= io_in_r_bypass_16_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_2_data_22 <= io_in_r_bypass_16_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_2_load_store_22 <= io_in_r_bypass_16_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_2_df_is_ws_22 <= io_in_r_bypass_16_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_2_stall_22 <= io_in_r_bypass_16_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_3_data_22 <= io_in_r_bypass_16_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_3_load_store_22 <= io_in_r_bypass_16_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_3_df_is_ws_22 <= io_in_r_bypass_16_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_3_stall_22 <= io_in_r_bypass_16_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_0_data_22 <= io_in_r_bypass_17_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_0_load_store_22 <= io_in_r_bypass_17_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_0_df_is_ws_22 <= io_in_r_bypass_17_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_0_stall_22 <= io_in_r_bypass_17_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_1_data_22 <= io_in_r_bypass_17_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_1_load_store_22 <= io_in_r_bypass_17_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_1_df_is_ws_22 <= io_in_r_bypass_17_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_1_stall_22 <= io_in_r_bypass_17_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_2_data_22 <= io_in_r_bypass_17_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_2_load_store_22 <= io_in_r_bypass_17_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_2_df_is_ws_22 <= io_in_r_bypass_17_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_2_stall_22 <= io_in_r_bypass_17_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_3_data_22 <= io_in_r_bypass_17_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_3_load_store_22 <= io_in_r_bypass_17_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_3_df_is_ws_22 <= io_in_r_bypass_17_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_3_stall_22 <= io_in_r_bypass_17_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_0_data_22 <= io_in_r_bypass_18_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_0_load_store_22 <= io_in_r_bypass_18_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_0_df_is_ws_22 <= io_in_r_bypass_18_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_0_stall_22 <= io_in_r_bypass_18_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_1_data_22 <= io_in_r_bypass_18_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_1_load_store_22 <= io_in_r_bypass_18_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_1_df_is_ws_22 <= io_in_r_bypass_18_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_1_stall_22 <= io_in_r_bypass_18_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_2_data_22 <= io_in_r_bypass_18_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_2_load_store_22 <= io_in_r_bypass_18_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_2_df_is_ws_22 <= io_in_r_bypass_18_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_2_stall_22 <= io_in_r_bypass_18_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_3_data_22 <= io_in_r_bypass_18_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_3_load_store_22 <= io_in_r_bypass_18_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_3_df_is_ws_22 <= io_in_r_bypass_18_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_3_stall_22 <= io_in_r_bypass_18_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_0_data_22 <= io_in_r_bypass_19_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_0_load_store_22 <= io_in_r_bypass_19_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_0_df_is_ws_22 <= io_in_r_bypass_19_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_0_stall_22 <= io_in_r_bypass_19_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_1_data_22 <= io_in_r_bypass_19_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_1_load_store_22 <= io_in_r_bypass_19_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_1_df_is_ws_22 <= io_in_r_bypass_19_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_1_stall_22 <= io_in_r_bypass_19_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_2_data_22 <= io_in_r_bypass_19_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_2_load_store_22 <= io_in_r_bypass_19_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_2_df_is_ws_22 <= io_in_r_bypass_19_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_2_stall_22 <= io_in_r_bypass_19_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_3_data_22 <= io_in_r_bypass_19_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_3_load_store_22 <= io_in_r_bypass_19_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_3_df_is_ws_22 <= io_in_r_bypass_19_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_3_stall_22 <= io_in_r_bypass_19_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_0_data_22 <= io_in_r_bypass_20_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_0_load_store_22 <= io_in_r_bypass_20_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_0_df_is_ws_22 <= io_in_r_bypass_20_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_0_stall_22 <= io_in_r_bypass_20_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_1_data_22 <= io_in_r_bypass_20_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_1_load_store_22 <= io_in_r_bypass_20_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_1_df_is_ws_22 <= io_in_r_bypass_20_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_1_stall_22 <= io_in_r_bypass_20_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_2_data_22 <= io_in_r_bypass_20_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_2_load_store_22 <= io_in_r_bypass_20_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_2_df_is_ws_22 <= io_in_r_bypass_20_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_2_stall_22 <= io_in_r_bypass_20_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_3_data_22 <= io_in_r_bypass_20_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_3_load_store_22 <= io_in_r_bypass_20_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_3_df_is_ws_22 <= io_in_r_bypass_20_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_3_stall_22 <= io_in_r_bypass_20_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_0_data_22 <= io_in_r_bypass_21_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_0_load_store_22 <= io_in_r_bypass_21_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_0_df_is_ws_22 <= io_in_r_bypass_21_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_0_stall_22 <= io_in_r_bypass_21_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_1_data_22 <= io_in_r_bypass_21_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_1_load_store_22 <= io_in_r_bypass_21_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_1_df_is_ws_22 <= io_in_r_bypass_21_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_1_stall_22 <= io_in_r_bypass_21_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_2_data_22 <= io_in_r_bypass_21_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_2_load_store_22 <= io_in_r_bypass_21_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_2_df_is_ws_22 <= io_in_r_bypass_21_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_2_stall_22 <= io_in_r_bypass_21_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_3_data_22 <= io_in_r_bypass_21_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_3_load_store_22 <= io_in_r_bypass_21_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_3_df_is_ws_22 <= io_in_r_bypass_21_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_3_stall_22 <= io_in_r_bypass_21_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_0_data_22 <= io_in_r_bypass_22_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_0_load_store_22 <= io_in_r_bypass_22_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_0_df_is_ws_22 <= io_in_r_bypass_22_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_0_stall_22 <= io_in_r_bypass_22_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_1_data_22 <= io_in_r_bypass_22_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_1_load_store_22 <= io_in_r_bypass_22_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_1_df_is_ws_22 <= io_in_r_bypass_22_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_1_stall_22 <= io_in_r_bypass_22_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_2_data_22 <= io_in_r_bypass_22_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_2_load_store_22 <= io_in_r_bypass_22_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_2_df_is_ws_22 <= io_in_r_bypass_22_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_2_stall_22 <= io_in_r_bypass_22_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_3_data_22 <= io_in_r_bypass_22_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_3_load_store_22 <= io_in_r_bypass_22_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_3_df_is_ws_22 <= io_in_r_bypass_22_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_3_stall_22 <= io_in_r_bypass_22_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_0_data_22 <= io_in_r_bypass_23_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_0_load_store_22 <= io_in_r_bypass_23_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_0_df_is_ws_22 <= io_in_r_bypass_23_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_0_stall_22 <= io_in_r_bypass_23_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_1_data_22 <= io_in_r_bypass_23_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_1_load_store_22 <= io_in_r_bypass_23_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_1_df_is_ws_22 <= io_in_r_bypass_23_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_1_stall_22 <= io_in_r_bypass_23_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_2_data_22 <= io_in_r_bypass_23_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_2_load_store_22 <= io_in_r_bypass_23_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_2_df_is_ws_22 <= io_in_r_bypass_23_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_2_stall_22 <= io_in_r_bypass_23_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_3_data_22 <= io_in_r_bypass_23_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_3_load_store_22 <= io_in_r_bypass_23_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_3_df_is_ws_22 <= io_in_r_bypass_23_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_3_stall_22 <= io_in_r_bypass_23_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_0_data_22 <= io_in_r_bypass_24_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_0_load_store_22 <= io_in_r_bypass_24_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_0_df_is_ws_22 <= io_in_r_bypass_24_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_0_stall_22 <= io_in_r_bypass_24_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_1_data_22 <= io_in_r_bypass_24_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_1_load_store_22 <= io_in_r_bypass_24_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_1_df_is_ws_22 <= io_in_r_bypass_24_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_1_stall_22 <= io_in_r_bypass_24_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_2_data_22 <= io_in_r_bypass_24_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_2_load_store_22 <= io_in_r_bypass_24_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_2_df_is_ws_22 <= io_in_r_bypass_24_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_2_stall_22 <= io_in_r_bypass_24_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_3_data_22 <= io_in_r_bypass_24_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_3_load_store_22 <= io_in_r_bypass_24_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_3_df_is_ws_22 <= io_in_r_bypass_24_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_3_stall_22 <= io_in_r_bypass_24_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_0_data_22 <= io_in_r_bypass_25_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_0_load_store_22 <= io_in_r_bypass_25_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_0_df_is_ws_22 <= io_in_r_bypass_25_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_0_stall_22 <= io_in_r_bypass_25_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_1_data_22 <= io_in_r_bypass_25_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_1_load_store_22 <= io_in_r_bypass_25_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_1_df_is_ws_22 <= io_in_r_bypass_25_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_1_stall_22 <= io_in_r_bypass_25_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_2_data_22 <= io_in_r_bypass_25_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_2_load_store_22 <= io_in_r_bypass_25_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_2_df_is_ws_22 <= io_in_r_bypass_25_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_2_stall_22 <= io_in_r_bypass_25_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_3_data_22 <= io_in_r_bypass_25_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_3_load_store_22 <= io_in_r_bypass_25_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_3_df_is_ws_22 <= io_in_r_bypass_25_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_3_stall_22 <= io_in_r_bypass_25_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_0_data_22 <= io_in_r_bypass_26_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_0_load_store_22 <= io_in_r_bypass_26_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_0_df_is_ws_22 <= io_in_r_bypass_26_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_0_stall_22 <= io_in_r_bypass_26_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_1_data_22 <= io_in_r_bypass_26_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_1_load_store_22 <= io_in_r_bypass_26_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_1_df_is_ws_22 <= io_in_r_bypass_26_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_1_stall_22 <= io_in_r_bypass_26_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_2_data_22 <= io_in_r_bypass_26_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_2_load_store_22 <= io_in_r_bypass_26_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_2_df_is_ws_22 <= io_in_r_bypass_26_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_2_stall_22 <= io_in_r_bypass_26_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_3_data_22 <= io_in_r_bypass_26_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_3_load_store_22 <= io_in_r_bypass_26_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_3_df_is_ws_22 <= io_in_r_bypass_26_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_3_stall_22 <= io_in_r_bypass_26_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_0_data_22 <= io_in_r_bypass_27_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_0_load_store_22 <= io_in_r_bypass_27_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_0_df_is_ws_22 <= io_in_r_bypass_27_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_0_stall_22 <= io_in_r_bypass_27_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_1_data_22 <= io_in_r_bypass_27_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_1_load_store_22 <= io_in_r_bypass_27_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_1_df_is_ws_22 <= io_in_r_bypass_27_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_1_stall_22 <= io_in_r_bypass_27_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_2_data_22 <= io_in_r_bypass_27_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_2_load_store_22 <= io_in_r_bypass_27_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_2_df_is_ws_22 <= io_in_r_bypass_27_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_2_stall_22 <= io_in_r_bypass_27_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_3_data_22 <= io_in_r_bypass_27_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_3_load_store_22 <= io_in_r_bypass_27_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_3_df_is_ws_22 <= io_in_r_bypass_27_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_3_stall_22 <= io_in_r_bypass_27_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_0_data_22 <= io_in_r_bypass_28_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_0_load_store_22 <= io_in_r_bypass_28_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_0_df_is_ws_22 <= io_in_r_bypass_28_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_0_stall_22 <= io_in_r_bypass_28_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_1_data_22 <= io_in_r_bypass_28_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_1_load_store_22 <= io_in_r_bypass_28_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_1_df_is_ws_22 <= io_in_r_bypass_28_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_1_stall_22 <= io_in_r_bypass_28_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_2_data_22 <= io_in_r_bypass_28_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_2_load_store_22 <= io_in_r_bypass_28_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_2_df_is_ws_22 <= io_in_r_bypass_28_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_2_stall_22 <= io_in_r_bypass_28_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_3_data_22 <= io_in_r_bypass_28_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_3_load_store_22 <= io_in_r_bypass_28_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_3_df_is_ws_22 <= io_in_r_bypass_28_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_3_stall_22 <= io_in_r_bypass_28_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_0_data_22 <= io_in_r_bypass_29_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_0_load_store_22 <= io_in_r_bypass_29_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_0_df_is_ws_22 <= io_in_r_bypass_29_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_0_stall_22 <= io_in_r_bypass_29_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_1_data_22 <= io_in_r_bypass_29_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_1_load_store_22 <= io_in_r_bypass_29_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_1_df_is_ws_22 <= io_in_r_bypass_29_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_1_stall_22 <= io_in_r_bypass_29_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_2_data_22 <= io_in_r_bypass_29_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_2_load_store_22 <= io_in_r_bypass_29_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_2_df_is_ws_22 <= io_in_r_bypass_29_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_2_stall_22 <= io_in_r_bypass_29_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_3_data_22 <= io_in_r_bypass_29_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_3_load_store_22 <= io_in_r_bypass_29_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_3_df_is_ws_22 <= io_in_r_bypass_29_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_3_stall_22 <= io_in_r_bypass_29_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_0_data_22 <= io_in_r_bypass_30_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_0_load_store_22 <= io_in_r_bypass_30_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_0_df_is_ws_22 <= io_in_r_bypass_30_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_0_stall_22 <= io_in_r_bypass_30_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_1_data_22 <= io_in_r_bypass_30_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_1_load_store_22 <= io_in_r_bypass_30_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_1_df_is_ws_22 <= io_in_r_bypass_30_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_1_stall_22 <= io_in_r_bypass_30_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_2_data_22 <= io_in_r_bypass_30_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_2_load_store_22 <= io_in_r_bypass_30_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_2_df_is_ws_22 <= io_in_r_bypass_30_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_2_stall_22 <= io_in_r_bypass_30_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_3_data_22 <= io_in_r_bypass_30_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_3_load_store_22 <= io_in_r_bypass_30_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_3_df_is_ws_22 <= io_in_r_bypass_30_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_3_stall_22 <= io_in_r_bypass_30_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_0_data_22 <= io_in_r_bypass_31_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_0_load_store_22 <= io_in_r_bypass_31_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_0_df_is_ws_22 <= io_in_r_bypass_31_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_0_stall_22 <= io_in_r_bypass_31_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_1_data_22 <= io_in_r_bypass_31_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_1_load_store_22 <= io_in_r_bypass_31_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_1_df_is_ws_22 <= io_in_r_bypass_31_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_1_stall_22 <= io_in_r_bypass_31_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_2_data_22 <= io_in_r_bypass_31_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_2_load_store_22 <= io_in_r_bypass_31_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_2_df_is_ws_22 <= io_in_r_bypass_31_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_2_stall_22 <= io_in_r_bypass_31_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_3_data_22 <= io_in_r_bypass_31_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_3_load_store_22 <= io_in_r_bypass_31_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_3_df_is_ws_22 <= io_in_r_bypass_31_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_3_stall_22 <= io_in_r_bypass_31_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_0_data_23 <= io_in_r_bypass_0_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_0_load_store_23 <= io_in_r_bypass_0_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_0_df_is_ws_23 <= io_in_r_bypass_0_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_0_stall_23 <= io_in_r_bypass_0_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_1_data_23 <= io_in_r_bypass_0_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_1_load_store_23 <= io_in_r_bypass_0_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_1_df_is_ws_23 <= io_in_r_bypass_0_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_1_stall_23 <= io_in_r_bypass_0_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_2_data_23 <= io_in_r_bypass_0_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_2_load_store_23 <= io_in_r_bypass_0_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_2_df_is_ws_23 <= io_in_r_bypass_0_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_2_stall_23 <= io_in_r_bypass_0_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_3_data_23 <= io_in_r_bypass_0_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_3_load_store_23 <= io_in_r_bypass_0_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_3_df_is_ws_23 <= io_in_r_bypass_0_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_3_stall_23 <= io_in_r_bypass_0_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_0_data_23 <= io_in_r_bypass_1_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_0_load_store_23 <= io_in_r_bypass_1_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_0_df_is_ws_23 <= io_in_r_bypass_1_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_0_stall_23 <= io_in_r_bypass_1_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_1_data_23 <= io_in_r_bypass_1_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_1_load_store_23 <= io_in_r_bypass_1_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_1_df_is_ws_23 <= io_in_r_bypass_1_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_1_stall_23 <= io_in_r_bypass_1_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_2_data_23 <= io_in_r_bypass_1_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_2_load_store_23 <= io_in_r_bypass_1_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_2_df_is_ws_23 <= io_in_r_bypass_1_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_2_stall_23 <= io_in_r_bypass_1_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_3_data_23 <= io_in_r_bypass_1_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_3_load_store_23 <= io_in_r_bypass_1_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_3_df_is_ws_23 <= io_in_r_bypass_1_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_3_stall_23 <= io_in_r_bypass_1_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_0_data_23 <= io_in_r_bypass_2_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_0_load_store_23 <= io_in_r_bypass_2_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_0_df_is_ws_23 <= io_in_r_bypass_2_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_0_stall_23 <= io_in_r_bypass_2_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_1_data_23 <= io_in_r_bypass_2_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_1_load_store_23 <= io_in_r_bypass_2_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_1_df_is_ws_23 <= io_in_r_bypass_2_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_1_stall_23 <= io_in_r_bypass_2_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_2_data_23 <= io_in_r_bypass_2_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_2_load_store_23 <= io_in_r_bypass_2_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_2_df_is_ws_23 <= io_in_r_bypass_2_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_2_stall_23 <= io_in_r_bypass_2_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_3_data_23 <= io_in_r_bypass_2_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_3_load_store_23 <= io_in_r_bypass_2_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_3_df_is_ws_23 <= io_in_r_bypass_2_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_3_stall_23 <= io_in_r_bypass_2_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_0_data_23 <= io_in_r_bypass_3_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_0_load_store_23 <= io_in_r_bypass_3_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_0_df_is_ws_23 <= io_in_r_bypass_3_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_0_stall_23 <= io_in_r_bypass_3_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_1_data_23 <= io_in_r_bypass_3_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_1_load_store_23 <= io_in_r_bypass_3_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_1_df_is_ws_23 <= io_in_r_bypass_3_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_1_stall_23 <= io_in_r_bypass_3_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_2_data_23 <= io_in_r_bypass_3_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_2_load_store_23 <= io_in_r_bypass_3_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_2_df_is_ws_23 <= io_in_r_bypass_3_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_2_stall_23 <= io_in_r_bypass_3_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_3_data_23 <= io_in_r_bypass_3_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_3_load_store_23 <= io_in_r_bypass_3_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_3_df_is_ws_23 <= io_in_r_bypass_3_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_3_stall_23 <= io_in_r_bypass_3_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_0_data_23 <= io_in_r_bypass_4_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_0_load_store_23 <= io_in_r_bypass_4_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_0_df_is_ws_23 <= io_in_r_bypass_4_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_0_stall_23 <= io_in_r_bypass_4_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_1_data_23 <= io_in_r_bypass_4_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_1_load_store_23 <= io_in_r_bypass_4_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_1_df_is_ws_23 <= io_in_r_bypass_4_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_1_stall_23 <= io_in_r_bypass_4_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_2_data_23 <= io_in_r_bypass_4_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_2_load_store_23 <= io_in_r_bypass_4_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_2_df_is_ws_23 <= io_in_r_bypass_4_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_2_stall_23 <= io_in_r_bypass_4_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_3_data_23 <= io_in_r_bypass_4_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_3_load_store_23 <= io_in_r_bypass_4_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_3_df_is_ws_23 <= io_in_r_bypass_4_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_3_stall_23 <= io_in_r_bypass_4_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_0_data_23 <= io_in_r_bypass_5_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_0_load_store_23 <= io_in_r_bypass_5_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_0_df_is_ws_23 <= io_in_r_bypass_5_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_0_stall_23 <= io_in_r_bypass_5_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_1_data_23 <= io_in_r_bypass_5_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_1_load_store_23 <= io_in_r_bypass_5_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_1_df_is_ws_23 <= io_in_r_bypass_5_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_1_stall_23 <= io_in_r_bypass_5_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_2_data_23 <= io_in_r_bypass_5_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_2_load_store_23 <= io_in_r_bypass_5_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_2_df_is_ws_23 <= io_in_r_bypass_5_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_2_stall_23 <= io_in_r_bypass_5_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_3_data_23 <= io_in_r_bypass_5_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_3_load_store_23 <= io_in_r_bypass_5_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_3_df_is_ws_23 <= io_in_r_bypass_5_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_3_stall_23 <= io_in_r_bypass_5_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_0_data_23 <= io_in_r_bypass_6_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_0_load_store_23 <= io_in_r_bypass_6_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_0_df_is_ws_23 <= io_in_r_bypass_6_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_0_stall_23 <= io_in_r_bypass_6_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_1_data_23 <= io_in_r_bypass_6_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_1_load_store_23 <= io_in_r_bypass_6_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_1_df_is_ws_23 <= io_in_r_bypass_6_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_1_stall_23 <= io_in_r_bypass_6_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_2_data_23 <= io_in_r_bypass_6_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_2_load_store_23 <= io_in_r_bypass_6_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_2_df_is_ws_23 <= io_in_r_bypass_6_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_2_stall_23 <= io_in_r_bypass_6_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_3_data_23 <= io_in_r_bypass_6_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_3_load_store_23 <= io_in_r_bypass_6_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_3_df_is_ws_23 <= io_in_r_bypass_6_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_3_stall_23 <= io_in_r_bypass_6_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_0_data_23 <= io_in_r_bypass_7_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_0_load_store_23 <= io_in_r_bypass_7_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_0_df_is_ws_23 <= io_in_r_bypass_7_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_0_stall_23 <= io_in_r_bypass_7_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_1_data_23 <= io_in_r_bypass_7_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_1_load_store_23 <= io_in_r_bypass_7_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_1_df_is_ws_23 <= io_in_r_bypass_7_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_1_stall_23 <= io_in_r_bypass_7_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_2_data_23 <= io_in_r_bypass_7_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_2_load_store_23 <= io_in_r_bypass_7_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_2_df_is_ws_23 <= io_in_r_bypass_7_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_2_stall_23 <= io_in_r_bypass_7_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_3_data_23 <= io_in_r_bypass_7_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_3_load_store_23 <= io_in_r_bypass_7_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_3_df_is_ws_23 <= io_in_r_bypass_7_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_3_stall_23 <= io_in_r_bypass_7_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_0_data_23 <= io_in_r_bypass_8_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_0_load_store_23 <= io_in_r_bypass_8_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_0_df_is_ws_23 <= io_in_r_bypass_8_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_0_stall_23 <= io_in_r_bypass_8_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_1_data_23 <= io_in_r_bypass_8_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_1_load_store_23 <= io_in_r_bypass_8_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_1_df_is_ws_23 <= io_in_r_bypass_8_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_1_stall_23 <= io_in_r_bypass_8_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_2_data_23 <= io_in_r_bypass_8_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_2_load_store_23 <= io_in_r_bypass_8_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_2_df_is_ws_23 <= io_in_r_bypass_8_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_2_stall_23 <= io_in_r_bypass_8_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_3_data_23 <= io_in_r_bypass_8_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_3_load_store_23 <= io_in_r_bypass_8_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_3_df_is_ws_23 <= io_in_r_bypass_8_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_3_stall_23 <= io_in_r_bypass_8_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_0_data_23 <= io_in_r_bypass_9_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_0_load_store_23 <= io_in_r_bypass_9_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_0_df_is_ws_23 <= io_in_r_bypass_9_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_0_stall_23 <= io_in_r_bypass_9_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_1_data_23 <= io_in_r_bypass_9_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_1_load_store_23 <= io_in_r_bypass_9_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_1_df_is_ws_23 <= io_in_r_bypass_9_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_1_stall_23 <= io_in_r_bypass_9_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_2_data_23 <= io_in_r_bypass_9_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_2_load_store_23 <= io_in_r_bypass_9_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_2_df_is_ws_23 <= io_in_r_bypass_9_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_2_stall_23 <= io_in_r_bypass_9_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_3_data_23 <= io_in_r_bypass_9_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_3_load_store_23 <= io_in_r_bypass_9_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_3_df_is_ws_23 <= io_in_r_bypass_9_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_3_stall_23 <= io_in_r_bypass_9_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_0_data_23 <= io_in_r_bypass_10_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_0_load_store_23 <= io_in_r_bypass_10_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_0_df_is_ws_23 <= io_in_r_bypass_10_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_0_stall_23 <= io_in_r_bypass_10_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_1_data_23 <= io_in_r_bypass_10_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_1_load_store_23 <= io_in_r_bypass_10_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_1_df_is_ws_23 <= io_in_r_bypass_10_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_1_stall_23 <= io_in_r_bypass_10_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_2_data_23 <= io_in_r_bypass_10_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_2_load_store_23 <= io_in_r_bypass_10_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_2_df_is_ws_23 <= io_in_r_bypass_10_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_2_stall_23 <= io_in_r_bypass_10_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_3_data_23 <= io_in_r_bypass_10_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_3_load_store_23 <= io_in_r_bypass_10_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_3_df_is_ws_23 <= io_in_r_bypass_10_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_3_stall_23 <= io_in_r_bypass_10_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_0_data_23 <= io_in_r_bypass_11_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_0_load_store_23 <= io_in_r_bypass_11_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_0_df_is_ws_23 <= io_in_r_bypass_11_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_0_stall_23 <= io_in_r_bypass_11_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_1_data_23 <= io_in_r_bypass_11_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_1_load_store_23 <= io_in_r_bypass_11_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_1_df_is_ws_23 <= io_in_r_bypass_11_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_1_stall_23 <= io_in_r_bypass_11_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_2_data_23 <= io_in_r_bypass_11_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_2_load_store_23 <= io_in_r_bypass_11_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_2_df_is_ws_23 <= io_in_r_bypass_11_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_2_stall_23 <= io_in_r_bypass_11_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_3_data_23 <= io_in_r_bypass_11_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_3_load_store_23 <= io_in_r_bypass_11_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_3_df_is_ws_23 <= io_in_r_bypass_11_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_3_stall_23 <= io_in_r_bypass_11_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_0_data_23 <= io_in_r_bypass_12_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_0_load_store_23 <= io_in_r_bypass_12_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_0_df_is_ws_23 <= io_in_r_bypass_12_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_0_stall_23 <= io_in_r_bypass_12_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_1_data_23 <= io_in_r_bypass_12_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_1_load_store_23 <= io_in_r_bypass_12_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_1_df_is_ws_23 <= io_in_r_bypass_12_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_1_stall_23 <= io_in_r_bypass_12_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_2_data_23 <= io_in_r_bypass_12_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_2_load_store_23 <= io_in_r_bypass_12_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_2_df_is_ws_23 <= io_in_r_bypass_12_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_2_stall_23 <= io_in_r_bypass_12_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_3_data_23 <= io_in_r_bypass_12_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_3_load_store_23 <= io_in_r_bypass_12_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_3_df_is_ws_23 <= io_in_r_bypass_12_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_3_stall_23 <= io_in_r_bypass_12_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_0_data_23 <= io_in_r_bypass_13_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_0_load_store_23 <= io_in_r_bypass_13_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_0_df_is_ws_23 <= io_in_r_bypass_13_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_0_stall_23 <= io_in_r_bypass_13_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_1_data_23 <= io_in_r_bypass_13_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_1_load_store_23 <= io_in_r_bypass_13_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_1_df_is_ws_23 <= io_in_r_bypass_13_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_1_stall_23 <= io_in_r_bypass_13_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_2_data_23 <= io_in_r_bypass_13_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_2_load_store_23 <= io_in_r_bypass_13_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_2_df_is_ws_23 <= io_in_r_bypass_13_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_2_stall_23 <= io_in_r_bypass_13_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_3_data_23 <= io_in_r_bypass_13_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_3_load_store_23 <= io_in_r_bypass_13_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_3_df_is_ws_23 <= io_in_r_bypass_13_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_3_stall_23 <= io_in_r_bypass_13_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_0_data_23 <= io_in_r_bypass_14_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_0_load_store_23 <= io_in_r_bypass_14_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_0_df_is_ws_23 <= io_in_r_bypass_14_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_0_stall_23 <= io_in_r_bypass_14_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_1_data_23 <= io_in_r_bypass_14_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_1_load_store_23 <= io_in_r_bypass_14_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_1_df_is_ws_23 <= io_in_r_bypass_14_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_1_stall_23 <= io_in_r_bypass_14_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_2_data_23 <= io_in_r_bypass_14_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_2_load_store_23 <= io_in_r_bypass_14_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_2_df_is_ws_23 <= io_in_r_bypass_14_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_2_stall_23 <= io_in_r_bypass_14_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_3_data_23 <= io_in_r_bypass_14_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_3_load_store_23 <= io_in_r_bypass_14_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_3_df_is_ws_23 <= io_in_r_bypass_14_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_3_stall_23 <= io_in_r_bypass_14_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_0_data_23 <= io_in_r_bypass_15_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_0_load_store_23 <= io_in_r_bypass_15_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_0_df_is_ws_23 <= io_in_r_bypass_15_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_0_stall_23 <= io_in_r_bypass_15_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_1_data_23 <= io_in_r_bypass_15_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_1_load_store_23 <= io_in_r_bypass_15_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_1_df_is_ws_23 <= io_in_r_bypass_15_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_1_stall_23 <= io_in_r_bypass_15_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_2_data_23 <= io_in_r_bypass_15_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_2_load_store_23 <= io_in_r_bypass_15_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_2_df_is_ws_23 <= io_in_r_bypass_15_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_2_stall_23 <= io_in_r_bypass_15_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_3_data_23 <= io_in_r_bypass_15_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_3_load_store_23 <= io_in_r_bypass_15_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_3_df_is_ws_23 <= io_in_r_bypass_15_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_3_stall_23 <= io_in_r_bypass_15_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_0_data_23 <= io_in_r_bypass_16_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_0_load_store_23 <= io_in_r_bypass_16_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_0_df_is_ws_23 <= io_in_r_bypass_16_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_0_stall_23 <= io_in_r_bypass_16_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_1_data_23 <= io_in_r_bypass_16_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_1_load_store_23 <= io_in_r_bypass_16_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_1_df_is_ws_23 <= io_in_r_bypass_16_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_1_stall_23 <= io_in_r_bypass_16_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_2_data_23 <= io_in_r_bypass_16_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_2_load_store_23 <= io_in_r_bypass_16_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_2_df_is_ws_23 <= io_in_r_bypass_16_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_2_stall_23 <= io_in_r_bypass_16_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_3_data_23 <= io_in_r_bypass_16_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_3_load_store_23 <= io_in_r_bypass_16_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_3_df_is_ws_23 <= io_in_r_bypass_16_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_3_stall_23 <= io_in_r_bypass_16_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_0_data_23 <= io_in_r_bypass_17_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_0_load_store_23 <= io_in_r_bypass_17_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_0_df_is_ws_23 <= io_in_r_bypass_17_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_0_stall_23 <= io_in_r_bypass_17_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_1_data_23 <= io_in_r_bypass_17_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_1_load_store_23 <= io_in_r_bypass_17_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_1_df_is_ws_23 <= io_in_r_bypass_17_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_1_stall_23 <= io_in_r_bypass_17_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_2_data_23 <= io_in_r_bypass_17_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_2_load_store_23 <= io_in_r_bypass_17_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_2_df_is_ws_23 <= io_in_r_bypass_17_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_2_stall_23 <= io_in_r_bypass_17_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_3_data_23 <= io_in_r_bypass_17_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_3_load_store_23 <= io_in_r_bypass_17_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_3_df_is_ws_23 <= io_in_r_bypass_17_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_3_stall_23 <= io_in_r_bypass_17_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_0_data_23 <= io_in_r_bypass_18_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_0_load_store_23 <= io_in_r_bypass_18_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_0_df_is_ws_23 <= io_in_r_bypass_18_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_0_stall_23 <= io_in_r_bypass_18_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_1_data_23 <= io_in_r_bypass_18_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_1_load_store_23 <= io_in_r_bypass_18_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_1_df_is_ws_23 <= io_in_r_bypass_18_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_1_stall_23 <= io_in_r_bypass_18_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_2_data_23 <= io_in_r_bypass_18_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_2_load_store_23 <= io_in_r_bypass_18_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_2_df_is_ws_23 <= io_in_r_bypass_18_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_2_stall_23 <= io_in_r_bypass_18_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_3_data_23 <= io_in_r_bypass_18_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_3_load_store_23 <= io_in_r_bypass_18_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_3_df_is_ws_23 <= io_in_r_bypass_18_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_3_stall_23 <= io_in_r_bypass_18_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_0_data_23 <= io_in_r_bypass_19_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_0_load_store_23 <= io_in_r_bypass_19_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_0_df_is_ws_23 <= io_in_r_bypass_19_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_0_stall_23 <= io_in_r_bypass_19_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_1_data_23 <= io_in_r_bypass_19_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_1_load_store_23 <= io_in_r_bypass_19_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_1_df_is_ws_23 <= io_in_r_bypass_19_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_1_stall_23 <= io_in_r_bypass_19_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_2_data_23 <= io_in_r_bypass_19_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_2_load_store_23 <= io_in_r_bypass_19_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_2_df_is_ws_23 <= io_in_r_bypass_19_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_2_stall_23 <= io_in_r_bypass_19_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_3_data_23 <= io_in_r_bypass_19_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_3_load_store_23 <= io_in_r_bypass_19_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_3_df_is_ws_23 <= io_in_r_bypass_19_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_3_stall_23 <= io_in_r_bypass_19_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_0_data_23 <= io_in_r_bypass_20_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_0_load_store_23 <= io_in_r_bypass_20_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_0_df_is_ws_23 <= io_in_r_bypass_20_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_0_stall_23 <= io_in_r_bypass_20_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_1_data_23 <= io_in_r_bypass_20_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_1_load_store_23 <= io_in_r_bypass_20_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_1_df_is_ws_23 <= io_in_r_bypass_20_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_1_stall_23 <= io_in_r_bypass_20_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_2_data_23 <= io_in_r_bypass_20_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_2_load_store_23 <= io_in_r_bypass_20_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_2_df_is_ws_23 <= io_in_r_bypass_20_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_2_stall_23 <= io_in_r_bypass_20_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_3_data_23 <= io_in_r_bypass_20_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_3_load_store_23 <= io_in_r_bypass_20_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_3_df_is_ws_23 <= io_in_r_bypass_20_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_3_stall_23 <= io_in_r_bypass_20_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_0_data_23 <= io_in_r_bypass_21_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_0_load_store_23 <= io_in_r_bypass_21_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_0_df_is_ws_23 <= io_in_r_bypass_21_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_0_stall_23 <= io_in_r_bypass_21_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_1_data_23 <= io_in_r_bypass_21_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_1_load_store_23 <= io_in_r_bypass_21_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_1_df_is_ws_23 <= io_in_r_bypass_21_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_1_stall_23 <= io_in_r_bypass_21_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_2_data_23 <= io_in_r_bypass_21_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_2_load_store_23 <= io_in_r_bypass_21_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_2_df_is_ws_23 <= io_in_r_bypass_21_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_2_stall_23 <= io_in_r_bypass_21_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_3_data_23 <= io_in_r_bypass_21_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_3_load_store_23 <= io_in_r_bypass_21_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_3_df_is_ws_23 <= io_in_r_bypass_21_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_3_stall_23 <= io_in_r_bypass_21_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_0_data_23 <= io_in_r_bypass_22_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_0_load_store_23 <= io_in_r_bypass_22_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_0_df_is_ws_23 <= io_in_r_bypass_22_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_0_stall_23 <= io_in_r_bypass_22_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_1_data_23 <= io_in_r_bypass_22_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_1_load_store_23 <= io_in_r_bypass_22_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_1_df_is_ws_23 <= io_in_r_bypass_22_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_1_stall_23 <= io_in_r_bypass_22_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_2_data_23 <= io_in_r_bypass_22_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_2_load_store_23 <= io_in_r_bypass_22_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_2_df_is_ws_23 <= io_in_r_bypass_22_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_2_stall_23 <= io_in_r_bypass_22_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_3_data_23 <= io_in_r_bypass_22_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_3_load_store_23 <= io_in_r_bypass_22_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_3_df_is_ws_23 <= io_in_r_bypass_22_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_3_stall_23 <= io_in_r_bypass_22_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_0_data_23 <= io_in_r_bypass_23_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_0_load_store_23 <= io_in_r_bypass_23_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_0_df_is_ws_23 <= io_in_r_bypass_23_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_0_stall_23 <= io_in_r_bypass_23_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_1_data_23 <= io_in_r_bypass_23_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_1_load_store_23 <= io_in_r_bypass_23_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_1_df_is_ws_23 <= io_in_r_bypass_23_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_1_stall_23 <= io_in_r_bypass_23_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_2_data_23 <= io_in_r_bypass_23_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_2_load_store_23 <= io_in_r_bypass_23_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_2_df_is_ws_23 <= io_in_r_bypass_23_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_2_stall_23 <= io_in_r_bypass_23_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_3_data_23 <= io_in_r_bypass_23_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_3_load_store_23 <= io_in_r_bypass_23_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_3_df_is_ws_23 <= io_in_r_bypass_23_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_3_stall_23 <= io_in_r_bypass_23_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_0_data_23 <= io_in_r_bypass_24_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_0_load_store_23 <= io_in_r_bypass_24_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_0_df_is_ws_23 <= io_in_r_bypass_24_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_0_stall_23 <= io_in_r_bypass_24_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_1_data_23 <= io_in_r_bypass_24_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_1_load_store_23 <= io_in_r_bypass_24_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_1_df_is_ws_23 <= io_in_r_bypass_24_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_1_stall_23 <= io_in_r_bypass_24_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_2_data_23 <= io_in_r_bypass_24_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_2_load_store_23 <= io_in_r_bypass_24_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_2_df_is_ws_23 <= io_in_r_bypass_24_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_2_stall_23 <= io_in_r_bypass_24_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_3_data_23 <= io_in_r_bypass_24_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_3_load_store_23 <= io_in_r_bypass_24_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_3_df_is_ws_23 <= io_in_r_bypass_24_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_3_stall_23 <= io_in_r_bypass_24_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_0_data_23 <= io_in_r_bypass_25_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_0_load_store_23 <= io_in_r_bypass_25_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_0_df_is_ws_23 <= io_in_r_bypass_25_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_0_stall_23 <= io_in_r_bypass_25_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_1_data_23 <= io_in_r_bypass_25_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_1_load_store_23 <= io_in_r_bypass_25_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_1_df_is_ws_23 <= io_in_r_bypass_25_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_1_stall_23 <= io_in_r_bypass_25_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_2_data_23 <= io_in_r_bypass_25_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_2_load_store_23 <= io_in_r_bypass_25_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_2_df_is_ws_23 <= io_in_r_bypass_25_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_2_stall_23 <= io_in_r_bypass_25_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_3_data_23 <= io_in_r_bypass_25_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_3_load_store_23 <= io_in_r_bypass_25_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_3_df_is_ws_23 <= io_in_r_bypass_25_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_3_stall_23 <= io_in_r_bypass_25_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_0_data_23 <= io_in_r_bypass_26_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_0_load_store_23 <= io_in_r_bypass_26_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_0_df_is_ws_23 <= io_in_r_bypass_26_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_0_stall_23 <= io_in_r_bypass_26_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_1_data_23 <= io_in_r_bypass_26_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_1_load_store_23 <= io_in_r_bypass_26_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_1_df_is_ws_23 <= io_in_r_bypass_26_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_1_stall_23 <= io_in_r_bypass_26_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_2_data_23 <= io_in_r_bypass_26_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_2_load_store_23 <= io_in_r_bypass_26_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_2_df_is_ws_23 <= io_in_r_bypass_26_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_2_stall_23 <= io_in_r_bypass_26_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_3_data_23 <= io_in_r_bypass_26_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_3_load_store_23 <= io_in_r_bypass_26_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_3_df_is_ws_23 <= io_in_r_bypass_26_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_3_stall_23 <= io_in_r_bypass_26_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_0_data_23 <= io_in_r_bypass_27_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_0_load_store_23 <= io_in_r_bypass_27_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_0_df_is_ws_23 <= io_in_r_bypass_27_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_0_stall_23 <= io_in_r_bypass_27_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_1_data_23 <= io_in_r_bypass_27_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_1_load_store_23 <= io_in_r_bypass_27_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_1_df_is_ws_23 <= io_in_r_bypass_27_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_1_stall_23 <= io_in_r_bypass_27_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_2_data_23 <= io_in_r_bypass_27_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_2_load_store_23 <= io_in_r_bypass_27_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_2_df_is_ws_23 <= io_in_r_bypass_27_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_2_stall_23 <= io_in_r_bypass_27_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_3_data_23 <= io_in_r_bypass_27_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_3_load_store_23 <= io_in_r_bypass_27_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_3_df_is_ws_23 <= io_in_r_bypass_27_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_3_stall_23 <= io_in_r_bypass_27_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_0_data_23 <= io_in_r_bypass_28_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_0_load_store_23 <= io_in_r_bypass_28_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_0_df_is_ws_23 <= io_in_r_bypass_28_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_0_stall_23 <= io_in_r_bypass_28_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_1_data_23 <= io_in_r_bypass_28_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_1_load_store_23 <= io_in_r_bypass_28_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_1_df_is_ws_23 <= io_in_r_bypass_28_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_1_stall_23 <= io_in_r_bypass_28_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_2_data_23 <= io_in_r_bypass_28_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_2_load_store_23 <= io_in_r_bypass_28_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_2_df_is_ws_23 <= io_in_r_bypass_28_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_2_stall_23 <= io_in_r_bypass_28_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_3_data_23 <= io_in_r_bypass_28_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_3_load_store_23 <= io_in_r_bypass_28_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_3_df_is_ws_23 <= io_in_r_bypass_28_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_3_stall_23 <= io_in_r_bypass_28_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_0_data_23 <= io_in_r_bypass_29_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_0_load_store_23 <= io_in_r_bypass_29_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_0_df_is_ws_23 <= io_in_r_bypass_29_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_0_stall_23 <= io_in_r_bypass_29_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_1_data_23 <= io_in_r_bypass_29_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_1_load_store_23 <= io_in_r_bypass_29_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_1_df_is_ws_23 <= io_in_r_bypass_29_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_1_stall_23 <= io_in_r_bypass_29_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_2_data_23 <= io_in_r_bypass_29_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_2_load_store_23 <= io_in_r_bypass_29_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_2_df_is_ws_23 <= io_in_r_bypass_29_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_2_stall_23 <= io_in_r_bypass_29_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_3_data_23 <= io_in_r_bypass_29_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_3_load_store_23 <= io_in_r_bypass_29_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_3_df_is_ws_23 <= io_in_r_bypass_29_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_3_stall_23 <= io_in_r_bypass_29_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_0_data_23 <= io_in_r_bypass_30_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_0_load_store_23 <= io_in_r_bypass_30_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_0_df_is_ws_23 <= io_in_r_bypass_30_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_0_stall_23 <= io_in_r_bypass_30_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_1_data_23 <= io_in_r_bypass_30_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_1_load_store_23 <= io_in_r_bypass_30_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_1_df_is_ws_23 <= io_in_r_bypass_30_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_1_stall_23 <= io_in_r_bypass_30_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_2_data_23 <= io_in_r_bypass_30_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_2_load_store_23 <= io_in_r_bypass_30_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_2_df_is_ws_23 <= io_in_r_bypass_30_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_2_stall_23 <= io_in_r_bypass_30_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_3_data_23 <= io_in_r_bypass_30_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_3_load_store_23 <= io_in_r_bypass_30_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_3_df_is_ws_23 <= io_in_r_bypass_30_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_3_stall_23 <= io_in_r_bypass_30_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_0_data_23 <= io_in_r_bypass_31_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_0_load_store_23 <= io_in_r_bypass_31_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_0_df_is_ws_23 <= io_in_r_bypass_31_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_0_stall_23 <= io_in_r_bypass_31_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_1_data_23 <= io_in_r_bypass_31_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_1_load_store_23 <= io_in_r_bypass_31_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_1_df_is_ws_23 <= io_in_r_bypass_31_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_1_stall_23 <= io_in_r_bypass_31_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_2_data_23 <= io_in_r_bypass_31_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_2_load_store_23 <= io_in_r_bypass_31_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_2_df_is_ws_23 <= io_in_r_bypass_31_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_2_stall_23 <= io_in_r_bypass_31_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_3_data_23 <= io_in_r_bypass_31_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_3_load_store_23 <= io_in_r_bypass_31_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_3_df_is_ws_23 <= io_in_r_bypass_31_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_3_stall_23 <= io_in_r_bypass_31_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_0_data_24 <= io_in_r_bypass_0_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_0_load_store_24 <= io_in_r_bypass_0_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_0_df_is_ws_24 <= io_in_r_bypass_0_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_0_stall_24 <= io_in_r_bypass_0_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_1_data_24 <= io_in_r_bypass_0_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_1_load_store_24 <= io_in_r_bypass_0_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_1_df_is_ws_24 <= io_in_r_bypass_0_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_1_stall_24 <= io_in_r_bypass_0_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_2_data_24 <= io_in_r_bypass_0_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_2_load_store_24 <= io_in_r_bypass_0_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_2_df_is_ws_24 <= io_in_r_bypass_0_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_2_stall_24 <= io_in_r_bypass_0_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_3_data_24 <= io_in_r_bypass_0_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_3_load_store_24 <= io_in_r_bypass_0_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_3_df_is_ws_24 <= io_in_r_bypass_0_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_3_stall_24 <= io_in_r_bypass_0_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_0_data_24 <= io_in_r_bypass_1_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_0_load_store_24 <= io_in_r_bypass_1_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_0_df_is_ws_24 <= io_in_r_bypass_1_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_0_stall_24 <= io_in_r_bypass_1_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_1_data_24 <= io_in_r_bypass_1_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_1_load_store_24 <= io_in_r_bypass_1_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_1_df_is_ws_24 <= io_in_r_bypass_1_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_1_stall_24 <= io_in_r_bypass_1_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_2_data_24 <= io_in_r_bypass_1_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_2_load_store_24 <= io_in_r_bypass_1_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_2_df_is_ws_24 <= io_in_r_bypass_1_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_2_stall_24 <= io_in_r_bypass_1_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_3_data_24 <= io_in_r_bypass_1_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_3_load_store_24 <= io_in_r_bypass_1_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_3_df_is_ws_24 <= io_in_r_bypass_1_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_3_stall_24 <= io_in_r_bypass_1_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_0_data_24 <= io_in_r_bypass_2_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_0_load_store_24 <= io_in_r_bypass_2_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_0_df_is_ws_24 <= io_in_r_bypass_2_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_0_stall_24 <= io_in_r_bypass_2_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_1_data_24 <= io_in_r_bypass_2_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_1_load_store_24 <= io_in_r_bypass_2_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_1_df_is_ws_24 <= io_in_r_bypass_2_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_1_stall_24 <= io_in_r_bypass_2_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_2_data_24 <= io_in_r_bypass_2_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_2_load_store_24 <= io_in_r_bypass_2_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_2_df_is_ws_24 <= io_in_r_bypass_2_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_2_stall_24 <= io_in_r_bypass_2_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_3_data_24 <= io_in_r_bypass_2_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_3_load_store_24 <= io_in_r_bypass_2_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_3_df_is_ws_24 <= io_in_r_bypass_2_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_3_stall_24 <= io_in_r_bypass_2_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_0_data_24 <= io_in_r_bypass_3_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_0_load_store_24 <= io_in_r_bypass_3_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_0_df_is_ws_24 <= io_in_r_bypass_3_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_0_stall_24 <= io_in_r_bypass_3_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_1_data_24 <= io_in_r_bypass_3_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_1_load_store_24 <= io_in_r_bypass_3_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_1_df_is_ws_24 <= io_in_r_bypass_3_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_1_stall_24 <= io_in_r_bypass_3_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_2_data_24 <= io_in_r_bypass_3_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_2_load_store_24 <= io_in_r_bypass_3_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_2_df_is_ws_24 <= io_in_r_bypass_3_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_2_stall_24 <= io_in_r_bypass_3_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_3_data_24 <= io_in_r_bypass_3_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_3_load_store_24 <= io_in_r_bypass_3_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_3_df_is_ws_24 <= io_in_r_bypass_3_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_3_stall_24 <= io_in_r_bypass_3_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_0_data_24 <= io_in_r_bypass_4_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_0_load_store_24 <= io_in_r_bypass_4_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_0_df_is_ws_24 <= io_in_r_bypass_4_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_0_stall_24 <= io_in_r_bypass_4_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_1_data_24 <= io_in_r_bypass_4_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_1_load_store_24 <= io_in_r_bypass_4_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_1_df_is_ws_24 <= io_in_r_bypass_4_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_1_stall_24 <= io_in_r_bypass_4_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_2_data_24 <= io_in_r_bypass_4_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_2_load_store_24 <= io_in_r_bypass_4_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_2_df_is_ws_24 <= io_in_r_bypass_4_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_2_stall_24 <= io_in_r_bypass_4_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_3_data_24 <= io_in_r_bypass_4_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_3_load_store_24 <= io_in_r_bypass_4_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_3_df_is_ws_24 <= io_in_r_bypass_4_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_3_stall_24 <= io_in_r_bypass_4_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_0_data_24 <= io_in_r_bypass_5_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_0_load_store_24 <= io_in_r_bypass_5_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_0_df_is_ws_24 <= io_in_r_bypass_5_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_0_stall_24 <= io_in_r_bypass_5_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_1_data_24 <= io_in_r_bypass_5_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_1_load_store_24 <= io_in_r_bypass_5_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_1_df_is_ws_24 <= io_in_r_bypass_5_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_1_stall_24 <= io_in_r_bypass_5_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_2_data_24 <= io_in_r_bypass_5_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_2_load_store_24 <= io_in_r_bypass_5_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_2_df_is_ws_24 <= io_in_r_bypass_5_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_2_stall_24 <= io_in_r_bypass_5_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_3_data_24 <= io_in_r_bypass_5_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_3_load_store_24 <= io_in_r_bypass_5_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_3_df_is_ws_24 <= io_in_r_bypass_5_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_3_stall_24 <= io_in_r_bypass_5_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_0_data_24 <= io_in_r_bypass_6_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_0_load_store_24 <= io_in_r_bypass_6_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_0_df_is_ws_24 <= io_in_r_bypass_6_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_0_stall_24 <= io_in_r_bypass_6_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_1_data_24 <= io_in_r_bypass_6_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_1_load_store_24 <= io_in_r_bypass_6_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_1_df_is_ws_24 <= io_in_r_bypass_6_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_1_stall_24 <= io_in_r_bypass_6_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_2_data_24 <= io_in_r_bypass_6_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_2_load_store_24 <= io_in_r_bypass_6_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_2_df_is_ws_24 <= io_in_r_bypass_6_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_2_stall_24 <= io_in_r_bypass_6_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_3_data_24 <= io_in_r_bypass_6_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_3_load_store_24 <= io_in_r_bypass_6_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_3_df_is_ws_24 <= io_in_r_bypass_6_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_3_stall_24 <= io_in_r_bypass_6_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_0_data_24 <= io_in_r_bypass_7_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_0_load_store_24 <= io_in_r_bypass_7_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_0_df_is_ws_24 <= io_in_r_bypass_7_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_0_stall_24 <= io_in_r_bypass_7_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_1_data_24 <= io_in_r_bypass_7_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_1_load_store_24 <= io_in_r_bypass_7_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_1_df_is_ws_24 <= io_in_r_bypass_7_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_1_stall_24 <= io_in_r_bypass_7_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_2_data_24 <= io_in_r_bypass_7_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_2_load_store_24 <= io_in_r_bypass_7_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_2_df_is_ws_24 <= io_in_r_bypass_7_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_2_stall_24 <= io_in_r_bypass_7_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_3_data_24 <= io_in_r_bypass_7_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_3_load_store_24 <= io_in_r_bypass_7_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_3_df_is_ws_24 <= io_in_r_bypass_7_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_3_stall_24 <= io_in_r_bypass_7_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_0_data_24 <= io_in_r_bypass_8_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_0_load_store_24 <= io_in_r_bypass_8_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_0_df_is_ws_24 <= io_in_r_bypass_8_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_0_stall_24 <= io_in_r_bypass_8_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_1_data_24 <= io_in_r_bypass_8_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_1_load_store_24 <= io_in_r_bypass_8_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_1_df_is_ws_24 <= io_in_r_bypass_8_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_1_stall_24 <= io_in_r_bypass_8_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_2_data_24 <= io_in_r_bypass_8_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_2_load_store_24 <= io_in_r_bypass_8_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_2_df_is_ws_24 <= io_in_r_bypass_8_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_2_stall_24 <= io_in_r_bypass_8_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_3_data_24 <= io_in_r_bypass_8_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_3_load_store_24 <= io_in_r_bypass_8_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_3_df_is_ws_24 <= io_in_r_bypass_8_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_3_stall_24 <= io_in_r_bypass_8_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_0_data_24 <= io_in_r_bypass_9_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_0_load_store_24 <= io_in_r_bypass_9_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_0_df_is_ws_24 <= io_in_r_bypass_9_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_0_stall_24 <= io_in_r_bypass_9_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_1_data_24 <= io_in_r_bypass_9_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_1_load_store_24 <= io_in_r_bypass_9_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_1_df_is_ws_24 <= io_in_r_bypass_9_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_1_stall_24 <= io_in_r_bypass_9_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_2_data_24 <= io_in_r_bypass_9_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_2_load_store_24 <= io_in_r_bypass_9_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_2_df_is_ws_24 <= io_in_r_bypass_9_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_2_stall_24 <= io_in_r_bypass_9_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_3_data_24 <= io_in_r_bypass_9_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_3_load_store_24 <= io_in_r_bypass_9_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_3_df_is_ws_24 <= io_in_r_bypass_9_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_3_stall_24 <= io_in_r_bypass_9_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_0_data_24 <= io_in_r_bypass_10_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_0_load_store_24 <= io_in_r_bypass_10_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_0_df_is_ws_24 <= io_in_r_bypass_10_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_0_stall_24 <= io_in_r_bypass_10_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_1_data_24 <= io_in_r_bypass_10_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_1_load_store_24 <= io_in_r_bypass_10_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_1_df_is_ws_24 <= io_in_r_bypass_10_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_1_stall_24 <= io_in_r_bypass_10_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_2_data_24 <= io_in_r_bypass_10_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_2_load_store_24 <= io_in_r_bypass_10_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_2_df_is_ws_24 <= io_in_r_bypass_10_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_2_stall_24 <= io_in_r_bypass_10_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_3_data_24 <= io_in_r_bypass_10_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_3_load_store_24 <= io_in_r_bypass_10_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_3_df_is_ws_24 <= io_in_r_bypass_10_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_3_stall_24 <= io_in_r_bypass_10_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_0_data_24 <= io_in_r_bypass_11_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_0_load_store_24 <= io_in_r_bypass_11_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_0_df_is_ws_24 <= io_in_r_bypass_11_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_0_stall_24 <= io_in_r_bypass_11_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_1_data_24 <= io_in_r_bypass_11_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_1_load_store_24 <= io_in_r_bypass_11_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_1_df_is_ws_24 <= io_in_r_bypass_11_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_1_stall_24 <= io_in_r_bypass_11_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_2_data_24 <= io_in_r_bypass_11_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_2_load_store_24 <= io_in_r_bypass_11_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_2_df_is_ws_24 <= io_in_r_bypass_11_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_2_stall_24 <= io_in_r_bypass_11_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_3_data_24 <= io_in_r_bypass_11_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_3_load_store_24 <= io_in_r_bypass_11_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_3_df_is_ws_24 <= io_in_r_bypass_11_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_3_stall_24 <= io_in_r_bypass_11_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_0_data_24 <= io_in_r_bypass_12_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_0_load_store_24 <= io_in_r_bypass_12_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_0_df_is_ws_24 <= io_in_r_bypass_12_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_0_stall_24 <= io_in_r_bypass_12_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_1_data_24 <= io_in_r_bypass_12_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_1_load_store_24 <= io_in_r_bypass_12_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_1_df_is_ws_24 <= io_in_r_bypass_12_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_1_stall_24 <= io_in_r_bypass_12_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_2_data_24 <= io_in_r_bypass_12_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_2_load_store_24 <= io_in_r_bypass_12_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_2_df_is_ws_24 <= io_in_r_bypass_12_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_2_stall_24 <= io_in_r_bypass_12_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_3_data_24 <= io_in_r_bypass_12_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_3_load_store_24 <= io_in_r_bypass_12_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_3_df_is_ws_24 <= io_in_r_bypass_12_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_3_stall_24 <= io_in_r_bypass_12_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_0_data_24 <= io_in_r_bypass_13_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_0_load_store_24 <= io_in_r_bypass_13_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_0_df_is_ws_24 <= io_in_r_bypass_13_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_0_stall_24 <= io_in_r_bypass_13_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_1_data_24 <= io_in_r_bypass_13_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_1_load_store_24 <= io_in_r_bypass_13_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_1_df_is_ws_24 <= io_in_r_bypass_13_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_1_stall_24 <= io_in_r_bypass_13_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_2_data_24 <= io_in_r_bypass_13_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_2_load_store_24 <= io_in_r_bypass_13_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_2_df_is_ws_24 <= io_in_r_bypass_13_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_2_stall_24 <= io_in_r_bypass_13_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_3_data_24 <= io_in_r_bypass_13_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_3_load_store_24 <= io_in_r_bypass_13_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_3_df_is_ws_24 <= io_in_r_bypass_13_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_3_stall_24 <= io_in_r_bypass_13_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_0_data_24 <= io_in_r_bypass_14_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_0_load_store_24 <= io_in_r_bypass_14_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_0_df_is_ws_24 <= io_in_r_bypass_14_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_0_stall_24 <= io_in_r_bypass_14_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_1_data_24 <= io_in_r_bypass_14_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_1_load_store_24 <= io_in_r_bypass_14_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_1_df_is_ws_24 <= io_in_r_bypass_14_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_1_stall_24 <= io_in_r_bypass_14_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_2_data_24 <= io_in_r_bypass_14_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_2_load_store_24 <= io_in_r_bypass_14_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_2_df_is_ws_24 <= io_in_r_bypass_14_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_2_stall_24 <= io_in_r_bypass_14_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_3_data_24 <= io_in_r_bypass_14_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_3_load_store_24 <= io_in_r_bypass_14_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_3_df_is_ws_24 <= io_in_r_bypass_14_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_3_stall_24 <= io_in_r_bypass_14_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_0_data_24 <= io_in_r_bypass_15_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_0_load_store_24 <= io_in_r_bypass_15_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_0_df_is_ws_24 <= io_in_r_bypass_15_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_0_stall_24 <= io_in_r_bypass_15_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_1_data_24 <= io_in_r_bypass_15_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_1_load_store_24 <= io_in_r_bypass_15_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_1_df_is_ws_24 <= io_in_r_bypass_15_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_1_stall_24 <= io_in_r_bypass_15_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_2_data_24 <= io_in_r_bypass_15_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_2_load_store_24 <= io_in_r_bypass_15_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_2_df_is_ws_24 <= io_in_r_bypass_15_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_2_stall_24 <= io_in_r_bypass_15_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_3_data_24 <= io_in_r_bypass_15_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_3_load_store_24 <= io_in_r_bypass_15_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_3_df_is_ws_24 <= io_in_r_bypass_15_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_3_stall_24 <= io_in_r_bypass_15_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_0_data_24 <= io_in_r_bypass_16_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_0_load_store_24 <= io_in_r_bypass_16_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_0_df_is_ws_24 <= io_in_r_bypass_16_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_0_stall_24 <= io_in_r_bypass_16_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_1_data_24 <= io_in_r_bypass_16_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_1_load_store_24 <= io_in_r_bypass_16_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_1_df_is_ws_24 <= io_in_r_bypass_16_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_1_stall_24 <= io_in_r_bypass_16_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_2_data_24 <= io_in_r_bypass_16_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_2_load_store_24 <= io_in_r_bypass_16_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_2_df_is_ws_24 <= io_in_r_bypass_16_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_2_stall_24 <= io_in_r_bypass_16_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_3_data_24 <= io_in_r_bypass_16_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_3_load_store_24 <= io_in_r_bypass_16_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_3_df_is_ws_24 <= io_in_r_bypass_16_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_3_stall_24 <= io_in_r_bypass_16_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_0_data_24 <= io_in_r_bypass_17_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_0_load_store_24 <= io_in_r_bypass_17_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_0_df_is_ws_24 <= io_in_r_bypass_17_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_0_stall_24 <= io_in_r_bypass_17_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_1_data_24 <= io_in_r_bypass_17_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_1_load_store_24 <= io_in_r_bypass_17_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_1_df_is_ws_24 <= io_in_r_bypass_17_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_1_stall_24 <= io_in_r_bypass_17_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_2_data_24 <= io_in_r_bypass_17_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_2_load_store_24 <= io_in_r_bypass_17_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_2_df_is_ws_24 <= io_in_r_bypass_17_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_2_stall_24 <= io_in_r_bypass_17_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_3_data_24 <= io_in_r_bypass_17_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_3_load_store_24 <= io_in_r_bypass_17_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_3_df_is_ws_24 <= io_in_r_bypass_17_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_3_stall_24 <= io_in_r_bypass_17_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_0_data_24 <= io_in_r_bypass_18_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_0_load_store_24 <= io_in_r_bypass_18_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_0_df_is_ws_24 <= io_in_r_bypass_18_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_0_stall_24 <= io_in_r_bypass_18_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_1_data_24 <= io_in_r_bypass_18_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_1_load_store_24 <= io_in_r_bypass_18_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_1_df_is_ws_24 <= io_in_r_bypass_18_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_1_stall_24 <= io_in_r_bypass_18_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_2_data_24 <= io_in_r_bypass_18_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_2_load_store_24 <= io_in_r_bypass_18_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_2_df_is_ws_24 <= io_in_r_bypass_18_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_2_stall_24 <= io_in_r_bypass_18_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_3_data_24 <= io_in_r_bypass_18_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_3_load_store_24 <= io_in_r_bypass_18_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_3_df_is_ws_24 <= io_in_r_bypass_18_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_3_stall_24 <= io_in_r_bypass_18_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_0_data_24 <= io_in_r_bypass_19_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_0_load_store_24 <= io_in_r_bypass_19_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_0_df_is_ws_24 <= io_in_r_bypass_19_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_0_stall_24 <= io_in_r_bypass_19_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_1_data_24 <= io_in_r_bypass_19_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_1_load_store_24 <= io_in_r_bypass_19_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_1_df_is_ws_24 <= io_in_r_bypass_19_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_1_stall_24 <= io_in_r_bypass_19_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_2_data_24 <= io_in_r_bypass_19_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_2_load_store_24 <= io_in_r_bypass_19_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_2_df_is_ws_24 <= io_in_r_bypass_19_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_2_stall_24 <= io_in_r_bypass_19_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_3_data_24 <= io_in_r_bypass_19_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_3_load_store_24 <= io_in_r_bypass_19_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_3_df_is_ws_24 <= io_in_r_bypass_19_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_3_stall_24 <= io_in_r_bypass_19_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_0_data_24 <= io_in_r_bypass_20_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_0_load_store_24 <= io_in_r_bypass_20_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_0_df_is_ws_24 <= io_in_r_bypass_20_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_0_stall_24 <= io_in_r_bypass_20_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_1_data_24 <= io_in_r_bypass_20_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_1_load_store_24 <= io_in_r_bypass_20_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_1_df_is_ws_24 <= io_in_r_bypass_20_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_1_stall_24 <= io_in_r_bypass_20_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_2_data_24 <= io_in_r_bypass_20_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_2_load_store_24 <= io_in_r_bypass_20_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_2_df_is_ws_24 <= io_in_r_bypass_20_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_2_stall_24 <= io_in_r_bypass_20_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_3_data_24 <= io_in_r_bypass_20_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_3_load_store_24 <= io_in_r_bypass_20_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_3_df_is_ws_24 <= io_in_r_bypass_20_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_3_stall_24 <= io_in_r_bypass_20_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_0_data_24 <= io_in_r_bypass_21_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_0_load_store_24 <= io_in_r_bypass_21_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_0_df_is_ws_24 <= io_in_r_bypass_21_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_0_stall_24 <= io_in_r_bypass_21_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_1_data_24 <= io_in_r_bypass_21_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_1_load_store_24 <= io_in_r_bypass_21_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_1_df_is_ws_24 <= io_in_r_bypass_21_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_1_stall_24 <= io_in_r_bypass_21_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_2_data_24 <= io_in_r_bypass_21_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_2_load_store_24 <= io_in_r_bypass_21_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_2_df_is_ws_24 <= io_in_r_bypass_21_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_2_stall_24 <= io_in_r_bypass_21_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_3_data_24 <= io_in_r_bypass_21_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_3_load_store_24 <= io_in_r_bypass_21_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_3_df_is_ws_24 <= io_in_r_bypass_21_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_3_stall_24 <= io_in_r_bypass_21_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_0_data_24 <= io_in_r_bypass_22_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_0_load_store_24 <= io_in_r_bypass_22_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_0_df_is_ws_24 <= io_in_r_bypass_22_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_0_stall_24 <= io_in_r_bypass_22_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_1_data_24 <= io_in_r_bypass_22_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_1_load_store_24 <= io_in_r_bypass_22_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_1_df_is_ws_24 <= io_in_r_bypass_22_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_1_stall_24 <= io_in_r_bypass_22_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_2_data_24 <= io_in_r_bypass_22_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_2_load_store_24 <= io_in_r_bypass_22_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_2_df_is_ws_24 <= io_in_r_bypass_22_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_2_stall_24 <= io_in_r_bypass_22_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_3_data_24 <= io_in_r_bypass_22_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_3_load_store_24 <= io_in_r_bypass_22_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_3_df_is_ws_24 <= io_in_r_bypass_22_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_3_stall_24 <= io_in_r_bypass_22_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_0_data_24 <= io_in_r_bypass_23_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_0_load_store_24 <= io_in_r_bypass_23_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_0_df_is_ws_24 <= io_in_r_bypass_23_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_0_stall_24 <= io_in_r_bypass_23_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_1_data_24 <= io_in_r_bypass_23_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_1_load_store_24 <= io_in_r_bypass_23_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_1_df_is_ws_24 <= io_in_r_bypass_23_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_1_stall_24 <= io_in_r_bypass_23_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_2_data_24 <= io_in_r_bypass_23_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_2_load_store_24 <= io_in_r_bypass_23_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_2_df_is_ws_24 <= io_in_r_bypass_23_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_2_stall_24 <= io_in_r_bypass_23_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_3_data_24 <= io_in_r_bypass_23_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_3_load_store_24 <= io_in_r_bypass_23_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_3_df_is_ws_24 <= io_in_r_bypass_23_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_3_stall_24 <= io_in_r_bypass_23_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_0_data_24 <= io_in_r_bypass_24_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_0_load_store_24 <= io_in_r_bypass_24_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_0_df_is_ws_24 <= io_in_r_bypass_24_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_0_stall_24 <= io_in_r_bypass_24_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_1_data_24 <= io_in_r_bypass_24_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_1_load_store_24 <= io_in_r_bypass_24_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_1_df_is_ws_24 <= io_in_r_bypass_24_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_1_stall_24 <= io_in_r_bypass_24_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_2_data_24 <= io_in_r_bypass_24_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_2_load_store_24 <= io_in_r_bypass_24_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_2_df_is_ws_24 <= io_in_r_bypass_24_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_2_stall_24 <= io_in_r_bypass_24_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_3_data_24 <= io_in_r_bypass_24_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_3_load_store_24 <= io_in_r_bypass_24_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_3_df_is_ws_24 <= io_in_r_bypass_24_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_3_stall_24 <= io_in_r_bypass_24_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_0_data_24 <= io_in_r_bypass_25_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_0_load_store_24 <= io_in_r_bypass_25_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_0_df_is_ws_24 <= io_in_r_bypass_25_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_0_stall_24 <= io_in_r_bypass_25_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_1_data_24 <= io_in_r_bypass_25_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_1_load_store_24 <= io_in_r_bypass_25_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_1_df_is_ws_24 <= io_in_r_bypass_25_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_1_stall_24 <= io_in_r_bypass_25_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_2_data_24 <= io_in_r_bypass_25_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_2_load_store_24 <= io_in_r_bypass_25_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_2_df_is_ws_24 <= io_in_r_bypass_25_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_2_stall_24 <= io_in_r_bypass_25_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_3_data_24 <= io_in_r_bypass_25_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_3_load_store_24 <= io_in_r_bypass_25_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_3_df_is_ws_24 <= io_in_r_bypass_25_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_3_stall_24 <= io_in_r_bypass_25_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_0_data_24 <= io_in_r_bypass_26_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_0_load_store_24 <= io_in_r_bypass_26_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_0_df_is_ws_24 <= io_in_r_bypass_26_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_0_stall_24 <= io_in_r_bypass_26_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_1_data_24 <= io_in_r_bypass_26_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_1_load_store_24 <= io_in_r_bypass_26_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_1_df_is_ws_24 <= io_in_r_bypass_26_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_1_stall_24 <= io_in_r_bypass_26_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_2_data_24 <= io_in_r_bypass_26_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_2_load_store_24 <= io_in_r_bypass_26_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_2_df_is_ws_24 <= io_in_r_bypass_26_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_2_stall_24 <= io_in_r_bypass_26_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_3_data_24 <= io_in_r_bypass_26_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_3_load_store_24 <= io_in_r_bypass_26_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_3_df_is_ws_24 <= io_in_r_bypass_26_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_3_stall_24 <= io_in_r_bypass_26_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_0_data_24 <= io_in_r_bypass_27_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_0_load_store_24 <= io_in_r_bypass_27_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_0_df_is_ws_24 <= io_in_r_bypass_27_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_0_stall_24 <= io_in_r_bypass_27_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_1_data_24 <= io_in_r_bypass_27_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_1_load_store_24 <= io_in_r_bypass_27_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_1_df_is_ws_24 <= io_in_r_bypass_27_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_1_stall_24 <= io_in_r_bypass_27_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_2_data_24 <= io_in_r_bypass_27_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_2_load_store_24 <= io_in_r_bypass_27_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_2_df_is_ws_24 <= io_in_r_bypass_27_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_2_stall_24 <= io_in_r_bypass_27_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_3_data_24 <= io_in_r_bypass_27_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_3_load_store_24 <= io_in_r_bypass_27_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_3_df_is_ws_24 <= io_in_r_bypass_27_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_3_stall_24 <= io_in_r_bypass_27_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_0_data_24 <= io_in_r_bypass_28_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_0_load_store_24 <= io_in_r_bypass_28_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_0_df_is_ws_24 <= io_in_r_bypass_28_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_0_stall_24 <= io_in_r_bypass_28_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_1_data_24 <= io_in_r_bypass_28_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_1_load_store_24 <= io_in_r_bypass_28_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_1_df_is_ws_24 <= io_in_r_bypass_28_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_1_stall_24 <= io_in_r_bypass_28_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_2_data_24 <= io_in_r_bypass_28_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_2_load_store_24 <= io_in_r_bypass_28_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_2_df_is_ws_24 <= io_in_r_bypass_28_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_2_stall_24 <= io_in_r_bypass_28_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_3_data_24 <= io_in_r_bypass_28_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_3_load_store_24 <= io_in_r_bypass_28_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_3_df_is_ws_24 <= io_in_r_bypass_28_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_3_stall_24 <= io_in_r_bypass_28_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_0_data_24 <= io_in_r_bypass_29_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_0_load_store_24 <= io_in_r_bypass_29_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_0_df_is_ws_24 <= io_in_r_bypass_29_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_0_stall_24 <= io_in_r_bypass_29_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_1_data_24 <= io_in_r_bypass_29_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_1_load_store_24 <= io_in_r_bypass_29_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_1_df_is_ws_24 <= io_in_r_bypass_29_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_1_stall_24 <= io_in_r_bypass_29_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_2_data_24 <= io_in_r_bypass_29_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_2_load_store_24 <= io_in_r_bypass_29_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_2_df_is_ws_24 <= io_in_r_bypass_29_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_2_stall_24 <= io_in_r_bypass_29_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_3_data_24 <= io_in_r_bypass_29_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_3_load_store_24 <= io_in_r_bypass_29_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_3_df_is_ws_24 <= io_in_r_bypass_29_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_3_stall_24 <= io_in_r_bypass_29_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_0_data_24 <= io_in_r_bypass_30_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_0_load_store_24 <= io_in_r_bypass_30_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_0_df_is_ws_24 <= io_in_r_bypass_30_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_0_stall_24 <= io_in_r_bypass_30_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_1_data_24 <= io_in_r_bypass_30_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_1_load_store_24 <= io_in_r_bypass_30_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_1_df_is_ws_24 <= io_in_r_bypass_30_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_1_stall_24 <= io_in_r_bypass_30_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_2_data_24 <= io_in_r_bypass_30_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_2_load_store_24 <= io_in_r_bypass_30_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_2_df_is_ws_24 <= io_in_r_bypass_30_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_2_stall_24 <= io_in_r_bypass_30_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_3_data_24 <= io_in_r_bypass_30_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_3_load_store_24 <= io_in_r_bypass_30_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_3_df_is_ws_24 <= io_in_r_bypass_30_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_3_stall_24 <= io_in_r_bypass_30_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_0_data_24 <= io_in_r_bypass_31_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_0_load_store_24 <= io_in_r_bypass_31_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_0_df_is_ws_24 <= io_in_r_bypass_31_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_0_stall_24 <= io_in_r_bypass_31_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_1_data_24 <= io_in_r_bypass_31_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_1_load_store_24 <= io_in_r_bypass_31_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_1_df_is_ws_24 <= io_in_r_bypass_31_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_1_stall_24 <= io_in_r_bypass_31_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_2_data_24 <= io_in_r_bypass_31_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_2_load_store_24 <= io_in_r_bypass_31_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_2_df_is_ws_24 <= io_in_r_bypass_31_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_2_stall_24 <= io_in_r_bypass_31_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_3_data_24 <= io_in_r_bypass_31_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_3_load_store_24 <= io_in_r_bypass_31_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_3_df_is_ws_24 <= io_in_r_bypass_31_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_3_stall_24 <= io_in_r_bypass_31_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_0_data_25 <= io_in_r_bypass_0_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_0_load_store_25 <= io_in_r_bypass_0_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_0_df_is_ws_25 <= io_in_r_bypass_0_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_0_stall_25 <= io_in_r_bypass_0_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_1_data_25 <= io_in_r_bypass_0_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_1_load_store_25 <= io_in_r_bypass_0_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_1_df_is_ws_25 <= io_in_r_bypass_0_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_1_stall_25 <= io_in_r_bypass_0_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_2_data_25 <= io_in_r_bypass_0_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_2_load_store_25 <= io_in_r_bypass_0_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_2_df_is_ws_25 <= io_in_r_bypass_0_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_2_stall_25 <= io_in_r_bypass_0_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_3_data_25 <= io_in_r_bypass_0_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_3_load_store_25 <= io_in_r_bypass_0_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_3_df_is_ws_25 <= io_in_r_bypass_0_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_3_stall_25 <= io_in_r_bypass_0_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_0_data_25 <= io_in_r_bypass_1_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_0_load_store_25 <= io_in_r_bypass_1_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_0_df_is_ws_25 <= io_in_r_bypass_1_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_0_stall_25 <= io_in_r_bypass_1_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_1_data_25 <= io_in_r_bypass_1_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_1_load_store_25 <= io_in_r_bypass_1_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_1_df_is_ws_25 <= io_in_r_bypass_1_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_1_stall_25 <= io_in_r_bypass_1_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_2_data_25 <= io_in_r_bypass_1_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_2_load_store_25 <= io_in_r_bypass_1_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_2_df_is_ws_25 <= io_in_r_bypass_1_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_2_stall_25 <= io_in_r_bypass_1_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_3_data_25 <= io_in_r_bypass_1_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_3_load_store_25 <= io_in_r_bypass_1_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_3_df_is_ws_25 <= io_in_r_bypass_1_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_3_stall_25 <= io_in_r_bypass_1_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_0_data_25 <= io_in_r_bypass_2_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_0_load_store_25 <= io_in_r_bypass_2_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_0_df_is_ws_25 <= io_in_r_bypass_2_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_0_stall_25 <= io_in_r_bypass_2_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_1_data_25 <= io_in_r_bypass_2_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_1_load_store_25 <= io_in_r_bypass_2_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_1_df_is_ws_25 <= io_in_r_bypass_2_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_1_stall_25 <= io_in_r_bypass_2_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_2_data_25 <= io_in_r_bypass_2_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_2_load_store_25 <= io_in_r_bypass_2_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_2_df_is_ws_25 <= io_in_r_bypass_2_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_2_stall_25 <= io_in_r_bypass_2_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_3_data_25 <= io_in_r_bypass_2_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_3_load_store_25 <= io_in_r_bypass_2_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_3_df_is_ws_25 <= io_in_r_bypass_2_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_3_stall_25 <= io_in_r_bypass_2_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_0_data_25 <= io_in_r_bypass_3_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_0_load_store_25 <= io_in_r_bypass_3_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_0_df_is_ws_25 <= io_in_r_bypass_3_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_0_stall_25 <= io_in_r_bypass_3_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_1_data_25 <= io_in_r_bypass_3_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_1_load_store_25 <= io_in_r_bypass_3_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_1_df_is_ws_25 <= io_in_r_bypass_3_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_1_stall_25 <= io_in_r_bypass_3_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_2_data_25 <= io_in_r_bypass_3_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_2_load_store_25 <= io_in_r_bypass_3_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_2_df_is_ws_25 <= io_in_r_bypass_3_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_2_stall_25 <= io_in_r_bypass_3_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_3_data_25 <= io_in_r_bypass_3_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_3_load_store_25 <= io_in_r_bypass_3_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_3_df_is_ws_25 <= io_in_r_bypass_3_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_3_stall_25 <= io_in_r_bypass_3_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_0_data_25 <= io_in_r_bypass_4_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_0_load_store_25 <= io_in_r_bypass_4_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_0_df_is_ws_25 <= io_in_r_bypass_4_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_0_stall_25 <= io_in_r_bypass_4_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_1_data_25 <= io_in_r_bypass_4_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_1_load_store_25 <= io_in_r_bypass_4_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_1_df_is_ws_25 <= io_in_r_bypass_4_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_1_stall_25 <= io_in_r_bypass_4_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_2_data_25 <= io_in_r_bypass_4_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_2_load_store_25 <= io_in_r_bypass_4_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_2_df_is_ws_25 <= io_in_r_bypass_4_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_2_stall_25 <= io_in_r_bypass_4_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_3_data_25 <= io_in_r_bypass_4_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_3_load_store_25 <= io_in_r_bypass_4_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_3_df_is_ws_25 <= io_in_r_bypass_4_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_3_stall_25 <= io_in_r_bypass_4_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_0_data_25 <= io_in_r_bypass_5_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_0_load_store_25 <= io_in_r_bypass_5_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_0_df_is_ws_25 <= io_in_r_bypass_5_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_0_stall_25 <= io_in_r_bypass_5_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_1_data_25 <= io_in_r_bypass_5_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_1_load_store_25 <= io_in_r_bypass_5_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_1_df_is_ws_25 <= io_in_r_bypass_5_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_1_stall_25 <= io_in_r_bypass_5_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_2_data_25 <= io_in_r_bypass_5_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_2_load_store_25 <= io_in_r_bypass_5_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_2_df_is_ws_25 <= io_in_r_bypass_5_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_2_stall_25 <= io_in_r_bypass_5_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_3_data_25 <= io_in_r_bypass_5_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_3_load_store_25 <= io_in_r_bypass_5_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_3_df_is_ws_25 <= io_in_r_bypass_5_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_3_stall_25 <= io_in_r_bypass_5_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_0_data_25 <= io_in_r_bypass_6_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_0_load_store_25 <= io_in_r_bypass_6_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_0_df_is_ws_25 <= io_in_r_bypass_6_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_0_stall_25 <= io_in_r_bypass_6_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_1_data_25 <= io_in_r_bypass_6_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_1_load_store_25 <= io_in_r_bypass_6_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_1_df_is_ws_25 <= io_in_r_bypass_6_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_1_stall_25 <= io_in_r_bypass_6_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_2_data_25 <= io_in_r_bypass_6_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_2_load_store_25 <= io_in_r_bypass_6_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_2_df_is_ws_25 <= io_in_r_bypass_6_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_2_stall_25 <= io_in_r_bypass_6_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_3_data_25 <= io_in_r_bypass_6_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_3_load_store_25 <= io_in_r_bypass_6_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_3_df_is_ws_25 <= io_in_r_bypass_6_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_3_stall_25 <= io_in_r_bypass_6_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_0_data_25 <= io_in_r_bypass_7_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_0_load_store_25 <= io_in_r_bypass_7_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_0_df_is_ws_25 <= io_in_r_bypass_7_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_0_stall_25 <= io_in_r_bypass_7_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_1_data_25 <= io_in_r_bypass_7_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_1_load_store_25 <= io_in_r_bypass_7_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_1_df_is_ws_25 <= io_in_r_bypass_7_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_1_stall_25 <= io_in_r_bypass_7_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_2_data_25 <= io_in_r_bypass_7_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_2_load_store_25 <= io_in_r_bypass_7_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_2_df_is_ws_25 <= io_in_r_bypass_7_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_2_stall_25 <= io_in_r_bypass_7_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_3_data_25 <= io_in_r_bypass_7_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_3_load_store_25 <= io_in_r_bypass_7_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_3_df_is_ws_25 <= io_in_r_bypass_7_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_3_stall_25 <= io_in_r_bypass_7_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_0_data_25 <= io_in_r_bypass_8_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_0_load_store_25 <= io_in_r_bypass_8_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_0_df_is_ws_25 <= io_in_r_bypass_8_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_0_stall_25 <= io_in_r_bypass_8_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_1_data_25 <= io_in_r_bypass_8_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_1_load_store_25 <= io_in_r_bypass_8_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_1_df_is_ws_25 <= io_in_r_bypass_8_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_1_stall_25 <= io_in_r_bypass_8_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_2_data_25 <= io_in_r_bypass_8_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_2_load_store_25 <= io_in_r_bypass_8_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_2_df_is_ws_25 <= io_in_r_bypass_8_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_2_stall_25 <= io_in_r_bypass_8_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_3_data_25 <= io_in_r_bypass_8_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_3_load_store_25 <= io_in_r_bypass_8_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_3_df_is_ws_25 <= io_in_r_bypass_8_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_3_stall_25 <= io_in_r_bypass_8_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_0_data_25 <= io_in_r_bypass_9_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_0_load_store_25 <= io_in_r_bypass_9_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_0_df_is_ws_25 <= io_in_r_bypass_9_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_0_stall_25 <= io_in_r_bypass_9_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_1_data_25 <= io_in_r_bypass_9_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_1_load_store_25 <= io_in_r_bypass_9_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_1_df_is_ws_25 <= io_in_r_bypass_9_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_1_stall_25 <= io_in_r_bypass_9_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_2_data_25 <= io_in_r_bypass_9_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_2_load_store_25 <= io_in_r_bypass_9_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_2_df_is_ws_25 <= io_in_r_bypass_9_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_2_stall_25 <= io_in_r_bypass_9_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_3_data_25 <= io_in_r_bypass_9_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_3_load_store_25 <= io_in_r_bypass_9_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_3_df_is_ws_25 <= io_in_r_bypass_9_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_3_stall_25 <= io_in_r_bypass_9_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_0_data_25 <= io_in_r_bypass_10_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_0_load_store_25 <= io_in_r_bypass_10_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_0_df_is_ws_25 <= io_in_r_bypass_10_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_0_stall_25 <= io_in_r_bypass_10_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_1_data_25 <= io_in_r_bypass_10_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_1_load_store_25 <= io_in_r_bypass_10_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_1_df_is_ws_25 <= io_in_r_bypass_10_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_1_stall_25 <= io_in_r_bypass_10_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_2_data_25 <= io_in_r_bypass_10_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_2_load_store_25 <= io_in_r_bypass_10_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_2_df_is_ws_25 <= io_in_r_bypass_10_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_2_stall_25 <= io_in_r_bypass_10_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_3_data_25 <= io_in_r_bypass_10_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_3_load_store_25 <= io_in_r_bypass_10_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_3_df_is_ws_25 <= io_in_r_bypass_10_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_3_stall_25 <= io_in_r_bypass_10_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_0_data_25 <= io_in_r_bypass_11_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_0_load_store_25 <= io_in_r_bypass_11_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_0_df_is_ws_25 <= io_in_r_bypass_11_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_0_stall_25 <= io_in_r_bypass_11_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_1_data_25 <= io_in_r_bypass_11_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_1_load_store_25 <= io_in_r_bypass_11_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_1_df_is_ws_25 <= io_in_r_bypass_11_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_1_stall_25 <= io_in_r_bypass_11_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_2_data_25 <= io_in_r_bypass_11_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_2_load_store_25 <= io_in_r_bypass_11_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_2_df_is_ws_25 <= io_in_r_bypass_11_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_2_stall_25 <= io_in_r_bypass_11_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_3_data_25 <= io_in_r_bypass_11_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_3_load_store_25 <= io_in_r_bypass_11_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_3_df_is_ws_25 <= io_in_r_bypass_11_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_3_stall_25 <= io_in_r_bypass_11_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_0_data_25 <= io_in_r_bypass_12_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_0_load_store_25 <= io_in_r_bypass_12_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_0_df_is_ws_25 <= io_in_r_bypass_12_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_0_stall_25 <= io_in_r_bypass_12_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_1_data_25 <= io_in_r_bypass_12_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_1_load_store_25 <= io_in_r_bypass_12_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_1_df_is_ws_25 <= io_in_r_bypass_12_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_1_stall_25 <= io_in_r_bypass_12_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_2_data_25 <= io_in_r_bypass_12_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_2_load_store_25 <= io_in_r_bypass_12_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_2_df_is_ws_25 <= io_in_r_bypass_12_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_2_stall_25 <= io_in_r_bypass_12_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_3_data_25 <= io_in_r_bypass_12_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_3_load_store_25 <= io_in_r_bypass_12_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_3_df_is_ws_25 <= io_in_r_bypass_12_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_3_stall_25 <= io_in_r_bypass_12_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_0_data_25 <= io_in_r_bypass_13_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_0_load_store_25 <= io_in_r_bypass_13_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_0_df_is_ws_25 <= io_in_r_bypass_13_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_0_stall_25 <= io_in_r_bypass_13_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_1_data_25 <= io_in_r_bypass_13_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_1_load_store_25 <= io_in_r_bypass_13_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_1_df_is_ws_25 <= io_in_r_bypass_13_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_1_stall_25 <= io_in_r_bypass_13_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_2_data_25 <= io_in_r_bypass_13_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_2_load_store_25 <= io_in_r_bypass_13_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_2_df_is_ws_25 <= io_in_r_bypass_13_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_2_stall_25 <= io_in_r_bypass_13_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_3_data_25 <= io_in_r_bypass_13_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_3_load_store_25 <= io_in_r_bypass_13_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_3_df_is_ws_25 <= io_in_r_bypass_13_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_3_stall_25 <= io_in_r_bypass_13_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_0_data_25 <= io_in_r_bypass_14_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_0_load_store_25 <= io_in_r_bypass_14_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_0_df_is_ws_25 <= io_in_r_bypass_14_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_0_stall_25 <= io_in_r_bypass_14_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_1_data_25 <= io_in_r_bypass_14_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_1_load_store_25 <= io_in_r_bypass_14_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_1_df_is_ws_25 <= io_in_r_bypass_14_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_1_stall_25 <= io_in_r_bypass_14_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_2_data_25 <= io_in_r_bypass_14_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_2_load_store_25 <= io_in_r_bypass_14_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_2_df_is_ws_25 <= io_in_r_bypass_14_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_2_stall_25 <= io_in_r_bypass_14_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_3_data_25 <= io_in_r_bypass_14_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_3_load_store_25 <= io_in_r_bypass_14_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_3_df_is_ws_25 <= io_in_r_bypass_14_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_3_stall_25 <= io_in_r_bypass_14_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_0_data_25 <= io_in_r_bypass_15_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_0_load_store_25 <= io_in_r_bypass_15_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_0_df_is_ws_25 <= io_in_r_bypass_15_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_0_stall_25 <= io_in_r_bypass_15_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_1_data_25 <= io_in_r_bypass_15_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_1_load_store_25 <= io_in_r_bypass_15_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_1_df_is_ws_25 <= io_in_r_bypass_15_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_1_stall_25 <= io_in_r_bypass_15_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_2_data_25 <= io_in_r_bypass_15_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_2_load_store_25 <= io_in_r_bypass_15_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_2_df_is_ws_25 <= io_in_r_bypass_15_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_2_stall_25 <= io_in_r_bypass_15_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_3_data_25 <= io_in_r_bypass_15_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_3_load_store_25 <= io_in_r_bypass_15_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_3_df_is_ws_25 <= io_in_r_bypass_15_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_3_stall_25 <= io_in_r_bypass_15_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_0_data_25 <= io_in_r_bypass_16_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_0_load_store_25 <= io_in_r_bypass_16_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_0_df_is_ws_25 <= io_in_r_bypass_16_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_0_stall_25 <= io_in_r_bypass_16_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_1_data_25 <= io_in_r_bypass_16_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_1_load_store_25 <= io_in_r_bypass_16_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_1_df_is_ws_25 <= io_in_r_bypass_16_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_1_stall_25 <= io_in_r_bypass_16_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_2_data_25 <= io_in_r_bypass_16_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_2_load_store_25 <= io_in_r_bypass_16_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_2_df_is_ws_25 <= io_in_r_bypass_16_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_2_stall_25 <= io_in_r_bypass_16_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_3_data_25 <= io_in_r_bypass_16_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_3_load_store_25 <= io_in_r_bypass_16_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_3_df_is_ws_25 <= io_in_r_bypass_16_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_3_stall_25 <= io_in_r_bypass_16_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_0_data_25 <= io_in_r_bypass_17_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_0_load_store_25 <= io_in_r_bypass_17_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_0_df_is_ws_25 <= io_in_r_bypass_17_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_0_stall_25 <= io_in_r_bypass_17_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_1_data_25 <= io_in_r_bypass_17_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_1_load_store_25 <= io_in_r_bypass_17_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_1_df_is_ws_25 <= io_in_r_bypass_17_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_1_stall_25 <= io_in_r_bypass_17_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_2_data_25 <= io_in_r_bypass_17_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_2_load_store_25 <= io_in_r_bypass_17_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_2_df_is_ws_25 <= io_in_r_bypass_17_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_2_stall_25 <= io_in_r_bypass_17_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_3_data_25 <= io_in_r_bypass_17_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_3_load_store_25 <= io_in_r_bypass_17_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_3_df_is_ws_25 <= io_in_r_bypass_17_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_3_stall_25 <= io_in_r_bypass_17_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_0_data_25 <= io_in_r_bypass_18_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_0_load_store_25 <= io_in_r_bypass_18_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_0_df_is_ws_25 <= io_in_r_bypass_18_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_0_stall_25 <= io_in_r_bypass_18_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_1_data_25 <= io_in_r_bypass_18_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_1_load_store_25 <= io_in_r_bypass_18_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_1_df_is_ws_25 <= io_in_r_bypass_18_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_1_stall_25 <= io_in_r_bypass_18_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_2_data_25 <= io_in_r_bypass_18_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_2_load_store_25 <= io_in_r_bypass_18_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_2_df_is_ws_25 <= io_in_r_bypass_18_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_2_stall_25 <= io_in_r_bypass_18_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_3_data_25 <= io_in_r_bypass_18_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_3_load_store_25 <= io_in_r_bypass_18_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_3_df_is_ws_25 <= io_in_r_bypass_18_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_3_stall_25 <= io_in_r_bypass_18_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_0_data_25 <= io_in_r_bypass_19_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_0_load_store_25 <= io_in_r_bypass_19_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_0_df_is_ws_25 <= io_in_r_bypass_19_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_0_stall_25 <= io_in_r_bypass_19_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_1_data_25 <= io_in_r_bypass_19_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_1_load_store_25 <= io_in_r_bypass_19_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_1_df_is_ws_25 <= io_in_r_bypass_19_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_1_stall_25 <= io_in_r_bypass_19_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_2_data_25 <= io_in_r_bypass_19_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_2_load_store_25 <= io_in_r_bypass_19_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_2_df_is_ws_25 <= io_in_r_bypass_19_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_2_stall_25 <= io_in_r_bypass_19_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_3_data_25 <= io_in_r_bypass_19_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_3_load_store_25 <= io_in_r_bypass_19_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_3_df_is_ws_25 <= io_in_r_bypass_19_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_3_stall_25 <= io_in_r_bypass_19_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_0_data_25 <= io_in_r_bypass_20_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_0_load_store_25 <= io_in_r_bypass_20_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_0_df_is_ws_25 <= io_in_r_bypass_20_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_0_stall_25 <= io_in_r_bypass_20_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_1_data_25 <= io_in_r_bypass_20_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_1_load_store_25 <= io_in_r_bypass_20_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_1_df_is_ws_25 <= io_in_r_bypass_20_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_1_stall_25 <= io_in_r_bypass_20_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_2_data_25 <= io_in_r_bypass_20_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_2_load_store_25 <= io_in_r_bypass_20_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_2_df_is_ws_25 <= io_in_r_bypass_20_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_2_stall_25 <= io_in_r_bypass_20_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_3_data_25 <= io_in_r_bypass_20_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_3_load_store_25 <= io_in_r_bypass_20_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_3_df_is_ws_25 <= io_in_r_bypass_20_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_3_stall_25 <= io_in_r_bypass_20_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_0_data_25 <= io_in_r_bypass_21_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_0_load_store_25 <= io_in_r_bypass_21_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_0_df_is_ws_25 <= io_in_r_bypass_21_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_0_stall_25 <= io_in_r_bypass_21_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_1_data_25 <= io_in_r_bypass_21_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_1_load_store_25 <= io_in_r_bypass_21_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_1_df_is_ws_25 <= io_in_r_bypass_21_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_1_stall_25 <= io_in_r_bypass_21_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_2_data_25 <= io_in_r_bypass_21_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_2_load_store_25 <= io_in_r_bypass_21_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_2_df_is_ws_25 <= io_in_r_bypass_21_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_2_stall_25 <= io_in_r_bypass_21_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_3_data_25 <= io_in_r_bypass_21_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_3_load_store_25 <= io_in_r_bypass_21_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_3_df_is_ws_25 <= io_in_r_bypass_21_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_3_stall_25 <= io_in_r_bypass_21_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_0_data_25 <= io_in_r_bypass_22_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_0_load_store_25 <= io_in_r_bypass_22_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_0_df_is_ws_25 <= io_in_r_bypass_22_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_0_stall_25 <= io_in_r_bypass_22_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_1_data_25 <= io_in_r_bypass_22_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_1_load_store_25 <= io_in_r_bypass_22_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_1_df_is_ws_25 <= io_in_r_bypass_22_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_1_stall_25 <= io_in_r_bypass_22_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_2_data_25 <= io_in_r_bypass_22_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_2_load_store_25 <= io_in_r_bypass_22_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_2_df_is_ws_25 <= io_in_r_bypass_22_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_2_stall_25 <= io_in_r_bypass_22_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_3_data_25 <= io_in_r_bypass_22_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_3_load_store_25 <= io_in_r_bypass_22_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_3_df_is_ws_25 <= io_in_r_bypass_22_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_3_stall_25 <= io_in_r_bypass_22_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_0_data_25 <= io_in_r_bypass_23_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_0_load_store_25 <= io_in_r_bypass_23_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_0_df_is_ws_25 <= io_in_r_bypass_23_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_0_stall_25 <= io_in_r_bypass_23_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_1_data_25 <= io_in_r_bypass_23_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_1_load_store_25 <= io_in_r_bypass_23_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_1_df_is_ws_25 <= io_in_r_bypass_23_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_1_stall_25 <= io_in_r_bypass_23_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_2_data_25 <= io_in_r_bypass_23_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_2_load_store_25 <= io_in_r_bypass_23_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_2_df_is_ws_25 <= io_in_r_bypass_23_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_2_stall_25 <= io_in_r_bypass_23_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_3_data_25 <= io_in_r_bypass_23_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_3_load_store_25 <= io_in_r_bypass_23_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_3_df_is_ws_25 <= io_in_r_bypass_23_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_3_stall_25 <= io_in_r_bypass_23_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_0_data_25 <= io_in_r_bypass_24_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_0_load_store_25 <= io_in_r_bypass_24_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_0_df_is_ws_25 <= io_in_r_bypass_24_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_0_stall_25 <= io_in_r_bypass_24_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_1_data_25 <= io_in_r_bypass_24_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_1_load_store_25 <= io_in_r_bypass_24_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_1_df_is_ws_25 <= io_in_r_bypass_24_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_1_stall_25 <= io_in_r_bypass_24_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_2_data_25 <= io_in_r_bypass_24_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_2_load_store_25 <= io_in_r_bypass_24_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_2_df_is_ws_25 <= io_in_r_bypass_24_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_2_stall_25 <= io_in_r_bypass_24_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_3_data_25 <= io_in_r_bypass_24_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_3_load_store_25 <= io_in_r_bypass_24_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_3_df_is_ws_25 <= io_in_r_bypass_24_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_3_stall_25 <= io_in_r_bypass_24_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_0_data_25 <= io_in_r_bypass_25_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_0_load_store_25 <= io_in_r_bypass_25_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_0_df_is_ws_25 <= io_in_r_bypass_25_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_0_stall_25 <= io_in_r_bypass_25_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_1_data_25 <= io_in_r_bypass_25_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_1_load_store_25 <= io_in_r_bypass_25_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_1_df_is_ws_25 <= io_in_r_bypass_25_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_1_stall_25 <= io_in_r_bypass_25_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_2_data_25 <= io_in_r_bypass_25_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_2_load_store_25 <= io_in_r_bypass_25_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_2_df_is_ws_25 <= io_in_r_bypass_25_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_2_stall_25 <= io_in_r_bypass_25_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_3_data_25 <= io_in_r_bypass_25_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_3_load_store_25 <= io_in_r_bypass_25_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_3_df_is_ws_25 <= io_in_r_bypass_25_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_3_stall_25 <= io_in_r_bypass_25_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_0_data_25 <= io_in_r_bypass_26_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_0_load_store_25 <= io_in_r_bypass_26_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_0_df_is_ws_25 <= io_in_r_bypass_26_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_0_stall_25 <= io_in_r_bypass_26_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_1_data_25 <= io_in_r_bypass_26_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_1_load_store_25 <= io_in_r_bypass_26_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_1_df_is_ws_25 <= io_in_r_bypass_26_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_1_stall_25 <= io_in_r_bypass_26_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_2_data_25 <= io_in_r_bypass_26_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_2_load_store_25 <= io_in_r_bypass_26_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_2_df_is_ws_25 <= io_in_r_bypass_26_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_2_stall_25 <= io_in_r_bypass_26_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_3_data_25 <= io_in_r_bypass_26_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_3_load_store_25 <= io_in_r_bypass_26_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_3_df_is_ws_25 <= io_in_r_bypass_26_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_3_stall_25 <= io_in_r_bypass_26_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_0_data_25 <= io_in_r_bypass_27_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_0_load_store_25 <= io_in_r_bypass_27_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_0_df_is_ws_25 <= io_in_r_bypass_27_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_0_stall_25 <= io_in_r_bypass_27_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_1_data_25 <= io_in_r_bypass_27_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_1_load_store_25 <= io_in_r_bypass_27_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_1_df_is_ws_25 <= io_in_r_bypass_27_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_1_stall_25 <= io_in_r_bypass_27_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_2_data_25 <= io_in_r_bypass_27_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_2_load_store_25 <= io_in_r_bypass_27_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_2_df_is_ws_25 <= io_in_r_bypass_27_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_2_stall_25 <= io_in_r_bypass_27_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_3_data_25 <= io_in_r_bypass_27_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_3_load_store_25 <= io_in_r_bypass_27_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_3_df_is_ws_25 <= io_in_r_bypass_27_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_3_stall_25 <= io_in_r_bypass_27_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_0_data_25 <= io_in_r_bypass_28_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_0_load_store_25 <= io_in_r_bypass_28_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_0_df_is_ws_25 <= io_in_r_bypass_28_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_0_stall_25 <= io_in_r_bypass_28_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_1_data_25 <= io_in_r_bypass_28_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_1_load_store_25 <= io_in_r_bypass_28_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_1_df_is_ws_25 <= io_in_r_bypass_28_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_1_stall_25 <= io_in_r_bypass_28_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_2_data_25 <= io_in_r_bypass_28_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_2_load_store_25 <= io_in_r_bypass_28_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_2_df_is_ws_25 <= io_in_r_bypass_28_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_2_stall_25 <= io_in_r_bypass_28_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_3_data_25 <= io_in_r_bypass_28_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_3_load_store_25 <= io_in_r_bypass_28_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_3_df_is_ws_25 <= io_in_r_bypass_28_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_3_stall_25 <= io_in_r_bypass_28_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_0_data_25 <= io_in_r_bypass_29_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_0_load_store_25 <= io_in_r_bypass_29_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_0_df_is_ws_25 <= io_in_r_bypass_29_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_0_stall_25 <= io_in_r_bypass_29_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_1_data_25 <= io_in_r_bypass_29_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_1_load_store_25 <= io_in_r_bypass_29_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_1_df_is_ws_25 <= io_in_r_bypass_29_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_1_stall_25 <= io_in_r_bypass_29_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_2_data_25 <= io_in_r_bypass_29_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_2_load_store_25 <= io_in_r_bypass_29_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_2_df_is_ws_25 <= io_in_r_bypass_29_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_2_stall_25 <= io_in_r_bypass_29_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_3_data_25 <= io_in_r_bypass_29_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_3_load_store_25 <= io_in_r_bypass_29_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_3_df_is_ws_25 <= io_in_r_bypass_29_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_3_stall_25 <= io_in_r_bypass_29_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_0_data_25 <= io_in_r_bypass_30_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_0_load_store_25 <= io_in_r_bypass_30_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_0_df_is_ws_25 <= io_in_r_bypass_30_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_0_stall_25 <= io_in_r_bypass_30_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_1_data_25 <= io_in_r_bypass_30_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_1_load_store_25 <= io_in_r_bypass_30_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_1_df_is_ws_25 <= io_in_r_bypass_30_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_1_stall_25 <= io_in_r_bypass_30_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_2_data_25 <= io_in_r_bypass_30_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_2_load_store_25 <= io_in_r_bypass_30_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_2_df_is_ws_25 <= io_in_r_bypass_30_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_2_stall_25 <= io_in_r_bypass_30_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_3_data_25 <= io_in_r_bypass_30_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_3_load_store_25 <= io_in_r_bypass_30_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_3_df_is_ws_25 <= io_in_r_bypass_30_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_3_stall_25 <= io_in_r_bypass_30_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_0_data_25 <= io_in_r_bypass_31_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_0_load_store_25 <= io_in_r_bypass_31_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_0_df_is_ws_25 <= io_in_r_bypass_31_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_0_stall_25 <= io_in_r_bypass_31_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_1_data_25 <= io_in_r_bypass_31_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_1_load_store_25 <= io_in_r_bypass_31_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_1_df_is_ws_25 <= io_in_r_bypass_31_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_1_stall_25 <= io_in_r_bypass_31_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_2_data_25 <= io_in_r_bypass_31_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_2_load_store_25 <= io_in_r_bypass_31_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_2_df_is_ws_25 <= io_in_r_bypass_31_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_2_stall_25 <= io_in_r_bypass_31_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_3_data_25 <= io_in_r_bypass_31_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_3_load_store_25 <= io_in_r_bypass_31_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_3_df_is_ws_25 <= io_in_r_bypass_31_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_3_stall_25 <= io_in_r_bypass_31_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_0_data_26 <= io_in_r_bypass_0_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_0_load_store_26 <= io_in_r_bypass_0_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_0_df_is_ws_26 <= io_in_r_bypass_0_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_0_stall_26 <= io_in_r_bypass_0_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_1_data_26 <= io_in_r_bypass_0_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_1_load_store_26 <= io_in_r_bypass_0_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_1_df_is_ws_26 <= io_in_r_bypass_0_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_1_stall_26 <= io_in_r_bypass_0_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_2_data_26 <= io_in_r_bypass_0_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_2_load_store_26 <= io_in_r_bypass_0_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_2_df_is_ws_26 <= io_in_r_bypass_0_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_2_stall_26 <= io_in_r_bypass_0_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_3_data_26 <= io_in_r_bypass_0_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_3_load_store_26 <= io_in_r_bypass_0_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_3_df_is_ws_26 <= io_in_r_bypass_0_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_3_stall_26 <= io_in_r_bypass_0_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_0_data_26 <= io_in_r_bypass_1_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_0_load_store_26 <= io_in_r_bypass_1_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_0_df_is_ws_26 <= io_in_r_bypass_1_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_0_stall_26 <= io_in_r_bypass_1_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_1_data_26 <= io_in_r_bypass_1_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_1_load_store_26 <= io_in_r_bypass_1_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_1_df_is_ws_26 <= io_in_r_bypass_1_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_1_stall_26 <= io_in_r_bypass_1_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_2_data_26 <= io_in_r_bypass_1_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_2_load_store_26 <= io_in_r_bypass_1_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_2_df_is_ws_26 <= io_in_r_bypass_1_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_2_stall_26 <= io_in_r_bypass_1_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_3_data_26 <= io_in_r_bypass_1_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_3_load_store_26 <= io_in_r_bypass_1_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_3_df_is_ws_26 <= io_in_r_bypass_1_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_3_stall_26 <= io_in_r_bypass_1_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_0_data_26 <= io_in_r_bypass_2_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_0_load_store_26 <= io_in_r_bypass_2_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_0_df_is_ws_26 <= io_in_r_bypass_2_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_0_stall_26 <= io_in_r_bypass_2_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_1_data_26 <= io_in_r_bypass_2_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_1_load_store_26 <= io_in_r_bypass_2_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_1_df_is_ws_26 <= io_in_r_bypass_2_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_1_stall_26 <= io_in_r_bypass_2_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_2_data_26 <= io_in_r_bypass_2_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_2_load_store_26 <= io_in_r_bypass_2_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_2_df_is_ws_26 <= io_in_r_bypass_2_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_2_stall_26 <= io_in_r_bypass_2_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_3_data_26 <= io_in_r_bypass_2_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_3_load_store_26 <= io_in_r_bypass_2_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_3_df_is_ws_26 <= io_in_r_bypass_2_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_3_stall_26 <= io_in_r_bypass_2_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_0_data_26 <= io_in_r_bypass_3_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_0_load_store_26 <= io_in_r_bypass_3_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_0_df_is_ws_26 <= io_in_r_bypass_3_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_0_stall_26 <= io_in_r_bypass_3_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_1_data_26 <= io_in_r_bypass_3_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_1_load_store_26 <= io_in_r_bypass_3_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_1_df_is_ws_26 <= io_in_r_bypass_3_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_1_stall_26 <= io_in_r_bypass_3_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_2_data_26 <= io_in_r_bypass_3_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_2_load_store_26 <= io_in_r_bypass_3_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_2_df_is_ws_26 <= io_in_r_bypass_3_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_2_stall_26 <= io_in_r_bypass_3_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_3_data_26 <= io_in_r_bypass_3_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_3_load_store_26 <= io_in_r_bypass_3_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_3_df_is_ws_26 <= io_in_r_bypass_3_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_3_stall_26 <= io_in_r_bypass_3_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_0_data_26 <= io_in_r_bypass_4_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_0_load_store_26 <= io_in_r_bypass_4_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_0_df_is_ws_26 <= io_in_r_bypass_4_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_0_stall_26 <= io_in_r_bypass_4_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_1_data_26 <= io_in_r_bypass_4_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_1_load_store_26 <= io_in_r_bypass_4_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_1_df_is_ws_26 <= io_in_r_bypass_4_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_1_stall_26 <= io_in_r_bypass_4_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_2_data_26 <= io_in_r_bypass_4_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_2_load_store_26 <= io_in_r_bypass_4_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_2_df_is_ws_26 <= io_in_r_bypass_4_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_2_stall_26 <= io_in_r_bypass_4_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_3_data_26 <= io_in_r_bypass_4_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_3_load_store_26 <= io_in_r_bypass_4_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_3_df_is_ws_26 <= io_in_r_bypass_4_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_3_stall_26 <= io_in_r_bypass_4_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_0_data_26 <= io_in_r_bypass_5_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_0_load_store_26 <= io_in_r_bypass_5_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_0_df_is_ws_26 <= io_in_r_bypass_5_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_0_stall_26 <= io_in_r_bypass_5_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_1_data_26 <= io_in_r_bypass_5_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_1_load_store_26 <= io_in_r_bypass_5_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_1_df_is_ws_26 <= io_in_r_bypass_5_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_1_stall_26 <= io_in_r_bypass_5_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_2_data_26 <= io_in_r_bypass_5_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_2_load_store_26 <= io_in_r_bypass_5_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_2_df_is_ws_26 <= io_in_r_bypass_5_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_2_stall_26 <= io_in_r_bypass_5_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_3_data_26 <= io_in_r_bypass_5_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_3_load_store_26 <= io_in_r_bypass_5_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_3_df_is_ws_26 <= io_in_r_bypass_5_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_3_stall_26 <= io_in_r_bypass_5_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_0_data_26 <= io_in_r_bypass_6_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_0_load_store_26 <= io_in_r_bypass_6_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_0_df_is_ws_26 <= io_in_r_bypass_6_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_0_stall_26 <= io_in_r_bypass_6_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_1_data_26 <= io_in_r_bypass_6_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_1_load_store_26 <= io_in_r_bypass_6_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_1_df_is_ws_26 <= io_in_r_bypass_6_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_1_stall_26 <= io_in_r_bypass_6_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_2_data_26 <= io_in_r_bypass_6_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_2_load_store_26 <= io_in_r_bypass_6_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_2_df_is_ws_26 <= io_in_r_bypass_6_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_2_stall_26 <= io_in_r_bypass_6_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_3_data_26 <= io_in_r_bypass_6_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_3_load_store_26 <= io_in_r_bypass_6_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_3_df_is_ws_26 <= io_in_r_bypass_6_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_3_stall_26 <= io_in_r_bypass_6_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_0_data_26 <= io_in_r_bypass_7_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_0_load_store_26 <= io_in_r_bypass_7_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_0_df_is_ws_26 <= io_in_r_bypass_7_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_0_stall_26 <= io_in_r_bypass_7_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_1_data_26 <= io_in_r_bypass_7_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_1_load_store_26 <= io_in_r_bypass_7_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_1_df_is_ws_26 <= io_in_r_bypass_7_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_1_stall_26 <= io_in_r_bypass_7_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_2_data_26 <= io_in_r_bypass_7_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_2_load_store_26 <= io_in_r_bypass_7_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_2_df_is_ws_26 <= io_in_r_bypass_7_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_2_stall_26 <= io_in_r_bypass_7_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_3_data_26 <= io_in_r_bypass_7_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_3_load_store_26 <= io_in_r_bypass_7_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_3_df_is_ws_26 <= io_in_r_bypass_7_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_3_stall_26 <= io_in_r_bypass_7_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_0_data_26 <= io_in_r_bypass_8_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_0_load_store_26 <= io_in_r_bypass_8_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_0_df_is_ws_26 <= io_in_r_bypass_8_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_0_stall_26 <= io_in_r_bypass_8_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_1_data_26 <= io_in_r_bypass_8_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_1_load_store_26 <= io_in_r_bypass_8_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_1_df_is_ws_26 <= io_in_r_bypass_8_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_1_stall_26 <= io_in_r_bypass_8_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_2_data_26 <= io_in_r_bypass_8_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_2_load_store_26 <= io_in_r_bypass_8_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_2_df_is_ws_26 <= io_in_r_bypass_8_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_2_stall_26 <= io_in_r_bypass_8_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_3_data_26 <= io_in_r_bypass_8_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_3_load_store_26 <= io_in_r_bypass_8_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_3_df_is_ws_26 <= io_in_r_bypass_8_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_3_stall_26 <= io_in_r_bypass_8_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_0_data_26 <= io_in_r_bypass_9_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_0_load_store_26 <= io_in_r_bypass_9_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_0_df_is_ws_26 <= io_in_r_bypass_9_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_0_stall_26 <= io_in_r_bypass_9_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_1_data_26 <= io_in_r_bypass_9_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_1_load_store_26 <= io_in_r_bypass_9_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_1_df_is_ws_26 <= io_in_r_bypass_9_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_1_stall_26 <= io_in_r_bypass_9_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_2_data_26 <= io_in_r_bypass_9_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_2_load_store_26 <= io_in_r_bypass_9_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_2_df_is_ws_26 <= io_in_r_bypass_9_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_2_stall_26 <= io_in_r_bypass_9_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_3_data_26 <= io_in_r_bypass_9_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_3_load_store_26 <= io_in_r_bypass_9_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_3_df_is_ws_26 <= io_in_r_bypass_9_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_3_stall_26 <= io_in_r_bypass_9_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_0_data_26 <= io_in_r_bypass_10_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_0_load_store_26 <= io_in_r_bypass_10_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_0_df_is_ws_26 <= io_in_r_bypass_10_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_0_stall_26 <= io_in_r_bypass_10_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_1_data_26 <= io_in_r_bypass_10_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_1_load_store_26 <= io_in_r_bypass_10_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_1_df_is_ws_26 <= io_in_r_bypass_10_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_1_stall_26 <= io_in_r_bypass_10_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_2_data_26 <= io_in_r_bypass_10_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_2_load_store_26 <= io_in_r_bypass_10_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_2_df_is_ws_26 <= io_in_r_bypass_10_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_2_stall_26 <= io_in_r_bypass_10_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_3_data_26 <= io_in_r_bypass_10_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_3_load_store_26 <= io_in_r_bypass_10_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_3_df_is_ws_26 <= io_in_r_bypass_10_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_3_stall_26 <= io_in_r_bypass_10_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_0_data_26 <= io_in_r_bypass_11_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_0_load_store_26 <= io_in_r_bypass_11_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_0_df_is_ws_26 <= io_in_r_bypass_11_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_0_stall_26 <= io_in_r_bypass_11_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_1_data_26 <= io_in_r_bypass_11_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_1_load_store_26 <= io_in_r_bypass_11_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_1_df_is_ws_26 <= io_in_r_bypass_11_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_1_stall_26 <= io_in_r_bypass_11_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_2_data_26 <= io_in_r_bypass_11_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_2_load_store_26 <= io_in_r_bypass_11_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_2_df_is_ws_26 <= io_in_r_bypass_11_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_2_stall_26 <= io_in_r_bypass_11_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_3_data_26 <= io_in_r_bypass_11_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_3_load_store_26 <= io_in_r_bypass_11_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_3_df_is_ws_26 <= io_in_r_bypass_11_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_3_stall_26 <= io_in_r_bypass_11_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_0_data_26 <= io_in_r_bypass_12_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_0_load_store_26 <= io_in_r_bypass_12_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_0_df_is_ws_26 <= io_in_r_bypass_12_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_0_stall_26 <= io_in_r_bypass_12_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_1_data_26 <= io_in_r_bypass_12_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_1_load_store_26 <= io_in_r_bypass_12_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_1_df_is_ws_26 <= io_in_r_bypass_12_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_1_stall_26 <= io_in_r_bypass_12_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_2_data_26 <= io_in_r_bypass_12_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_2_load_store_26 <= io_in_r_bypass_12_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_2_df_is_ws_26 <= io_in_r_bypass_12_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_2_stall_26 <= io_in_r_bypass_12_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_3_data_26 <= io_in_r_bypass_12_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_3_load_store_26 <= io_in_r_bypass_12_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_3_df_is_ws_26 <= io_in_r_bypass_12_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_3_stall_26 <= io_in_r_bypass_12_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_0_data_26 <= io_in_r_bypass_13_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_0_load_store_26 <= io_in_r_bypass_13_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_0_df_is_ws_26 <= io_in_r_bypass_13_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_0_stall_26 <= io_in_r_bypass_13_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_1_data_26 <= io_in_r_bypass_13_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_1_load_store_26 <= io_in_r_bypass_13_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_1_df_is_ws_26 <= io_in_r_bypass_13_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_1_stall_26 <= io_in_r_bypass_13_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_2_data_26 <= io_in_r_bypass_13_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_2_load_store_26 <= io_in_r_bypass_13_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_2_df_is_ws_26 <= io_in_r_bypass_13_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_2_stall_26 <= io_in_r_bypass_13_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_3_data_26 <= io_in_r_bypass_13_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_3_load_store_26 <= io_in_r_bypass_13_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_3_df_is_ws_26 <= io_in_r_bypass_13_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_3_stall_26 <= io_in_r_bypass_13_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_0_data_26 <= io_in_r_bypass_14_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_0_load_store_26 <= io_in_r_bypass_14_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_0_df_is_ws_26 <= io_in_r_bypass_14_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_0_stall_26 <= io_in_r_bypass_14_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_1_data_26 <= io_in_r_bypass_14_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_1_load_store_26 <= io_in_r_bypass_14_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_1_df_is_ws_26 <= io_in_r_bypass_14_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_1_stall_26 <= io_in_r_bypass_14_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_2_data_26 <= io_in_r_bypass_14_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_2_load_store_26 <= io_in_r_bypass_14_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_2_df_is_ws_26 <= io_in_r_bypass_14_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_2_stall_26 <= io_in_r_bypass_14_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_3_data_26 <= io_in_r_bypass_14_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_3_load_store_26 <= io_in_r_bypass_14_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_3_df_is_ws_26 <= io_in_r_bypass_14_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_3_stall_26 <= io_in_r_bypass_14_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_0_data_26 <= io_in_r_bypass_15_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_0_load_store_26 <= io_in_r_bypass_15_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_0_df_is_ws_26 <= io_in_r_bypass_15_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_0_stall_26 <= io_in_r_bypass_15_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_1_data_26 <= io_in_r_bypass_15_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_1_load_store_26 <= io_in_r_bypass_15_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_1_df_is_ws_26 <= io_in_r_bypass_15_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_1_stall_26 <= io_in_r_bypass_15_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_2_data_26 <= io_in_r_bypass_15_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_2_load_store_26 <= io_in_r_bypass_15_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_2_df_is_ws_26 <= io_in_r_bypass_15_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_2_stall_26 <= io_in_r_bypass_15_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_3_data_26 <= io_in_r_bypass_15_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_3_load_store_26 <= io_in_r_bypass_15_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_3_df_is_ws_26 <= io_in_r_bypass_15_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_3_stall_26 <= io_in_r_bypass_15_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_0_data_26 <= io_in_r_bypass_16_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_0_load_store_26 <= io_in_r_bypass_16_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_0_df_is_ws_26 <= io_in_r_bypass_16_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_0_stall_26 <= io_in_r_bypass_16_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_1_data_26 <= io_in_r_bypass_16_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_1_load_store_26 <= io_in_r_bypass_16_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_1_df_is_ws_26 <= io_in_r_bypass_16_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_1_stall_26 <= io_in_r_bypass_16_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_2_data_26 <= io_in_r_bypass_16_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_2_load_store_26 <= io_in_r_bypass_16_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_2_df_is_ws_26 <= io_in_r_bypass_16_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_2_stall_26 <= io_in_r_bypass_16_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_3_data_26 <= io_in_r_bypass_16_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_3_load_store_26 <= io_in_r_bypass_16_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_3_df_is_ws_26 <= io_in_r_bypass_16_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_3_stall_26 <= io_in_r_bypass_16_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_0_data_26 <= io_in_r_bypass_17_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_0_load_store_26 <= io_in_r_bypass_17_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_0_df_is_ws_26 <= io_in_r_bypass_17_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_0_stall_26 <= io_in_r_bypass_17_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_1_data_26 <= io_in_r_bypass_17_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_1_load_store_26 <= io_in_r_bypass_17_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_1_df_is_ws_26 <= io_in_r_bypass_17_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_1_stall_26 <= io_in_r_bypass_17_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_2_data_26 <= io_in_r_bypass_17_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_2_load_store_26 <= io_in_r_bypass_17_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_2_df_is_ws_26 <= io_in_r_bypass_17_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_2_stall_26 <= io_in_r_bypass_17_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_3_data_26 <= io_in_r_bypass_17_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_3_load_store_26 <= io_in_r_bypass_17_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_3_df_is_ws_26 <= io_in_r_bypass_17_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_3_stall_26 <= io_in_r_bypass_17_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_0_data_26 <= io_in_r_bypass_18_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_0_load_store_26 <= io_in_r_bypass_18_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_0_df_is_ws_26 <= io_in_r_bypass_18_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_0_stall_26 <= io_in_r_bypass_18_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_1_data_26 <= io_in_r_bypass_18_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_1_load_store_26 <= io_in_r_bypass_18_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_1_df_is_ws_26 <= io_in_r_bypass_18_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_1_stall_26 <= io_in_r_bypass_18_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_2_data_26 <= io_in_r_bypass_18_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_2_load_store_26 <= io_in_r_bypass_18_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_2_df_is_ws_26 <= io_in_r_bypass_18_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_2_stall_26 <= io_in_r_bypass_18_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_3_data_26 <= io_in_r_bypass_18_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_3_load_store_26 <= io_in_r_bypass_18_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_3_df_is_ws_26 <= io_in_r_bypass_18_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_3_stall_26 <= io_in_r_bypass_18_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_0_data_26 <= io_in_r_bypass_19_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_0_load_store_26 <= io_in_r_bypass_19_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_0_df_is_ws_26 <= io_in_r_bypass_19_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_0_stall_26 <= io_in_r_bypass_19_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_1_data_26 <= io_in_r_bypass_19_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_1_load_store_26 <= io_in_r_bypass_19_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_1_df_is_ws_26 <= io_in_r_bypass_19_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_1_stall_26 <= io_in_r_bypass_19_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_2_data_26 <= io_in_r_bypass_19_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_2_load_store_26 <= io_in_r_bypass_19_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_2_df_is_ws_26 <= io_in_r_bypass_19_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_2_stall_26 <= io_in_r_bypass_19_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_3_data_26 <= io_in_r_bypass_19_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_3_load_store_26 <= io_in_r_bypass_19_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_3_df_is_ws_26 <= io_in_r_bypass_19_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_3_stall_26 <= io_in_r_bypass_19_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_0_data_26 <= io_in_r_bypass_20_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_0_load_store_26 <= io_in_r_bypass_20_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_0_df_is_ws_26 <= io_in_r_bypass_20_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_0_stall_26 <= io_in_r_bypass_20_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_1_data_26 <= io_in_r_bypass_20_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_1_load_store_26 <= io_in_r_bypass_20_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_1_df_is_ws_26 <= io_in_r_bypass_20_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_1_stall_26 <= io_in_r_bypass_20_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_2_data_26 <= io_in_r_bypass_20_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_2_load_store_26 <= io_in_r_bypass_20_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_2_df_is_ws_26 <= io_in_r_bypass_20_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_2_stall_26 <= io_in_r_bypass_20_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_3_data_26 <= io_in_r_bypass_20_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_3_load_store_26 <= io_in_r_bypass_20_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_3_df_is_ws_26 <= io_in_r_bypass_20_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_3_stall_26 <= io_in_r_bypass_20_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_0_data_26 <= io_in_r_bypass_21_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_0_load_store_26 <= io_in_r_bypass_21_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_0_df_is_ws_26 <= io_in_r_bypass_21_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_0_stall_26 <= io_in_r_bypass_21_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_1_data_26 <= io_in_r_bypass_21_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_1_load_store_26 <= io_in_r_bypass_21_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_1_df_is_ws_26 <= io_in_r_bypass_21_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_1_stall_26 <= io_in_r_bypass_21_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_2_data_26 <= io_in_r_bypass_21_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_2_load_store_26 <= io_in_r_bypass_21_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_2_df_is_ws_26 <= io_in_r_bypass_21_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_2_stall_26 <= io_in_r_bypass_21_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_3_data_26 <= io_in_r_bypass_21_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_3_load_store_26 <= io_in_r_bypass_21_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_3_df_is_ws_26 <= io_in_r_bypass_21_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_3_stall_26 <= io_in_r_bypass_21_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_0_data_26 <= io_in_r_bypass_22_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_0_load_store_26 <= io_in_r_bypass_22_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_0_df_is_ws_26 <= io_in_r_bypass_22_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_0_stall_26 <= io_in_r_bypass_22_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_1_data_26 <= io_in_r_bypass_22_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_1_load_store_26 <= io_in_r_bypass_22_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_1_df_is_ws_26 <= io_in_r_bypass_22_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_1_stall_26 <= io_in_r_bypass_22_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_2_data_26 <= io_in_r_bypass_22_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_2_load_store_26 <= io_in_r_bypass_22_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_2_df_is_ws_26 <= io_in_r_bypass_22_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_2_stall_26 <= io_in_r_bypass_22_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_3_data_26 <= io_in_r_bypass_22_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_3_load_store_26 <= io_in_r_bypass_22_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_3_df_is_ws_26 <= io_in_r_bypass_22_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_3_stall_26 <= io_in_r_bypass_22_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_0_data_26 <= io_in_r_bypass_23_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_0_load_store_26 <= io_in_r_bypass_23_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_0_df_is_ws_26 <= io_in_r_bypass_23_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_0_stall_26 <= io_in_r_bypass_23_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_1_data_26 <= io_in_r_bypass_23_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_1_load_store_26 <= io_in_r_bypass_23_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_1_df_is_ws_26 <= io_in_r_bypass_23_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_1_stall_26 <= io_in_r_bypass_23_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_2_data_26 <= io_in_r_bypass_23_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_2_load_store_26 <= io_in_r_bypass_23_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_2_df_is_ws_26 <= io_in_r_bypass_23_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_2_stall_26 <= io_in_r_bypass_23_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_3_data_26 <= io_in_r_bypass_23_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_3_load_store_26 <= io_in_r_bypass_23_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_3_df_is_ws_26 <= io_in_r_bypass_23_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_3_stall_26 <= io_in_r_bypass_23_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_0_data_26 <= io_in_r_bypass_24_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_0_load_store_26 <= io_in_r_bypass_24_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_0_df_is_ws_26 <= io_in_r_bypass_24_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_0_stall_26 <= io_in_r_bypass_24_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_1_data_26 <= io_in_r_bypass_24_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_1_load_store_26 <= io_in_r_bypass_24_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_1_df_is_ws_26 <= io_in_r_bypass_24_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_1_stall_26 <= io_in_r_bypass_24_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_2_data_26 <= io_in_r_bypass_24_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_2_load_store_26 <= io_in_r_bypass_24_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_2_df_is_ws_26 <= io_in_r_bypass_24_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_2_stall_26 <= io_in_r_bypass_24_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_3_data_26 <= io_in_r_bypass_24_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_3_load_store_26 <= io_in_r_bypass_24_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_3_df_is_ws_26 <= io_in_r_bypass_24_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_3_stall_26 <= io_in_r_bypass_24_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_0_data_26 <= io_in_r_bypass_25_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_0_load_store_26 <= io_in_r_bypass_25_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_0_df_is_ws_26 <= io_in_r_bypass_25_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_0_stall_26 <= io_in_r_bypass_25_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_1_data_26 <= io_in_r_bypass_25_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_1_load_store_26 <= io_in_r_bypass_25_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_1_df_is_ws_26 <= io_in_r_bypass_25_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_1_stall_26 <= io_in_r_bypass_25_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_2_data_26 <= io_in_r_bypass_25_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_2_load_store_26 <= io_in_r_bypass_25_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_2_df_is_ws_26 <= io_in_r_bypass_25_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_2_stall_26 <= io_in_r_bypass_25_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_3_data_26 <= io_in_r_bypass_25_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_3_load_store_26 <= io_in_r_bypass_25_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_3_df_is_ws_26 <= io_in_r_bypass_25_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_3_stall_26 <= io_in_r_bypass_25_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_0_data_26 <= io_in_r_bypass_26_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_0_load_store_26 <= io_in_r_bypass_26_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_0_df_is_ws_26 <= io_in_r_bypass_26_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_0_stall_26 <= io_in_r_bypass_26_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_1_data_26 <= io_in_r_bypass_26_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_1_load_store_26 <= io_in_r_bypass_26_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_1_df_is_ws_26 <= io_in_r_bypass_26_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_1_stall_26 <= io_in_r_bypass_26_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_2_data_26 <= io_in_r_bypass_26_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_2_load_store_26 <= io_in_r_bypass_26_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_2_df_is_ws_26 <= io_in_r_bypass_26_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_2_stall_26 <= io_in_r_bypass_26_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_3_data_26 <= io_in_r_bypass_26_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_3_load_store_26 <= io_in_r_bypass_26_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_3_df_is_ws_26 <= io_in_r_bypass_26_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_3_stall_26 <= io_in_r_bypass_26_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_0_data_26 <= io_in_r_bypass_27_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_0_load_store_26 <= io_in_r_bypass_27_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_0_df_is_ws_26 <= io_in_r_bypass_27_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_0_stall_26 <= io_in_r_bypass_27_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_1_data_26 <= io_in_r_bypass_27_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_1_load_store_26 <= io_in_r_bypass_27_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_1_df_is_ws_26 <= io_in_r_bypass_27_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_1_stall_26 <= io_in_r_bypass_27_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_2_data_26 <= io_in_r_bypass_27_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_2_load_store_26 <= io_in_r_bypass_27_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_2_df_is_ws_26 <= io_in_r_bypass_27_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_2_stall_26 <= io_in_r_bypass_27_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_3_data_26 <= io_in_r_bypass_27_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_3_load_store_26 <= io_in_r_bypass_27_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_3_df_is_ws_26 <= io_in_r_bypass_27_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_3_stall_26 <= io_in_r_bypass_27_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_0_data_26 <= io_in_r_bypass_28_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_0_load_store_26 <= io_in_r_bypass_28_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_0_df_is_ws_26 <= io_in_r_bypass_28_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_0_stall_26 <= io_in_r_bypass_28_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_1_data_26 <= io_in_r_bypass_28_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_1_load_store_26 <= io_in_r_bypass_28_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_1_df_is_ws_26 <= io_in_r_bypass_28_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_1_stall_26 <= io_in_r_bypass_28_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_2_data_26 <= io_in_r_bypass_28_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_2_load_store_26 <= io_in_r_bypass_28_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_2_df_is_ws_26 <= io_in_r_bypass_28_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_2_stall_26 <= io_in_r_bypass_28_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_3_data_26 <= io_in_r_bypass_28_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_3_load_store_26 <= io_in_r_bypass_28_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_3_df_is_ws_26 <= io_in_r_bypass_28_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_3_stall_26 <= io_in_r_bypass_28_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_0_data_26 <= io_in_r_bypass_29_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_0_load_store_26 <= io_in_r_bypass_29_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_0_df_is_ws_26 <= io_in_r_bypass_29_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_0_stall_26 <= io_in_r_bypass_29_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_1_data_26 <= io_in_r_bypass_29_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_1_load_store_26 <= io_in_r_bypass_29_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_1_df_is_ws_26 <= io_in_r_bypass_29_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_1_stall_26 <= io_in_r_bypass_29_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_2_data_26 <= io_in_r_bypass_29_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_2_load_store_26 <= io_in_r_bypass_29_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_2_df_is_ws_26 <= io_in_r_bypass_29_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_2_stall_26 <= io_in_r_bypass_29_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_3_data_26 <= io_in_r_bypass_29_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_3_load_store_26 <= io_in_r_bypass_29_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_3_df_is_ws_26 <= io_in_r_bypass_29_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_3_stall_26 <= io_in_r_bypass_29_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_0_data_26 <= io_in_r_bypass_30_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_0_load_store_26 <= io_in_r_bypass_30_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_0_df_is_ws_26 <= io_in_r_bypass_30_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_0_stall_26 <= io_in_r_bypass_30_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_1_data_26 <= io_in_r_bypass_30_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_1_load_store_26 <= io_in_r_bypass_30_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_1_df_is_ws_26 <= io_in_r_bypass_30_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_1_stall_26 <= io_in_r_bypass_30_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_2_data_26 <= io_in_r_bypass_30_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_2_load_store_26 <= io_in_r_bypass_30_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_2_df_is_ws_26 <= io_in_r_bypass_30_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_2_stall_26 <= io_in_r_bypass_30_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_3_data_26 <= io_in_r_bypass_30_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_3_load_store_26 <= io_in_r_bypass_30_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_3_df_is_ws_26 <= io_in_r_bypass_30_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_3_stall_26 <= io_in_r_bypass_30_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_0_data_26 <= io_in_r_bypass_31_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_0_load_store_26 <= io_in_r_bypass_31_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_0_df_is_ws_26 <= io_in_r_bypass_31_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_0_stall_26 <= io_in_r_bypass_31_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_1_data_26 <= io_in_r_bypass_31_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_1_load_store_26 <= io_in_r_bypass_31_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_1_df_is_ws_26 <= io_in_r_bypass_31_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_1_stall_26 <= io_in_r_bypass_31_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_2_data_26 <= io_in_r_bypass_31_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_2_load_store_26 <= io_in_r_bypass_31_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_2_df_is_ws_26 <= io_in_r_bypass_31_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_2_stall_26 <= io_in_r_bypass_31_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_3_data_26 <= io_in_r_bypass_31_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_3_load_store_26 <= io_in_r_bypass_31_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_3_df_is_ws_26 <= io_in_r_bypass_31_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_3_stall_26 <= io_in_r_bypass_31_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_0_data_27 <= io_in_r_bypass_0_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_0_load_store_27 <= io_in_r_bypass_0_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_0_df_is_ws_27 <= io_in_r_bypass_0_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_0_stall_27 <= io_in_r_bypass_0_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_1_data_27 <= io_in_r_bypass_0_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_1_load_store_27 <= io_in_r_bypass_0_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_1_df_is_ws_27 <= io_in_r_bypass_0_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_1_stall_27 <= io_in_r_bypass_0_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_2_data_27 <= io_in_r_bypass_0_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_2_load_store_27 <= io_in_r_bypass_0_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_2_df_is_ws_27 <= io_in_r_bypass_0_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_2_stall_27 <= io_in_r_bypass_0_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_3_data_27 <= io_in_r_bypass_0_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_3_load_store_27 <= io_in_r_bypass_0_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_3_df_is_ws_27 <= io_in_r_bypass_0_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_3_stall_27 <= io_in_r_bypass_0_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_0_data_27 <= io_in_r_bypass_1_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_0_load_store_27 <= io_in_r_bypass_1_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_0_df_is_ws_27 <= io_in_r_bypass_1_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_0_stall_27 <= io_in_r_bypass_1_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_1_data_27 <= io_in_r_bypass_1_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_1_load_store_27 <= io_in_r_bypass_1_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_1_df_is_ws_27 <= io_in_r_bypass_1_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_1_stall_27 <= io_in_r_bypass_1_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_2_data_27 <= io_in_r_bypass_1_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_2_load_store_27 <= io_in_r_bypass_1_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_2_df_is_ws_27 <= io_in_r_bypass_1_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_2_stall_27 <= io_in_r_bypass_1_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_3_data_27 <= io_in_r_bypass_1_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_3_load_store_27 <= io_in_r_bypass_1_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_3_df_is_ws_27 <= io_in_r_bypass_1_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_3_stall_27 <= io_in_r_bypass_1_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_0_data_27 <= io_in_r_bypass_2_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_0_load_store_27 <= io_in_r_bypass_2_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_0_df_is_ws_27 <= io_in_r_bypass_2_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_0_stall_27 <= io_in_r_bypass_2_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_1_data_27 <= io_in_r_bypass_2_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_1_load_store_27 <= io_in_r_bypass_2_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_1_df_is_ws_27 <= io_in_r_bypass_2_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_1_stall_27 <= io_in_r_bypass_2_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_2_data_27 <= io_in_r_bypass_2_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_2_load_store_27 <= io_in_r_bypass_2_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_2_df_is_ws_27 <= io_in_r_bypass_2_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_2_stall_27 <= io_in_r_bypass_2_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_3_data_27 <= io_in_r_bypass_2_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_3_load_store_27 <= io_in_r_bypass_2_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_3_df_is_ws_27 <= io_in_r_bypass_2_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_3_stall_27 <= io_in_r_bypass_2_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_0_data_27 <= io_in_r_bypass_3_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_0_load_store_27 <= io_in_r_bypass_3_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_0_df_is_ws_27 <= io_in_r_bypass_3_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_0_stall_27 <= io_in_r_bypass_3_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_1_data_27 <= io_in_r_bypass_3_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_1_load_store_27 <= io_in_r_bypass_3_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_1_df_is_ws_27 <= io_in_r_bypass_3_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_1_stall_27 <= io_in_r_bypass_3_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_2_data_27 <= io_in_r_bypass_3_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_2_load_store_27 <= io_in_r_bypass_3_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_2_df_is_ws_27 <= io_in_r_bypass_3_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_2_stall_27 <= io_in_r_bypass_3_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_3_data_27 <= io_in_r_bypass_3_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_3_load_store_27 <= io_in_r_bypass_3_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_3_df_is_ws_27 <= io_in_r_bypass_3_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_3_stall_27 <= io_in_r_bypass_3_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_0_data_27 <= io_in_r_bypass_4_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_0_load_store_27 <= io_in_r_bypass_4_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_0_df_is_ws_27 <= io_in_r_bypass_4_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_0_stall_27 <= io_in_r_bypass_4_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_1_data_27 <= io_in_r_bypass_4_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_1_load_store_27 <= io_in_r_bypass_4_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_1_df_is_ws_27 <= io_in_r_bypass_4_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_1_stall_27 <= io_in_r_bypass_4_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_2_data_27 <= io_in_r_bypass_4_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_2_load_store_27 <= io_in_r_bypass_4_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_2_df_is_ws_27 <= io_in_r_bypass_4_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_2_stall_27 <= io_in_r_bypass_4_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_3_data_27 <= io_in_r_bypass_4_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_3_load_store_27 <= io_in_r_bypass_4_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_3_df_is_ws_27 <= io_in_r_bypass_4_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_3_stall_27 <= io_in_r_bypass_4_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_0_data_27 <= io_in_r_bypass_5_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_0_load_store_27 <= io_in_r_bypass_5_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_0_df_is_ws_27 <= io_in_r_bypass_5_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_0_stall_27 <= io_in_r_bypass_5_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_1_data_27 <= io_in_r_bypass_5_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_1_load_store_27 <= io_in_r_bypass_5_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_1_df_is_ws_27 <= io_in_r_bypass_5_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_1_stall_27 <= io_in_r_bypass_5_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_2_data_27 <= io_in_r_bypass_5_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_2_load_store_27 <= io_in_r_bypass_5_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_2_df_is_ws_27 <= io_in_r_bypass_5_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_2_stall_27 <= io_in_r_bypass_5_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_3_data_27 <= io_in_r_bypass_5_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_3_load_store_27 <= io_in_r_bypass_5_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_3_df_is_ws_27 <= io_in_r_bypass_5_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_3_stall_27 <= io_in_r_bypass_5_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_0_data_27 <= io_in_r_bypass_6_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_0_load_store_27 <= io_in_r_bypass_6_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_0_df_is_ws_27 <= io_in_r_bypass_6_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_0_stall_27 <= io_in_r_bypass_6_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_1_data_27 <= io_in_r_bypass_6_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_1_load_store_27 <= io_in_r_bypass_6_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_1_df_is_ws_27 <= io_in_r_bypass_6_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_1_stall_27 <= io_in_r_bypass_6_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_2_data_27 <= io_in_r_bypass_6_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_2_load_store_27 <= io_in_r_bypass_6_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_2_df_is_ws_27 <= io_in_r_bypass_6_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_2_stall_27 <= io_in_r_bypass_6_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_3_data_27 <= io_in_r_bypass_6_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_3_load_store_27 <= io_in_r_bypass_6_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_3_df_is_ws_27 <= io_in_r_bypass_6_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_3_stall_27 <= io_in_r_bypass_6_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_0_data_27 <= io_in_r_bypass_7_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_0_load_store_27 <= io_in_r_bypass_7_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_0_df_is_ws_27 <= io_in_r_bypass_7_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_0_stall_27 <= io_in_r_bypass_7_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_1_data_27 <= io_in_r_bypass_7_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_1_load_store_27 <= io_in_r_bypass_7_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_1_df_is_ws_27 <= io_in_r_bypass_7_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_1_stall_27 <= io_in_r_bypass_7_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_2_data_27 <= io_in_r_bypass_7_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_2_load_store_27 <= io_in_r_bypass_7_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_2_df_is_ws_27 <= io_in_r_bypass_7_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_2_stall_27 <= io_in_r_bypass_7_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_3_data_27 <= io_in_r_bypass_7_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_3_load_store_27 <= io_in_r_bypass_7_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_3_df_is_ws_27 <= io_in_r_bypass_7_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_3_stall_27 <= io_in_r_bypass_7_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_0_data_27 <= io_in_r_bypass_8_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_0_load_store_27 <= io_in_r_bypass_8_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_0_df_is_ws_27 <= io_in_r_bypass_8_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_0_stall_27 <= io_in_r_bypass_8_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_1_data_27 <= io_in_r_bypass_8_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_1_load_store_27 <= io_in_r_bypass_8_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_1_df_is_ws_27 <= io_in_r_bypass_8_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_1_stall_27 <= io_in_r_bypass_8_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_2_data_27 <= io_in_r_bypass_8_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_2_load_store_27 <= io_in_r_bypass_8_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_2_df_is_ws_27 <= io_in_r_bypass_8_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_2_stall_27 <= io_in_r_bypass_8_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_3_data_27 <= io_in_r_bypass_8_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_3_load_store_27 <= io_in_r_bypass_8_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_3_df_is_ws_27 <= io_in_r_bypass_8_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_3_stall_27 <= io_in_r_bypass_8_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_0_data_27 <= io_in_r_bypass_9_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_0_load_store_27 <= io_in_r_bypass_9_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_0_df_is_ws_27 <= io_in_r_bypass_9_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_0_stall_27 <= io_in_r_bypass_9_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_1_data_27 <= io_in_r_bypass_9_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_1_load_store_27 <= io_in_r_bypass_9_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_1_df_is_ws_27 <= io_in_r_bypass_9_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_1_stall_27 <= io_in_r_bypass_9_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_2_data_27 <= io_in_r_bypass_9_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_2_load_store_27 <= io_in_r_bypass_9_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_2_df_is_ws_27 <= io_in_r_bypass_9_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_2_stall_27 <= io_in_r_bypass_9_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_3_data_27 <= io_in_r_bypass_9_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_3_load_store_27 <= io_in_r_bypass_9_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_3_df_is_ws_27 <= io_in_r_bypass_9_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_3_stall_27 <= io_in_r_bypass_9_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_0_data_27 <= io_in_r_bypass_10_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_0_load_store_27 <= io_in_r_bypass_10_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_0_df_is_ws_27 <= io_in_r_bypass_10_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_0_stall_27 <= io_in_r_bypass_10_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_1_data_27 <= io_in_r_bypass_10_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_1_load_store_27 <= io_in_r_bypass_10_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_1_df_is_ws_27 <= io_in_r_bypass_10_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_1_stall_27 <= io_in_r_bypass_10_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_2_data_27 <= io_in_r_bypass_10_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_2_load_store_27 <= io_in_r_bypass_10_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_2_df_is_ws_27 <= io_in_r_bypass_10_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_2_stall_27 <= io_in_r_bypass_10_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_3_data_27 <= io_in_r_bypass_10_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_3_load_store_27 <= io_in_r_bypass_10_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_3_df_is_ws_27 <= io_in_r_bypass_10_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_3_stall_27 <= io_in_r_bypass_10_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_0_data_27 <= io_in_r_bypass_11_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_0_load_store_27 <= io_in_r_bypass_11_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_0_df_is_ws_27 <= io_in_r_bypass_11_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_0_stall_27 <= io_in_r_bypass_11_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_1_data_27 <= io_in_r_bypass_11_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_1_load_store_27 <= io_in_r_bypass_11_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_1_df_is_ws_27 <= io_in_r_bypass_11_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_1_stall_27 <= io_in_r_bypass_11_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_2_data_27 <= io_in_r_bypass_11_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_2_load_store_27 <= io_in_r_bypass_11_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_2_df_is_ws_27 <= io_in_r_bypass_11_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_2_stall_27 <= io_in_r_bypass_11_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_3_data_27 <= io_in_r_bypass_11_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_3_load_store_27 <= io_in_r_bypass_11_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_3_df_is_ws_27 <= io_in_r_bypass_11_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_3_stall_27 <= io_in_r_bypass_11_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_0_data_27 <= io_in_r_bypass_12_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_0_load_store_27 <= io_in_r_bypass_12_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_0_df_is_ws_27 <= io_in_r_bypass_12_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_0_stall_27 <= io_in_r_bypass_12_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_1_data_27 <= io_in_r_bypass_12_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_1_load_store_27 <= io_in_r_bypass_12_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_1_df_is_ws_27 <= io_in_r_bypass_12_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_1_stall_27 <= io_in_r_bypass_12_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_2_data_27 <= io_in_r_bypass_12_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_2_load_store_27 <= io_in_r_bypass_12_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_2_df_is_ws_27 <= io_in_r_bypass_12_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_2_stall_27 <= io_in_r_bypass_12_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_3_data_27 <= io_in_r_bypass_12_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_3_load_store_27 <= io_in_r_bypass_12_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_3_df_is_ws_27 <= io_in_r_bypass_12_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_3_stall_27 <= io_in_r_bypass_12_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_0_data_27 <= io_in_r_bypass_13_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_0_load_store_27 <= io_in_r_bypass_13_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_0_df_is_ws_27 <= io_in_r_bypass_13_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_0_stall_27 <= io_in_r_bypass_13_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_1_data_27 <= io_in_r_bypass_13_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_1_load_store_27 <= io_in_r_bypass_13_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_1_df_is_ws_27 <= io_in_r_bypass_13_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_1_stall_27 <= io_in_r_bypass_13_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_2_data_27 <= io_in_r_bypass_13_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_2_load_store_27 <= io_in_r_bypass_13_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_2_df_is_ws_27 <= io_in_r_bypass_13_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_2_stall_27 <= io_in_r_bypass_13_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_3_data_27 <= io_in_r_bypass_13_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_3_load_store_27 <= io_in_r_bypass_13_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_3_df_is_ws_27 <= io_in_r_bypass_13_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_3_stall_27 <= io_in_r_bypass_13_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_0_data_27 <= io_in_r_bypass_14_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_0_load_store_27 <= io_in_r_bypass_14_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_0_df_is_ws_27 <= io_in_r_bypass_14_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_0_stall_27 <= io_in_r_bypass_14_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_1_data_27 <= io_in_r_bypass_14_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_1_load_store_27 <= io_in_r_bypass_14_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_1_df_is_ws_27 <= io_in_r_bypass_14_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_1_stall_27 <= io_in_r_bypass_14_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_2_data_27 <= io_in_r_bypass_14_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_2_load_store_27 <= io_in_r_bypass_14_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_2_df_is_ws_27 <= io_in_r_bypass_14_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_2_stall_27 <= io_in_r_bypass_14_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_3_data_27 <= io_in_r_bypass_14_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_3_load_store_27 <= io_in_r_bypass_14_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_3_df_is_ws_27 <= io_in_r_bypass_14_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_3_stall_27 <= io_in_r_bypass_14_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_0_data_27 <= io_in_r_bypass_15_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_0_load_store_27 <= io_in_r_bypass_15_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_0_df_is_ws_27 <= io_in_r_bypass_15_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_0_stall_27 <= io_in_r_bypass_15_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_1_data_27 <= io_in_r_bypass_15_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_1_load_store_27 <= io_in_r_bypass_15_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_1_df_is_ws_27 <= io_in_r_bypass_15_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_1_stall_27 <= io_in_r_bypass_15_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_2_data_27 <= io_in_r_bypass_15_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_2_load_store_27 <= io_in_r_bypass_15_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_2_df_is_ws_27 <= io_in_r_bypass_15_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_2_stall_27 <= io_in_r_bypass_15_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_3_data_27 <= io_in_r_bypass_15_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_3_load_store_27 <= io_in_r_bypass_15_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_3_df_is_ws_27 <= io_in_r_bypass_15_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_3_stall_27 <= io_in_r_bypass_15_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_0_data_27 <= io_in_r_bypass_16_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_0_load_store_27 <= io_in_r_bypass_16_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_0_df_is_ws_27 <= io_in_r_bypass_16_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_0_stall_27 <= io_in_r_bypass_16_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_1_data_27 <= io_in_r_bypass_16_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_1_load_store_27 <= io_in_r_bypass_16_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_1_df_is_ws_27 <= io_in_r_bypass_16_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_1_stall_27 <= io_in_r_bypass_16_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_2_data_27 <= io_in_r_bypass_16_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_2_load_store_27 <= io_in_r_bypass_16_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_2_df_is_ws_27 <= io_in_r_bypass_16_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_2_stall_27 <= io_in_r_bypass_16_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_3_data_27 <= io_in_r_bypass_16_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_3_load_store_27 <= io_in_r_bypass_16_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_3_df_is_ws_27 <= io_in_r_bypass_16_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_3_stall_27 <= io_in_r_bypass_16_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_0_data_27 <= io_in_r_bypass_17_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_0_load_store_27 <= io_in_r_bypass_17_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_0_df_is_ws_27 <= io_in_r_bypass_17_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_0_stall_27 <= io_in_r_bypass_17_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_1_data_27 <= io_in_r_bypass_17_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_1_load_store_27 <= io_in_r_bypass_17_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_1_df_is_ws_27 <= io_in_r_bypass_17_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_1_stall_27 <= io_in_r_bypass_17_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_2_data_27 <= io_in_r_bypass_17_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_2_load_store_27 <= io_in_r_bypass_17_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_2_df_is_ws_27 <= io_in_r_bypass_17_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_2_stall_27 <= io_in_r_bypass_17_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_3_data_27 <= io_in_r_bypass_17_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_3_load_store_27 <= io_in_r_bypass_17_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_3_df_is_ws_27 <= io_in_r_bypass_17_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_3_stall_27 <= io_in_r_bypass_17_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_0_data_27 <= io_in_r_bypass_18_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_0_load_store_27 <= io_in_r_bypass_18_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_0_df_is_ws_27 <= io_in_r_bypass_18_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_0_stall_27 <= io_in_r_bypass_18_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_1_data_27 <= io_in_r_bypass_18_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_1_load_store_27 <= io_in_r_bypass_18_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_1_df_is_ws_27 <= io_in_r_bypass_18_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_1_stall_27 <= io_in_r_bypass_18_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_2_data_27 <= io_in_r_bypass_18_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_2_load_store_27 <= io_in_r_bypass_18_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_2_df_is_ws_27 <= io_in_r_bypass_18_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_2_stall_27 <= io_in_r_bypass_18_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_3_data_27 <= io_in_r_bypass_18_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_3_load_store_27 <= io_in_r_bypass_18_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_3_df_is_ws_27 <= io_in_r_bypass_18_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_3_stall_27 <= io_in_r_bypass_18_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_0_data_27 <= io_in_r_bypass_19_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_0_load_store_27 <= io_in_r_bypass_19_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_0_df_is_ws_27 <= io_in_r_bypass_19_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_0_stall_27 <= io_in_r_bypass_19_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_1_data_27 <= io_in_r_bypass_19_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_1_load_store_27 <= io_in_r_bypass_19_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_1_df_is_ws_27 <= io_in_r_bypass_19_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_1_stall_27 <= io_in_r_bypass_19_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_2_data_27 <= io_in_r_bypass_19_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_2_load_store_27 <= io_in_r_bypass_19_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_2_df_is_ws_27 <= io_in_r_bypass_19_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_2_stall_27 <= io_in_r_bypass_19_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_3_data_27 <= io_in_r_bypass_19_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_3_load_store_27 <= io_in_r_bypass_19_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_3_df_is_ws_27 <= io_in_r_bypass_19_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_3_stall_27 <= io_in_r_bypass_19_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_0_data_27 <= io_in_r_bypass_20_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_0_load_store_27 <= io_in_r_bypass_20_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_0_df_is_ws_27 <= io_in_r_bypass_20_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_0_stall_27 <= io_in_r_bypass_20_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_1_data_27 <= io_in_r_bypass_20_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_1_load_store_27 <= io_in_r_bypass_20_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_1_df_is_ws_27 <= io_in_r_bypass_20_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_1_stall_27 <= io_in_r_bypass_20_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_2_data_27 <= io_in_r_bypass_20_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_2_load_store_27 <= io_in_r_bypass_20_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_2_df_is_ws_27 <= io_in_r_bypass_20_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_2_stall_27 <= io_in_r_bypass_20_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_3_data_27 <= io_in_r_bypass_20_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_3_load_store_27 <= io_in_r_bypass_20_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_3_df_is_ws_27 <= io_in_r_bypass_20_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_3_stall_27 <= io_in_r_bypass_20_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_0_data_27 <= io_in_r_bypass_21_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_0_load_store_27 <= io_in_r_bypass_21_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_0_df_is_ws_27 <= io_in_r_bypass_21_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_0_stall_27 <= io_in_r_bypass_21_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_1_data_27 <= io_in_r_bypass_21_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_1_load_store_27 <= io_in_r_bypass_21_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_1_df_is_ws_27 <= io_in_r_bypass_21_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_1_stall_27 <= io_in_r_bypass_21_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_2_data_27 <= io_in_r_bypass_21_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_2_load_store_27 <= io_in_r_bypass_21_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_2_df_is_ws_27 <= io_in_r_bypass_21_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_2_stall_27 <= io_in_r_bypass_21_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_3_data_27 <= io_in_r_bypass_21_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_3_load_store_27 <= io_in_r_bypass_21_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_3_df_is_ws_27 <= io_in_r_bypass_21_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_3_stall_27 <= io_in_r_bypass_21_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_0_data_27 <= io_in_r_bypass_22_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_0_load_store_27 <= io_in_r_bypass_22_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_0_df_is_ws_27 <= io_in_r_bypass_22_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_0_stall_27 <= io_in_r_bypass_22_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_1_data_27 <= io_in_r_bypass_22_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_1_load_store_27 <= io_in_r_bypass_22_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_1_df_is_ws_27 <= io_in_r_bypass_22_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_1_stall_27 <= io_in_r_bypass_22_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_2_data_27 <= io_in_r_bypass_22_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_2_load_store_27 <= io_in_r_bypass_22_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_2_df_is_ws_27 <= io_in_r_bypass_22_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_2_stall_27 <= io_in_r_bypass_22_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_3_data_27 <= io_in_r_bypass_22_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_3_load_store_27 <= io_in_r_bypass_22_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_3_df_is_ws_27 <= io_in_r_bypass_22_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_3_stall_27 <= io_in_r_bypass_22_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_0_data_27 <= io_in_r_bypass_23_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_0_load_store_27 <= io_in_r_bypass_23_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_0_df_is_ws_27 <= io_in_r_bypass_23_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_0_stall_27 <= io_in_r_bypass_23_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_1_data_27 <= io_in_r_bypass_23_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_1_load_store_27 <= io_in_r_bypass_23_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_1_df_is_ws_27 <= io_in_r_bypass_23_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_1_stall_27 <= io_in_r_bypass_23_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_2_data_27 <= io_in_r_bypass_23_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_2_load_store_27 <= io_in_r_bypass_23_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_2_df_is_ws_27 <= io_in_r_bypass_23_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_2_stall_27 <= io_in_r_bypass_23_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_3_data_27 <= io_in_r_bypass_23_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_3_load_store_27 <= io_in_r_bypass_23_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_3_df_is_ws_27 <= io_in_r_bypass_23_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_3_stall_27 <= io_in_r_bypass_23_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_0_data_27 <= io_in_r_bypass_24_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_0_load_store_27 <= io_in_r_bypass_24_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_0_df_is_ws_27 <= io_in_r_bypass_24_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_0_stall_27 <= io_in_r_bypass_24_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_1_data_27 <= io_in_r_bypass_24_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_1_load_store_27 <= io_in_r_bypass_24_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_1_df_is_ws_27 <= io_in_r_bypass_24_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_1_stall_27 <= io_in_r_bypass_24_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_2_data_27 <= io_in_r_bypass_24_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_2_load_store_27 <= io_in_r_bypass_24_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_2_df_is_ws_27 <= io_in_r_bypass_24_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_2_stall_27 <= io_in_r_bypass_24_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_3_data_27 <= io_in_r_bypass_24_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_3_load_store_27 <= io_in_r_bypass_24_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_3_df_is_ws_27 <= io_in_r_bypass_24_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_3_stall_27 <= io_in_r_bypass_24_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_0_data_27 <= io_in_r_bypass_25_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_0_load_store_27 <= io_in_r_bypass_25_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_0_df_is_ws_27 <= io_in_r_bypass_25_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_0_stall_27 <= io_in_r_bypass_25_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_1_data_27 <= io_in_r_bypass_25_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_1_load_store_27 <= io_in_r_bypass_25_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_1_df_is_ws_27 <= io_in_r_bypass_25_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_1_stall_27 <= io_in_r_bypass_25_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_2_data_27 <= io_in_r_bypass_25_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_2_load_store_27 <= io_in_r_bypass_25_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_2_df_is_ws_27 <= io_in_r_bypass_25_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_2_stall_27 <= io_in_r_bypass_25_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_3_data_27 <= io_in_r_bypass_25_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_3_load_store_27 <= io_in_r_bypass_25_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_3_df_is_ws_27 <= io_in_r_bypass_25_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_3_stall_27 <= io_in_r_bypass_25_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_0_data_27 <= io_in_r_bypass_26_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_0_load_store_27 <= io_in_r_bypass_26_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_0_df_is_ws_27 <= io_in_r_bypass_26_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_0_stall_27 <= io_in_r_bypass_26_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_1_data_27 <= io_in_r_bypass_26_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_1_load_store_27 <= io_in_r_bypass_26_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_1_df_is_ws_27 <= io_in_r_bypass_26_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_1_stall_27 <= io_in_r_bypass_26_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_2_data_27 <= io_in_r_bypass_26_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_2_load_store_27 <= io_in_r_bypass_26_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_2_df_is_ws_27 <= io_in_r_bypass_26_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_2_stall_27 <= io_in_r_bypass_26_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_3_data_27 <= io_in_r_bypass_26_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_3_load_store_27 <= io_in_r_bypass_26_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_3_df_is_ws_27 <= io_in_r_bypass_26_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_3_stall_27 <= io_in_r_bypass_26_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_0_data_27 <= io_in_r_bypass_27_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_0_load_store_27 <= io_in_r_bypass_27_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_0_df_is_ws_27 <= io_in_r_bypass_27_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_0_stall_27 <= io_in_r_bypass_27_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_1_data_27 <= io_in_r_bypass_27_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_1_load_store_27 <= io_in_r_bypass_27_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_1_df_is_ws_27 <= io_in_r_bypass_27_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_1_stall_27 <= io_in_r_bypass_27_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_2_data_27 <= io_in_r_bypass_27_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_2_load_store_27 <= io_in_r_bypass_27_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_2_df_is_ws_27 <= io_in_r_bypass_27_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_2_stall_27 <= io_in_r_bypass_27_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_3_data_27 <= io_in_r_bypass_27_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_3_load_store_27 <= io_in_r_bypass_27_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_3_df_is_ws_27 <= io_in_r_bypass_27_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_3_stall_27 <= io_in_r_bypass_27_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_0_data_27 <= io_in_r_bypass_28_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_0_load_store_27 <= io_in_r_bypass_28_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_0_df_is_ws_27 <= io_in_r_bypass_28_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_0_stall_27 <= io_in_r_bypass_28_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_1_data_27 <= io_in_r_bypass_28_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_1_load_store_27 <= io_in_r_bypass_28_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_1_df_is_ws_27 <= io_in_r_bypass_28_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_1_stall_27 <= io_in_r_bypass_28_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_2_data_27 <= io_in_r_bypass_28_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_2_load_store_27 <= io_in_r_bypass_28_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_2_df_is_ws_27 <= io_in_r_bypass_28_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_2_stall_27 <= io_in_r_bypass_28_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_3_data_27 <= io_in_r_bypass_28_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_3_load_store_27 <= io_in_r_bypass_28_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_3_df_is_ws_27 <= io_in_r_bypass_28_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_3_stall_27 <= io_in_r_bypass_28_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_0_data_27 <= io_in_r_bypass_29_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_0_load_store_27 <= io_in_r_bypass_29_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_0_df_is_ws_27 <= io_in_r_bypass_29_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_0_stall_27 <= io_in_r_bypass_29_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_1_data_27 <= io_in_r_bypass_29_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_1_load_store_27 <= io_in_r_bypass_29_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_1_df_is_ws_27 <= io_in_r_bypass_29_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_1_stall_27 <= io_in_r_bypass_29_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_2_data_27 <= io_in_r_bypass_29_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_2_load_store_27 <= io_in_r_bypass_29_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_2_df_is_ws_27 <= io_in_r_bypass_29_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_2_stall_27 <= io_in_r_bypass_29_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_3_data_27 <= io_in_r_bypass_29_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_3_load_store_27 <= io_in_r_bypass_29_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_3_df_is_ws_27 <= io_in_r_bypass_29_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_3_stall_27 <= io_in_r_bypass_29_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_0_data_27 <= io_in_r_bypass_30_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_0_load_store_27 <= io_in_r_bypass_30_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_0_df_is_ws_27 <= io_in_r_bypass_30_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_0_stall_27 <= io_in_r_bypass_30_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_1_data_27 <= io_in_r_bypass_30_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_1_load_store_27 <= io_in_r_bypass_30_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_1_df_is_ws_27 <= io_in_r_bypass_30_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_1_stall_27 <= io_in_r_bypass_30_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_2_data_27 <= io_in_r_bypass_30_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_2_load_store_27 <= io_in_r_bypass_30_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_2_df_is_ws_27 <= io_in_r_bypass_30_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_2_stall_27 <= io_in_r_bypass_30_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_3_data_27 <= io_in_r_bypass_30_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_3_load_store_27 <= io_in_r_bypass_30_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_3_df_is_ws_27 <= io_in_r_bypass_30_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_3_stall_27 <= io_in_r_bypass_30_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_0_data_27 <= io_in_r_bypass_31_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_0_load_store_27 <= io_in_r_bypass_31_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_0_df_is_ws_27 <= io_in_r_bypass_31_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_0_stall_27 <= io_in_r_bypass_31_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_1_data_27 <= io_in_r_bypass_31_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_1_load_store_27 <= io_in_r_bypass_31_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_1_df_is_ws_27 <= io_in_r_bypass_31_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_1_stall_27 <= io_in_r_bypass_31_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_2_data_27 <= io_in_r_bypass_31_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_2_load_store_27 <= io_in_r_bypass_31_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_2_df_is_ws_27 <= io_in_r_bypass_31_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_2_stall_27 <= io_in_r_bypass_31_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_3_data_27 <= io_in_r_bypass_31_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_3_load_store_27 <= io_in_r_bypass_31_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_3_df_is_ws_27 <= io_in_r_bypass_31_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_3_stall_27 <= io_in_r_bypass_31_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_0_data_28 <= io_in_r_bypass_0_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_0_load_store_28 <= io_in_r_bypass_0_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_0_df_is_ws_28 <= io_in_r_bypass_0_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_0_stall_28 <= io_in_r_bypass_0_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_1_data_28 <= io_in_r_bypass_0_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_1_load_store_28 <= io_in_r_bypass_0_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_1_df_is_ws_28 <= io_in_r_bypass_0_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_1_stall_28 <= io_in_r_bypass_0_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_2_data_28 <= io_in_r_bypass_0_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_2_load_store_28 <= io_in_r_bypass_0_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_2_df_is_ws_28 <= io_in_r_bypass_0_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_2_stall_28 <= io_in_r_bypass_0_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_3_data_28 <= io_in_r_bypass_0_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_3_load_store_28 <= io_in_r_bypass_0_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_3_df_is_ws_28 <= io_in_r_bypass_0_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_3_stall_28 <= io_in_r_bypass_0_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_0_data_28 <= io_in_r_bypass_1_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_0_load_store_28 <= io_in_r_bypass_1_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_0_df_is_ws_28 <= io_in_r_bypass_1_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_0_stall_28 <= io_in_r_bypass_1_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_1_data_28 <= io_in_r_bypass_1_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_1_load_store_28 <= io_in_r_bypass_1_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_1_df_is_ws_28 <= io_in_r_bypass_1_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_1_stall_28 <= io_in_r_bypass_1_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_2_data_28 <= io_in_r_bypass_1_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_2_load_store_28 <= io_in_r_bypass_1_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_2_df_is_ws_28 <= io_in_r_bypass_1_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_2_stall_28 <= io_in_r_bypass_1_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_3_data_28 <= io_in_r_bypass_1_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_3_load_store_28 <= io_in_r_bypass_1_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_3_df_is_ws_28 <= io_in_r_bypass_1_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_3_stall_28 <= io_in_r_bypass_1_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_0_data_28 <= io_in_r_bypass_2_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_0_load_store_28 <= io_in_r_bypass_2_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_0_df_is_ws_28 <= io_in_r_bypass_2_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_0_stall_28 <= io_in_r_bypass_2_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_1_data_28 <= io_in_r_bypass_2_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_1_load_store_28 <= io_in_r_bypass_2_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_1_df_is_ws_28 <= io_in_r_bypass_2_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_1_stall_28 <= io_in_r_bypass_2_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_2_data_28 <= io_in_r_bypass_2_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_2_load_store_28 <= io_in_r_bypass_2_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_2_df_is_ws_28 <= io_in_r_bypass_2_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_2_stall_28 <= io_in_r_bypass_2_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_3_data_28 <= io_in_r_bypass_2_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_3_load_store_28 <= io_in_r_bypass_2_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_3_df_is_ws_28 <= io_in_r_bypass_2_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_3_stall_28 <= io_in_r_bypass_2_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_0_data_28 <= io_in_r_bypass_3_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_0_load_store_28 <= io_in_r_bypass_3_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_0_df_is_ws_28 <= io_in_r_bypass_3_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_0_stall_28 <= io_in_r_bypass_3_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_1_data_28 <= io_in_r_bypass_3_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_1_load_store_28 <= io_in_r_bypass_3_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_1_df_is_ws_28 <= io_in_r_bypass_3_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_1_stall_28 <= io_in_r_bypass_3_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_2_data_28 <= io_in_r_bypass_3_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_2_load_store_28 <= io_in_r_bypass_3_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_2_df_is_ws_28 <= io_in_r_bypass_3_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_2_stall_28 <= io_in_r_bypass_3_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_3_data_28 <= io_in_r_bypass_3_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_3_load_store_28 <= io_in_r_bypass_3_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_3_df_is_ws_28 <= io_in_r_bypass_3_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_3_stall_28 <= io_in_r_bypass_3_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_0_data_28 <= io_in_r_bypass_4_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_0_load_store_28 <= io_in_r_bypass_4_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_0_df_is_ws_28 <= io_in_r_bypass_4_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_0_stall_28 <= io_in_r_bypass_4_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_1_data_28 <= io_in_r_bypass_4_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_1_load_store_28 <= io_in_r_bypass_4_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_1_df_is_ws_28 <= io_in_r_bypass_4_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_1_stall_28 <= io_in_r_bypass_4_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_2_data_28 <= io_in_r_bypass_4_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_2_load_store_28 <= io_in_r_bypass_4_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_2_df_is_ws_28 <= io_in_r_bypass_4_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_2_stall_28 <= io_in_r_bypass_4_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_3_data_28 <= io_in_r_bypass_4_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_3_load_store_28 <= io_in_r_bypass_4_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_3_df_is_ws_28 <= io_in_r_bypass_4_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_3_stall_28 <= io_in_r_bypass_4_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_0_data_28 <= io_in_r_bypass_5_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_0_load_store_28 <= io_in_r_bypass_5_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_0_df_is_ws_28 <= io_in_r_bypass_5_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_0_stall_28 <= io_in_r_bypass_5_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_1_data_28 <= io_in_r_bypass_5_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_1_load_store_28 <= io_in_r_bypass_5_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_1_df_is_ws_28 <= io_in_r_bypass_5_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_1_stall_28 <= io_in_r_bypass_5_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_2_data_28 <= io_in_r_bypass_5_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_2_load_store_28 <= io_in_r_bypass_5_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_2_df_is_ws_28 <= io_in_r_bypass_5_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_2_stall_28 <= io_in_r_bypass_5_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_3_data_28 <= io_in_r_bypass_5_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_3_load_store_28 <= io_in_r_bypass_5_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_3_df_is_ws_28 <= io_in_r_bypass_5_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_3_stall_28 <= io_in_r_bypass_5_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_0_data_28 <= io_in_r_bypass_6_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_0_load_store_28 <= io_in_r_bypass_6_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_0_df_is_ws_28 <= io_in_r_bypass_6_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_0_stall_28 <= io_in_r_bypass_6_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_1_data_28 <= io_in_r_bypass_6_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_1_load_store_28 <= io_in_r_bypass_6_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_1_df_is_ws_28 <= io_in_r_bypass_6_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_1_stall_28 <= io_in_r_bypass_6_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_2_data_28 <= io_in_r_bypass_6_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_2_load_store_28 <= io_in_r_bypass_6_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_2_df_is_ws_28 <= io_in_r_bypass_6_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_2_stall_28 <= io_in_r_bypass_6_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_3_data_28 <= io_in_r_bypass_6_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_3_load_store_28 <= io_in_r_bypass_6_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_3_df_is_ws_28 <= io_in_r_bypass_6_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_3_stall_28 <= io_in_r_bypass_6_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_0_data_28 <= io_in_r_bypass_7_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_0_load_store_28 <= io_in_r_bypass_7_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_0_df_is_ws_28 <= io_in_r_bypass_7_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_0_stall_28 <= io_in_r_bypass_7_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_1_data_28 <= io_in_r_bypass_7_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_1_load_store_28 <= io_in_r_bypass_7_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_1_df_is_ws_28 <= io_in_r_bypass_7_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_1_stall_28 <= io_in_r_bypass_7_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_2_data_28 <= io_in_r_bypass_7_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_2_load_store_28 <= io_in_r_bypass_7_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_2_df_is_ws_28 <= io_in_r_bypass_7_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_2_stall_28 <= io_in_r_bypass_7_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_3_data_28 <= io_in_r_bypass_7_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_3_load_store_28 <= io_in_r_bypass_7_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_3_df_is_ws_28 <= io_in_r_bypass_7_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_3_stall_28 <= io_in_r_bypass_7_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_0_data_28 <= io_in_r_bypass_8_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_0_load_store_28 <= io_in_r_bypass_8_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_0_df_is_ws_28 <= io_in_r_bypass_8_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_0_stall_28 <= io_in_r_bypass_8_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_1_data_28 <= io_in_r_bypass_8_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_1_load_store_28 <= io_in_r_bypass_8_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_1_df_is_ws_28 <= io_in_r_bypass_8_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_1_stall_28 <= io_in_r_bypass_8_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_2_data_28 <= io_in_r_bypass_8_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_2_load_store_28 <= io_in_r_bypass_8_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_2_df_is_ws_28 <= io_in_r_bypass_8_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_2_stall_28 <= io_in_r_bypass_8_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_3_data_28 <= io_in_r_bypass_8_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_3_load_store_28 <= io_in_r_bypass_8_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_3_df_is_ws_28 <= io_in_r_bypass_8_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_3_stall_28 <= io_in_r_bypass_8_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_0_data_28 <= io_in_r_bypass_9_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_0_load_store_28 <= io_in_r_bypass_9_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_0_df_is_ws_28 <= io_in_r_bypass_9_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_0_stall_28 <= io_in_r_bypass_9_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_1_data_28 <= io_in_r_bypass_9_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_1_load_store_28 <= io_in_r_bypass_9_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_1_df_is_ws_28 <= io_in_r_bypass_9_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_1_stall_28 <= io_in_r_bypass_9_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_2_data_28 <= io_in_r_bypass_9_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_2_load_store_28 <= io_in_r_bypass_9_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_2_df_is_ws_28 <= io_in_r_bypass_9_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_2_stall_28 <= io_in_r_bypass_9_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_3_data_28 <= io_in_r_bypass_9_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_3_load_store_28 <= io_in_r_bypass_9_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_3_df_is_ws_28 <= io_in_r_bypass_9_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_3_stall_28 <= io_in_r_bypass_9_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_0_data_28 <= io_in_r_bypass_10_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_0_load_store_28 <= io_in_r_bypass_10_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_0_df_is_ws_28 <= io_in_r_bypass_10_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_0_stall_28 <= io_in_r_bypass_10_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_1_data_28 <= io_in_r_bypass_10_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_1_load_store_28 <= io_in_r_bypass_10_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_1_df_is_ws_28 <= io_in_r_bypass_10_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_1_stall_28 <= io_in_r_bypass_10_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_2_data_28 <= io_in_r_bypass_10_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_2_load_store_28 <= io_in_r_bypass_10_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_2_df_is_ws_28 <= io_in_r_bypass_10_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_2_stall_28 <= io_in_r_bypass_10_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_3_data_28 <= io_in_r_bypass_10_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_3_load_store_28 <= io_in_r_bypass_10_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_3_df_is_ws_28 <= io_in_r_bypass_10_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_3_stall_28 <= io_in_r_bypass_10_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_0_data_28 <= io_in_r_bypass_11_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_0_load_store_28 <= io_in_r_bypass_11_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_0_df_is_ws_28 <= io_in_r_bypass_11_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_0_stall_28 <= io_in_r_bypass_11_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_1_data_28 <= io_in_r_bypass_11_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_1_load_store_28 <= io_in_r_bypass_11_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_1_df_is_ws_28 <= io_in_r_bypass_11_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_1_stall_28 <= io_in_r_bypass_11_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_2_data_28 <= io_in_r_bypass_11_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_2_load_store_28 <= io_in_r_bypass_11_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_2_df_is_ws_28 <= io_in_r_bypass_11_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_2_stall_28 <= io_in_r_bypass_11_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_3_data_28 <= io_in_r_bypass_11_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_3_load_store_28 <= io_in_r_bypass_11_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_3_df_is_ws_28 <= io_in_r_bypass_11_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_3_stall_28 <= io_in_r_bypass_11_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_0_data_28 <= io_in_r_bypass_12_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_0_load_store_28 <= io_in_r_bypass_12_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_0_df_is_ws_28 <= io_in_r_bypass_12_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_0_stall_28 <= io_in_r_bypass_12_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_1_data_28 <= io_in_r_bypass_12_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_1_load_store_28 <= io_in_r_bypass_12_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_1_df_is_ws_28 <= io_in_r_bypass_12_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_1_stall_28 <= io_in_r_bypass_12_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_2_data_28 <= io_in_r_bypass_12_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_2_load_store_28 <= io_in_r_bypass_12_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_2_df_is_ws_28 <= io_in_r_bypass_12_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_2_stall_28 <= io_in_r_bypass_12_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_3_data_28 <= io_in_r_bypass_12_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_3_load_store_28 <= io_in_r_bypass_12_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_3_df_is_ws_28 <= io_in_r_bypass_12_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_3_stall_28 <= io_in_r_bypass_12_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_0_data_28 <= io_in_r_bypass_13_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_0_load_store_28 <= io_in_r_bypass_13_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_0_df_is_ws_28 <= io_in_r_bypass_13_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_0_stall_28 <= io_in_r_bypass_13_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_1_data_28 <= io_in_r_bypass_13_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_1_load_store_28 <= io_in_r_bypass_13_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_1_df_is_ws_28 <= io_in_r_bypass_13_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_1_stall_28 <= io_in_r_bypass_13_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_2_data_28 <= io_in_r_bypass_13_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_2_load_store_28 <= io_in_r_bypass_13_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_2_df_is_ws_28 <= io_in_r_bypass_13_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_2_stall_28 <= io_in_r_bypass_13_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_3_data_28 <= io_in_r_bypass_13_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_3_load_store_28 <= io_in_r_bypass_13_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_3_df_is_ws_28 <= io_in_r_bypass_13_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_3_stall_28 <= io_in_r_bypass_13_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_0_data_28 <= io_in_r_bypass_14_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_0_load_store_28 <= io_in_r_bypass_14_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_0_df_is_ws_28 <= io_in_r_bypass_14_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_0_stall_28 <= io_in_r_bypass_14_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_1_data_28 <= io_in_r_bypass_14_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_1_load_store_28 <= io_in_r_bypass_14_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_1_df_is_ws_28 <= io_in_r_bypass_14_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_1_stall_28 <= io_in_r_bypass_14_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_2_data_28 <= io_in_r_bypass_14_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_2_load_store_28 <= io_in_r_bypass_14_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_2_df_is_ws_28 <= io_in_r_bypass_14_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_2_stall_28 <= io_in_r_bypass_14_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_3_data_28 <= io_in_r_bypass_14_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_3_load_store_28 <= io_in_r_bypass_14_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_3_df_is_ws_28 <= io_in_r_bypass_14_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_3_stall_28 <= io_in_r_bypass_14_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_0_data_28 <= io_in_r_bypass_15_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_0_load_store_28 <= io_in_r_bypass_15_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_0_df_is_ws_28 <= io_in_r_bypass_15_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_0_stall_28 <= io_in_r_bypass_15_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_1_data_28 <= io_in_r_bypass_15_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_1_load_store_28 <= io_in_r_bypass_15_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_1_df_is_ws_28 <= io_in_r_bypass_15_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_1_stall_28 <= io_in_r_bypass_15_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_2_data_28 <= io_in_r_bypass_15_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_2_load_store_28 <= io_in_r_bypass_15_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_2_df_is_ws_28 <= io_in_r_bypass_15_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_2_stall_28 <= io_in_r_bypass_15_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_3_data_28 <= io_in_r_bypass_15_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_3_load_store_28 <= io_in_r_bypass_15_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_3_df_is_ws_28 <= io_in_r_bypass_15_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_3_stall_28 <= io_in_r_bypass_15_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_0_data_28 <= io_in_r_bypass_16_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_0_load_store_28 <= io_in_r_bypass_16_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_0_df_is_ws_28 <= io_in_r_bypass_16_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_0_stall_28 <= io_in_r_bypass_16_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_1_data_28 <= io_in_r_bypass_16_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_1_load_store_28 <= io_in_r_bypass_16_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_1_df_is_ws_28 <= io_in_r_bypass_16_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_1_stall_28 <= io_in_r_bypass_16_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_2_data_28 <= io_in_r_bypass_16_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_2_load_store_28 <= io_in_r_bypass_16_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_2_df_is_ws_28 <= io_in_r_bypass_16_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_2_stall_28 <= io_in_r_bypass_16_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_3_data_28 <= io_in_r_bypass_16_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_3_load_store_28 <= io_in_r_bypass_16_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_3_df_is_ws_28 <= io_in_r_bypass_16_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_3_stall_28 <= io_in_r_bypass_16_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_0_data_28 <= io_in_r_bypass_17_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_0_load_store_28 <= io_in_r_bypass_17_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_0_df_is_ws_28 <= io_in_r_bypass_17_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_0_stall_28 <= io_in_r_bypass_17_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_1_data_28 <= io_in_r_bypass_17_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_1_load_store_28 <= io_in_r_bypass_17_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_1_df_is_ws_28 <= io_in_r_bypass_17_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_1_stall_28 <= io_in_r_bypass_17_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_2_data_28 <= io_in_r_bypass_17_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_2_load_store_28 <= io_in_r_bypass_17_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_2_df_is_ws_28 <= io_in_r_bypass_17_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_2_stall_28 <= io_in_r_bypass_17_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_3_data_28 <= io_in_r_bypass_17_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_3_load_store_28 <= io_in_r_bypass_17_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_3_df_is_ws_28 <= io_in_r_bypass_17_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_3_stall_28 <= io_in_r_bypass_17_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_0_data_28 <= io_in_r_bypass_18_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_0_load_store_28 <= io_in_r_bypass_18_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_0_df_is_ws_28 <= io_in_r_bypass_18_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_0_stall_28 <= io_in_r_bypass_18_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_1_data_28 <= io_in_r_bypass_18_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_1_load_store_28 <= io_in_r_bypass_18_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_1_df_is_ws_28 <= io_in_r_bypass_18_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_1_stall_28 <= io_in_r_bypass_18_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_2_data_28 <= io_in_r_bypass_18_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_2_load_store_28 <= io_in_r_bypass_18_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_2_df_is_ws_28 <= io_in_r_bypass_18_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_2_stall_28 <= io_in_r_bypass_18_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_3_data_28 <= io_in_r_bypass_18_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_3_load_store_28 <= io_in_r_bypass_18_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_3_df_is_ws_28 <= io_in_r_bypass_18_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_3_stall_28 <= io_in_r_bypass_18_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_0_data_28 <= io_in_r_bypass_19_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_0_load_store_28 <= io_in_r_bypass_19_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_0_df_is_ws_28 <= io_in_r_bypass_19_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_0_stall_28 <= io_in_r_bypass_19_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_1_data_28 <= io_in_r_bypass_19_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_1_load_store_28 <= io_in_r_bypass_19_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_1_df_is_ws_28 <= io_in_r_bypass_19_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_1_stall_28 <= io_in_r_bypass_19_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_2_data_28 <= io_in_r_bypass_19_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_2_load_store_28 <= io_in_r_bypass_19_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_2_df_is_ws_28 <= io_in_r_bypass_19_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_2_stall_28 <= io_in_r_bypass_19_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_3_data_28 <= io_in_r_bypass_19_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_3_load_store_28 <= io_in_r_bypass_19_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_3_df_is_ws_28 <= io_in_r_bypass_19_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_3_stall_28 <= io_in_r_bypass_19_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_0_data_28 <= io_in_r_bypass_20_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_0_load_store_28 <= io_in_r_bypass_20_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_0_df_is_ws_28 <= io_in_r_bypass_20_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_0_stall_28 <= io_in_r_bypass_20_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_1_data_28 <= io_in_r_bypass_20_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_1_load_store_28 <= io_in_r_bypass_20_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_1_df_is_ws_28 <= io_in_r_bypass_20_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_1_stall_28 <= io_in_r_bypass_20_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_2_data_28 <= io_in_r_bypass_20_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_2_load_store_28 <= io_in_r_bypass_20_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_2_df_is_ws_28 <= io_in_r_bypass_20_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_2_stall_28 <= io_in_r_bypass_20_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_3_data_28 <= io_in_r_bypass_20_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_3_load_store_28 <= io_in_r_bypass_20_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_3_df_is_ws_28 <= io_in_r_bypass_20_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_3_stall_28 <= io_in_r_bypass_20_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_0_data_28 <= io_in_r_bypass_21_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_0_load_store_28 <= io_in_r_bypass_21_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_0_df_is_ws_28 <= io_in_r_bypass_21_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_0_stall_28 <= io_in_r_bypass_21_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_1_data_28 <= io_in_r_bypass_21_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_1_load_store_28 <= io_in_r_bypass_21_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_1_df_is_ws_28 <= io_in_r_bypass_21_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_1_stall_28 <= io_in_r_bypass_21_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_2_data_28 <= io_in_r_bypass_21_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_2_load_store_28 <= io_in_r_bypass_21_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_2_df_is_ws_28 <= io_in_r_bypass_21_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_2_stall_28 <= io_in_r_bypass_21_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_3_data_28 <= io_in_r_bypass_21_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_3_load_store_28 <= io_in_r_bypass_21_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_3_df_is_ws_28 <= io_in_r_bypass_21_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_3_stall_28 <= io_in_r_bypass_21_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_0_data_28 <= io_in_r_bypass_22_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_0_load_store_28 <= io_in_r_bypass_22_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_0_df_is_ws_28 <= io_in_r_bypass_22_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_0_stall_28 <= io_in_r_bypass_22_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_1_data_28 <= io_in_r_bypass_22_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_1_load_store_28 <= io_in_r_bypass_22_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_1_df_is_ws_28 <= io_in_r_bypass_22_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_1_stall_28 <= io_in_r_bypass_22_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_2_data_28 <= io_in_r_bypass_22_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_2_load_store_28 <= io_in_r_bypass_22_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_2_df_is_ws_28 <= io_in_r_bypass_22_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_2_stall_28 <= io_in_r_bypass_22_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_3_data_28 <= io_in_r_bypass_22_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_3_load_store_28 <= io_in_r_bypass_22_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_3_df_is_ws_28 <= io_in_r_bypass_22_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_3_stall_28 <= io_in_r_bypass_22_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_0_data_28 <= io_in_r_bypass_23_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_0_load_store_28 <= io_in_r_bypass_23_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_0_df_is_ws_28 <= io_in_r_bypass_23_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_0_stall_28 <= io_in_r_bypass_23_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_1_data_28 <= io_in_r_bypass_23_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_1_load_store_28 <= io_in_r_bypass_23_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_1_df_is_ws_28 <= io_in_r_bypass_23_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_1_stall_28 <= io_in_r_bypass_23_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_2_data_28 <= io_in_r_bypass_23_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_2_load_store_28 <= io_in_r_bypass_23_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_2_df_is_ws_28 <= io_in_r_bypass_23_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_2_stall_28 <= io_in_r_bypass_23_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_3_data_28 <= io_in_r_bypass_23_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_3_load_store_28 <= io_in_r_bypass_23_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_3_df_is_ws_28 <= io_in_r_bypass_23_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_3_stall_28 <= io_in_r_bypass_23_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_0_data_28 <= io_in_r_bypass_24_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_0_load_store_28 <= io_in_r_bypass_24_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_0_df_is_ws_28 <= io_in_r_bypass_24_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_0_stall_28 <= io_in_r_bypass_24_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_1_data_28 <= io_in_r_bypass_24_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_1_load_store_28 <= io_in_r_bypass_24_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_1_df_is_ws_28 <= io_in_r_bypass_24_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_1_stall_28 <= io_in_r_bypass_24_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_2_data_28 <= io_in_r_bypass_24_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_2_load_store_28 <= io_in_r_bypass_24_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_2_df_is_ws_28 <= io_in_r_bypass_24_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_2_stall_28 <= io_in_r_bypass_24_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_3_data_28 <= io_in_r_bypass_24_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_3_load_store_28 <= io_in_r_bypass_24_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_3_df_is_ws_28 <= io_in_r_bypass_24_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_3_stall_28 <= io_in_r_bypass_24_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_0_data_28 <= io_in_r_bypass_25_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_0_load_store_28 <= io_in_r_bypass_25_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_0_df_is_ws_28 <= io_in_r_bypass_25_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_0_stall_28 <= io_in_r_bypass_25_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_1_data_28 <= io_in_r_bypass_25_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_1_load_store_28 <= io_in_r_bypass_25_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_1_df_is_ws_28 <= io_in_r_bypass_25_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_1_stall_28 <= io_in_r_bypass_25_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_2_data_28 <= io_in_r_bypass_25_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_2_load_store_28 <= io_in_r_bypass_25_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_2_df_is_ws_28 <= io_in_r_bypass_25_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_2_stall_28 <= io_in_r_bypass_25_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_3_data_28 <= io_in_r_bypass_25_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_3_load_store_28 <= io_in_r_bypass_25_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_3_df_is_ws_28 <= io_in_r_bypass_25_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_3_stall_28 <= io_in_r_bypass_25_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_0_data_28 <= io_in_r_bypass_26_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_0_load_store_28 <= io_in_r_bypass_26_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_0_df_is_ws_28 <= io_in_r_bypass_26_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_0_stall_28 <= io_in_r_bypass_26_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_1_data_28 <= io_in_r_bypass_26_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_1_load_store_28 <= io_in_r_bypass_26_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_1_df_is_ws_28 <= io_in_r_bypass_26_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_1_stall_28 <= io_in_r_bypass_26_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_2_data_28 <= io_in_r_bypass_26_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_2_load_store_28 <= io_in_r_bypass_26_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_2_df_is_ws_28 <= io_in_r_bypass_26_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_2_stall_28 <= io_in_r_bypass_26_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_3_data_28 <= io_in_r_bypass_26_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_3_load_store_28 <= io_in_r_bypass_26_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_3_df_is_ws_28 <= io_in_r_bypass_26_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_3_stall_28 <= io_in_r_bypass_26_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_0_data_28 <= io_in_r_bypass_27_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_0_load_store_28 <= io_in_r_bypass_27_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_0_df_is_ws_28 <= io_in_r_bypass_27_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_0_stall_28 <= io_in_r_bypass_27_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_1_data_28 <= io_in_r_bypass_27_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_1_load_store_28 <= io_in_r_bypass_27_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_1_df_is_ws_28 <= io_in_r_bypass_27_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_1_stall_28 <= io_in_r_bypass_27_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_2_data_28 <= io_in_r_bypass_27_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_2_load_store_28 <= io_in_r_bypass_27_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_2_df_is_ws_28 <= io_in_r_bypass_27_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_2_stall_28 <= io_in_r_bypass_27_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_3_data_28 <= io_in_r_bypass_27_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_3_load_store_28 <= io_in_r_bypass_27_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_3_df_is_ws_28 <= io_in_r_bypass_27_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_3_stall_28 <= io_in_r_bypass_27_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_0_data_28 <= io_in_r_bypass_28_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_0_load_store_28 <= io_in_r_bypass_28_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_0_df_is_ws_28 <= io_in_r_bypass_28_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_0_stall_28 <= io_in_r_bypass_28_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_1_data_28 <= io_in_r_bypass_28_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_1_load_store_28 <= io_in_r_bypass_28_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_1_df_is_ws_28 <= io_in_r_bypass_28_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_1_stall_28 <= io_in_r_bypass_28_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_2_data_28 <= io_in_r_bypass_28_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_2_load_store_28 <= io_in_r_bypass_28_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_2_df_is_ws_28 <= io_in_r_bypass_28_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_2_stall_28 <= io_in_r_bypass_28_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_3_data_28 <= io_in_r_bypass_28_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_3_load_store_28 <= io_in_r_bypass_28_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_3_df_is_ws_28 <= io_in_r_bypass_28_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_3_stall_28 <= io_in_r_bypass_28_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_0_data_28 <= io_in_r_bypass_29_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_0_load_store_28 <= io_in_r_bypass_29_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_0_df_is_ws_28 <= io_in_r_bypass_29_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_0_stall_28 <= io_in_r_bypass_29_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_1_data_28 <= io_in_r_bypass_29_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_1_load_store_28 <= io_in_r_bypass_29_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_1_df_is_ws_28 <= io_in_r_bypass_29_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_1_stall_28 <= io_in_r_bypass_29_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_2_data_28 <= io_in_r_bypass_29_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_2_load_store_28 <= io_in_r_bypass_29_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_2_df_is_ws_28 <= io_in_r_bypass_29_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_2_stall_28 <= io_in_r_bypass_29_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_3_data_28 <= io_in_r_bypass_29_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_3_load_store_28 <= io_in_r_bypass_29_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_3_df_is_ws_28 <= io_in_r_bypass_29_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_3_stall_28 <= io_in_r_bypass_29_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_0_data_28 <= io_in_r_bypass_30_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_0_load_store_28 <= io_in_r_bypass_30_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_0_df_is_ws_28 <= io_in_r_bypass_30_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_0_stall_28 <= io_in_r_bypass_30_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_1_data_28 <= io_in_r_bypass_30_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_1_load_store_28 <= io_in_r_bypass_30_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_1_df_is_ws_28 <= io_in_r_bypass_30_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_1_stall_28 <= io_in_r_bypass_30_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_2_data_28 <= io_in_r_bypass_30_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_2_load_store_28 <= io_in_r_bypass_30_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_2_df_is_ws_28 <= io_in_r_bypass_30_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_2_stall_28 <= io_in_r_bypass_30_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_3_data_28 <= io_in_r_bypass_30_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_3_load_store_28 <= io_in_r_bypass_30_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_3_df_is_ws_28 <= io_in_r_bypass_30_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_3_stall_28 <= io_in_r_bypass_30_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_0_data_28 <= io_in_r_bypass_31_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_0_load_store_28 <= io_in_r_bypass_31_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_0_df_is_ws_28 <= io_in_r_bypass_31_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_0_stall_28 <= io_in_r_bypass_31_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_1_data_28 <= io_in_r_bypass_31_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_1_load_store_28 <= io_in_r_bypass_31_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_1_df_is_ws_28 <= io_in_r_bypass_31_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_1_stall_28 <= io_in_r_bypass_31_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_2_data_28 <= io_in_r_bypass_31_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_2_load_store_28 <= io_in_r_bypass_31_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_2_df_is_ws_28 <= io_in_r_bypass_31_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_2_stall_28 <= io_in_r_bypass_31_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_3_data_28 <= io_in_r_bypass_31_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_3_load_store_28 <= io_in_r_bypass_31_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_3_df_is_ws_28 <= io_in_r_bypass_31_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_3_stall_28 <= io_in_r_bypass_31_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_0_data_29 <= io_in_r_bypass_0_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_0_load_store_29 <= io_in_r_bypass_0_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_0_df_is_ws_29 <= io_in_r_bypass_0_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_0_stall_29 <= io_in_r_bypass_0_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_1_data_29 <= io_in_r_bypass_0_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_1_load_store_29 <= io_in_r_bypass_0_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_1_df_is_ws_29 <= io_in_r_bypass_0_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_1_stall_29 <= io_in_r_bypass_0_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_2_data_29 <= io_in_r_bypass_0_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_2_load_store_29 <= io_in_r_bypass_0_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_2_df_is_ws_29 <= io_in_r_bypass_0_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_2_stall_29 <= io_in_r_bypass_0_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_3_data_29 <= io_in_r_bypass_0_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_3_load_store_29 <= io_in_r_bypass_0_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_3_df_is_ws_29 <= io_in_r_bypass_0_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_3_stall_29 <= io_in_r_bypass_0_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_0_data_29 <= io_in_r_bypass_1_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_0_load_store_29 <= io_in_r_bypass_1_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_0_df_is_ws_29 <= io_in_r_bypass_1_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_0_stall_29 <= io_in_r_bypass_1_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_1_data_29 <= io_in_r_bypass_1_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_1_load_store_29 <= io_in_r_bypass_1_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_1_df_is_ws_29 <= io_in_r_bypass_1_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_1_stall_29 <= io_in_r_bypass_1_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_2_data_29 <= io_in_r_bypass_1_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_2_load_store_29 <= io_in_r_bypass_1_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_2_df_is_ws_29 <= io_in_r_bypass_1_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_2_stall_29 <= io_in_r_bypass_1_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_3_data_29 <= io_in_r_bypass_1_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_3_load_store_29 <= io_in_r_bypass_1_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_3_df_is_ws_29 <= io_in_r_bypass_1_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_3_stall_29 <= io_in_r_bypass_1_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_0_data_29 <= io_in_r_bypass_2_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_0_load_store_29 <= io_in_r_bypass_2_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_0_df_is_ws_29 <= io_in_r_bypass_2_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_0_stall_29 <= io_in_r_bypass_2_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_1_data_29 <= io_in_r_bypass_2_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_1_load_store_29 <= io_in_r_bypass_2_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_1_df_is_ws_29 <= io_in_r_bypass_2_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_1_stall_29 <= io_in_r_bypass_2_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_2_data_29 <= io_in_r_bypass_2_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_2_load_store_29 <= io_in_r_bypass_2_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_2_df_is_ws_29 <= io_in_r_bypass_2_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_2_stall_29 <= io_in_r_bypass_2_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_3_data_29 <= io_in_r_bypass_2_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_3_load_store_29 <= io_in_r_bypass_2_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_3_df_is_ws_29 <= io_in_r_bypass_2_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_3_stall_29 <= io_in_r_bypass_2_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_0_data_29 <= io_in_r_bypass_3_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_0_load_store_29 <= io_in_r_bypass_3_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_0_df_is_ws_29 <= io_in_r_bypass_3_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_0_stall_29 <= io_in_r_bypass_3_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_1_data_29 <= io_in_r_bypass_3_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_1_load_store_29 <= io_in_r_bypass_3_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_1_df_is_ws_29 <= io_in_r_bypass_3_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_1_stall_29 <= io_in_r_bypass_3_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_2_data_29 <= io_in_r_bypass_3_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_2_load_store_29 <= io_in_r_bypass_3_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_2_df_is_ws_29 <= io_in_r_bypass_3_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_2_stall_29 <= io_in_r_bypass_3_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_3_data_29 <= io_in_r_bypass_3_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_3_load_store_29 <= io_in_r_bypass_3_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_3_df_is_ws_29 <= io_in_r_bypass_3_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_3_stall_29 <= io_in_r_bypass_3_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_0_data_29 <= io_in_r_bypass_4_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_0_load_store_29 <= io_in_r_bypass_4_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_0_df_is_ws_29 <= io_in_r_bypass_4_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_0_stall_29 <= io_in_r_bypass_4_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_1_data_29 <= io_in_r_bypass_4_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_1_load_store_29 <= io_in_r_bypass_4_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_1_df_is_ws_29 <= io_in_r_bypass_4_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_1_stall_29 <= io_in_r_bypass_4_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_2_data_29 <= io_in_r_bypass_4_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_2_load_store_29 <= io_in_r_bypass_4_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_2_df_is_ws_29 <= io_in_r_bypass_4_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_2_stall_29 <= io_in_r_bypass_4_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_3_data_29 <= io_in_r_bypass_4_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_3_load_store_29 <= io_in_r_bypass_4_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_3_df_is_ws_29 <= io_in_r_bypass_4_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_3_stall_29 <= io_in_r_bypass_4_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_0_data_29 <= io_in_r_bypass_5_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_0_load_store_29 <= io_in_r_bypass_5_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_0_df_is_ws_29 <= io_in_r_bypass_5_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_0_stall_29 <= io_in_r_bypass_5_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_1_data_29 <= io_in_r_bypass_5_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_1_load_store_29 <= io_in_r_bypass_5_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_1_df_is_ws_29 <= io_in_r_bypass_5_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_1_stall_29 <= io_in_r_bypass_5_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_2_data_29 <= io_in_r_bypass_5_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_2_load_store_29 <= io_in_r_bypass_5_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_2_df_is_ws_29 <= io_in_r_bypass_5_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_2_stall_29 <= io_in_r_bypass_5_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_3_data_29 <= io_in_r_bypass_5_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_3_load_store_29 <= io_in_r_bypass_5_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_3_df_is_ws_29 <= io_in_r_bypass_5_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_3_stall_29 <= io_in_r_bypass_5_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_0_data_29 <= io_in_r_bypass_6_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_0_load_store_29 <= io_in_r_bypass_6_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_0_df_is_ws_29 <= io_in_r_bypass_6_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_0_stall_29 <= io_in_r_bypass_6_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_1_data_29 <= io_in_r_bypass_6_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_1_load_store_29 <= io_in_r_bypass_6_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_1_df_is_ws_29 <= io_in_r_bypass_6_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_1_stall_29 <= io_in_r_bypass_6_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_2_data_29 <= io_in_r_bypass_6_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_2_load_store_29 <= io_in_r_bypass_6_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_2_df_is_ws_29 <= io_in_r_bypass_6_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_2_stall_29 <= io_in_r_bypass_6_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_3_data_29 <= io_in_r_bypass_6_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_3_load_store_29 <= io_in_r_bypass_6_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_3_df_is_ws_29 <= io_in_r_bypass_6_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_3_stall_29 <= io_in_r_bypass_6_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_0_data_29 <= io_in_r_bypass_7_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_0_load_store_29 <= io_in_r_bypass_7_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_0_df_is_ws_29 <= io_in_r_bypass_7_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_0_stall_29 <= io_in_r_bypass_7_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_1_data_29 <= io_in_r_bypass_7_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_1_load_store_29 <= io_in_r_bypass_7_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_1_df_is_ws_29 <= io_in_r_bypass_7_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_1_stall_29 <= io_in_r_bypass_7_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_2_data_29 <= io_in_r_bypass_7_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_2_load_store_29 <= io_in_r_bypass_7_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_2_df_is_ws_29 <= io_in_r_bypass_7_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_2_stall_29 <= io_in_r_bypass_7_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_3_data_29 <= io_in_r_bypass_7_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_3_load_store_29 <= io_in_r_bypass_7_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_3_df_is_ws_29 <= io_in_r_bypass_7_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_3_stall_29 <= io_in_r_bypass_7_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_0_data_29 <= io_in_r_bypass_8_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_0_load_store_29 <= io_in_r_bypass_8_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_0_df_is_ws_29 <= io_in_r_bypass_8_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_0_stall_29 <= io_in_r_bypass_8_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_1_data_29 <= io_in_r_bypass_8_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_1_load_store_29 <= io_in_r_bypass_8_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_1_df_is_ws_29 <= io_in_r_bypass_8_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_1_stall_29 <= io_in_r_bypass_8_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_2_data_29 <= io_in_r_bypass_8_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_2_load_store_29 <= io_in_r_bypass_8_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_2_df_is_ws_29 <= io_in_r_bypass_8_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_2_stall_29 <= io_in_r_bypass_8_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_3_data_29 <= io_in_r_bypass_8_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_3_load_store_29 <= io_in_r_bypass_8_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_3_df_is_ws_29 <= io_in_r_bypass_8_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_3_stall_29 <= io_in_r_bypass_8_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_0_data_29 <= io_in_r_bypass_9_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_0_load_store_29 <= io_in_r_bypass_9_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_0_df_is_ws_29 <= io_in_r_bypass_9_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_0_stall_29 <= io_in_r_bypass_9_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_1_data_29 <= io_in_r_bypass_9_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_1_load_store_29 <= io_in_r_bypass_9_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_1_df_is_ws_29 <= io_in_r_bypass_9_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_1_stall_29 <= io_in_r_bypass_9_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_2_data_29 <= io_in_r_bypass_9_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_2_load_store_29 <= io_in_r_bypass_9_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_2_df_is_ws_29 <= io_in_r_bypass_9_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_2_stall_29 <= io_in_r_bypass_9_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_3_data_29 <= io_in_r_bypass_9_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_3_load_store_29 <= io_in_r_bypass_9_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_3_df_is_ws_29 <= io_in_r_bypass_9_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_3_stall_29 <= io_in_r_bypass_9_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_0_data_29 <= io_in_r_bypass_10_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_0_load_store_29 <= io_in_r_bypass_10_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_0_df_is_ws_29 <= io_in_r_bypass_10_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_0_stall_29 <= io_in_r_bypass_10_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_1_data_29 <= io_in_r_bypass_10_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_1_load_store_29 <= io_in_r_bypass_10_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_1_df_is_ws_29 <= io_in_r_bypass_10_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_1_stall_29 <= io_in_r_bypass_10_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_2_data_29 <= io_in_r_bypass_10_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_2_load_store_29 <= io_in_r_bypass_10_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_2_df_is_ws_29 <= io_in_r_bypass_10_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_2_stall_29 <= io_in_r_bypass_10_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_3_data_29 <= io_in_r_bypass_10_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_3_load_store_29 <= io_in_r_bypass_10_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_3_df_is_ws_29 <= io_in_r_bypass_10_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_3_stall_29 <= io_in_r_bypass_10_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_0_data_29 <= io_in_r_bypass_11_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_0_load_store_29 <= io_in_r_bypass_11_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_0_df_is_ws_29 <= io_in_r_bypass_11_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_0_stall_29 <= io_in_r_bypass_11_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_1_data_29 <= io_in_r_bypass_11_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_1_load_store_29 <= io_in_r_bypass_11_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_1_df_is_ws_29 <= io_in_r_bypass_11_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_1_stall_29 <= io_in_r_bypass_11_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_2_data_29 <= io_in_r_bypass_11_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_2_load_store_29 <= io_in_r_bypass_11_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_2_df_is_ws_29 <= io_in_r_bypass_11_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_2_stall_29 <= io_in_r_bypass_11_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_3_data_29 <= io_in_r_bypass_11_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_3_load_store_29 <= io_in_r_bypass_11_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_3_df_is_ws_29 <= io_in_r_bypass_11_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_3_stall_29 <= io_in_r_bypass_11_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_0_data_29 <= io_in_r_bypass_12_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_0_load_store_29 <= io_in_r_bypass_12_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_0_df_is_ws_29 <= io_in_r_bypass_12_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_0_stall_29 <= io_in_r_bypass_12_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_1_data_29 <= io_in_r_bypass_12_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_1_load_store_29 <= io_in_r_bypass_12_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_1_df_is_ws_29 <= io_in_r_bypass_12_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_1_stall_29 <= io_in_r_bypass_12_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_2_data_29 <= io_in_r_bypass_12_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_2_load_store_29 <= io_in_r_bypass_12_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_2_df_is_ws_29 <= io_in_r_bypass_12_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_2_stall_29 <= io_in_r_bypass_12_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_3_data_29 <= io_in_r_bypass_12_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_3_load_store_29 <= io_in_r_bypass_12_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_3_df_is_ws_29 <= io_in_r_bypass_12_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_3_stall_29 <= io_in_r_bypass_12_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_0_data_29 <= io_in_r_bypass_13_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_0_load_store_29 <= io_in_r_bypass_13_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_0_df_is_ws_29 <= io_in_r_bypass_13_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_0_stall_29 <= io_in_r_bypass_13_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_1_data_29 <= io_in_r_bypass_13_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_1_load_store_29 <= io_in_r_bypass_13_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_1_df_is_ws_29 <= io_in_r_bypass_13_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_1_stall_29 <= io_in_r_bypass_13_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_2_data_29 <= io_in_r_bypass_13_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_2_load_store_29 <= io_in_r_bypass_13_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_2_df_is_ws_29 <= io_in_r_bypass_13_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_2_stall_29 <= io_in_r_bypass_13_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_3_data_29 <= io_in_r_bypass_13_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_3_load_store_29 <= io_in_r_bypass_13_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_3_df_is_ws_29 <= io_in_r_bypass_13_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_3_stall_29 <= io_in_r_bypass_13_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_0_data_29 <= io_in_r_bypass_14_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_0_load_store_29 <= io_in_r_bypass_14_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_0_df_is_ws_29 <= io_in_r_bypass_14_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_0_stall_29 <= io_in_r_bypass_14_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_1_data_29 <= io_in_r_bypass_14_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_1_load_store_29 <= io_in_r_bypass_14_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_1_df_is_ws_29 <= io_in_r_bypass_14_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_1_stall_29 <= io_in_r_bypass_14_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_2_data_29 <= io_in_r_bypass_14_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_2_load_store_29 <= io_in_r_bypass_14_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_2_df_is_ws_29 <= io_in_r_bypass_14_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_2_stall_29 <= io_in_r_bypass_14_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_3_data_29 <= io_in_r_bypass_14_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_3_load_store_29 <= io_in_r_bypass_14_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_3_df_is_ws_29 <= io_in_r_bypass_14_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_3_stall_29 <= io_in_r_bypass_14_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_0_data_29 <= io_in_r_bypass_15_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_0_load_store_29 <= io_in_r_bypass_15_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_0_df_is_ws_29 <= io_in_r_bypass_15_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_0_stall_29 <= io_in_r_bypass_15_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_1_data_29 <= io_in_r_bypass_15_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_1_load_store_29 <= io_in_r_bypass_15_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_1_df_is_ws_29 <= io_in_r_bypass_15_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_1_stall_29 <= io_in_r_bypass_15_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_2_data_29 <= io_in_r_bypass_15_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_2_load_store_29 <= io_in_r_bypass_15_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_2_df_is_ws_29 <= io_in_r_bypass_15_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_2_stall_29 <= io_in_r_bypass_15_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_3_data_29 <= io_in_r_bypass_15_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_3_load_store_29 <= io_in_r_bypass_15_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_3_df_is_ws_29 <= io_in_r_bypass_15_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_3_stall_29 <= io_in_r_bypass_15_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_0_data_29 <= io_in_r_bypass_16_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_0_load_store_29 <= io_in_r_bypass_16_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_0_df_is_ws_29 <= io_in_r_bypass_16_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_0_stall_29 <= io_in_r_bypass_16_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_1_data_29 <= io_in_r_bypass_16_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_1_load_store_29 <= io_in_r_bypass_16_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_1_df_is_ws_29 <= io_in_r_bypass_16_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_1_stall_29 <= io_in_r_bypass_16_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_2_data_29 <= io_in_r_bypass_16_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_2_load_store_29 <= io_in_r_bypass_16_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_2_df_is_ws_29 <= io_in_r_bypass_16_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_2_stall_29 <= io_in_r_bypass_16_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_3_data_29 <= io_in_r_bypass_16_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_3_load_store_29 <= io_in_r_bypass_16_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_3_df_is_ws_29 <= io_in_r_bypass_16_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_3_stall_29 <= io_in_r_bypass_16_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_0_data_29 <= io_in_r_bypass_17_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_0_load_store_29 <= io_in_r_bypass_17_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_0_df_is_ws_29 <= io_in_r_bypass_17_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_0_stall_29 <= io_in_r_bypass_17_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_1_data_29 <= io_in_r_bypass_17_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_1_load_store_29 <= io_in_r_bypass_17_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_1_df_is_ws_29 <= io_in_r_bypass_17_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_1_stall_29 <= io_in_r_bypass_17_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_2_data_29 <= io_in_r_bypass_17_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_2_load_store_29 <= io_in_r_bypass_17_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_2_df_is_ws_29 <= io_in_r_bypass_17_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_2_stall_29 <= io_in_r_bypass_17_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_3_data_29 <= io_in_r_bypass_17_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_3_load_store_29 <= io_in_r_bypass_17_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_3_df_is_ws_29 <= io_in_r_bypass_17_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_3_stall_29 <= io_in_r_bypass_17_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_0_data_29 <= io_in_r_bypass_18_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_0_load_store_29 <= io_in_r_bypass_18_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_0_df_is_ws_29 <= io_in_r_bypass_18_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_0_stall_29 <= io_in_r_bypass_18_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_1_data_29 <= io_in_r_bypass_18_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_1_load_store_29 <= io_in_r_bypass_18_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_1_df_is_ws_29 <= io_in_r_bypass_18_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_1_stall_29 <= io_in_r_bypass_18_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_2_data_29 <= io_in_r_bypass_18_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_2_load_store_29 <= io_in_r_bypass_18_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_2_df_is_ws_29 <= io_in_r_bypass_18_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_2_stall_29 <= io_in_r_bypass_18_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_3_data_29 <= io_in_r_bypass_18_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_3_load_store_29 <= io_in_r_bypass_18_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_3_df_is_ws_29 <= io_in_r_bypass_18_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_3_stall_29 <= io_in_r_bypass_18_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_0_data_29 <= io_in_r_bypass_19_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_0_load_store_29 <= io_in_r_bypass_19_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_0_df_is_ws_29 <= io_in_r_bypass_19_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_0_stall_29 <= io_in_r_bypass_19_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_1_data_29 <= io_in_r_bypass_19_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_1_load_store_29 <= io_in_r_bypass_19_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_1_df_is_ws_29 <= io_in_r_bypass_19_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_1_stall_29 <= io_in_r_bypass_19_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_2_data_29 <= io_in_r_bypass_19_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_2_load_store_29 <= io_in_r_bypass_19_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_2_df_is_ws_29 <= io_in_r_bypass_19_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_2_stall_29 <= io_in_r_bypass_19_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_3_data_29 <= io_in_r_bypass_19_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_3_load_store_29 <= io_in_r_bypass_19_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_3_df_is_ws_29 <= io_in_r_bypass_19_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_3_stall_29 <= io_in_r_bypass_19_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_0_data_29 <= io_in_r_bypass_20_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_0_load_store_29 <= io_in_r_bypass_20_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_0_df_is_ws_29 <= io_in_r_bypass_20_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_0_stall_29 <= io_in_r_bypass_20_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_1_data_29 <= io_in_r_bypass_20_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_1_load_store_29 <= io_in_r_bypass_20_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_1_df_is_ws_29 <= io_in_r_bypass_20_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_1_stall_29 <= io_in_r_bypass_20_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_2_data_29 <= io_in_r_bypass_20_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_2_load_store_29 <= io_in_r_bypass_20_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_2_df_is_ws_29 <= io_in_r_bypass_20_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_2_stall_29 <= io_in_r_bypass_20_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_3_data_29 <= io_in_r_bypass_20_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_3_load_store_29 <= io_in_r_bypass_20_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_3_df_is_ws_29 <= io_in_r_bypass_20_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_3_stall_29 <= io_in_r_bypass_20_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_0_data_29 <= io_in_r_bypass_21_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_0_load_store_29 <= io_in_r_bypass_21_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_0_df_is_ws_29 <= io_in_r_bypass_21_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_0_stall_29 <= io_in_r_bypass_21_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_1_data_29 <= io_in_r_bypass_21_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_1_load_store_29 <= io_in_r_bypass_21_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_1_df_is_ws_29 <= io_in_r_bypass_21_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_1_stall_29 <= io_in_r_bypass_21_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_2_data_29 <= io_in_r_bypass_21_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_2_load_store_29 <= io_in_r_bypass_21_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_2_df_is_ws_29 <= io_in_r_bypass_21_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_2_stall_29 <= io_in_r_bypass_21_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_3_data_29 <= io_in_r_bypass_21_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_3_load_store_29 <= io_in_r_bypass_21_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_3_df_is_ws_29 <= io_in_r_bypass_21_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_3_stall_29 <= io_in_r_bypass_21_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_0_data_29 <= io_in_r_bypass_22_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_0_load_store_29 <= io_in_r_bypass_22_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_0_df_is_ws_29 <= io_in_r_bypass_22_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_0_stall_29 <= io_in_r_bypass_22_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_1_data_29 <= io_in_r_bypass_22_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_1_load_store_29 <= io_in_r_bypass_22_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_1_df_is_ws_29 <= io_in_r_bypass_22_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_1_stall_29 <= io_in_r_bypass_22_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_2_data_29 <= io_in_r_bypass_22_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_2_load_store_29 <= io_in_r_bypass_22_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_2_df_is_ws_29 <= io_in_r_bypass_22_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_2_stall_29 <= io_in_r_bypass_22_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_3_data_29 <= io_in_r_bypass_22_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_3_load_store_29 <= io_in_r_bypass_22_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_3_df_is_ws_29 <= io_in_r_bypass_22_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_3_stall_29 <= io_in_r_bypass_22_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_0_data_29 <= io_in_r_bypass_23_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_0_load_store_29 <= io_in_r_bypass_23_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_0_df_is_ws_29 <= io_in_r_bypass_23_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_0_stall_29 <= io_in_r_bypass_23_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_1_data_29 <= io_in_r_bypass_23_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_1_load_store_29 <= io_in_r_bypass_23_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_1_df_is_ws_29 <= io_in_r_bypass_23_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_1_stall_29 <= io_in_r_bypass_23_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_2_data_29 <= io_in_r_bypass_23_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_2_load_store_29 <= io_in_r_bypass_23_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_2_df_is_ws_29 <= io_in_r_bypass_23_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_2_stall_29 <= io_in_r_bypass_23_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_3_data_29 <= io_in_r_bypass_23_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_3_load_store_29 <= io_in_r_bypass_23_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_3_df_is_ws_29 <= io_in_r_bypass_23_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_3_stall_29 <= io_in_r_bypass_23_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_0_data_29 <= io_in_r_bypass_24_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_0_load_store_29 <= io_in_r_bypass_24_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_0_df_is_ws_29 <= io_in_r_bypass_24_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_0_stall_29 <= io_in_r_bypass_24_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_1_data_29 <= io_in_r_bypass_24_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_1_load_store_29 <= io_in_r_bypass_24_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_1_df_is_ws_29 <= io_in_r_bypass_24_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_1_stall_29 <= io_in_r_bypass_24_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_2_data_29 <= io_in_r_bypass_24_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_2_load_store_29 <= io_in_r_bypass_24_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_2_df_is_ws_29 <= io_in_r_bypass_24_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_2_stall_29 <= io_in_r_bypass_24_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_3_data_29 <= io_in_r_bypass_24_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_3_load_store_29 <= io_in_r_bypass_24_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_3_df_is_ws_29 <= io_in_r_bypass_24_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_3_stall_29 <= io_in_r_bypass_24_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_0_data_29 <= io_in_r_bypass_25_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_0_load_store_29 <= io_in_r_bypass_25_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_0_df_is_ws_29 <= io_in_r_bypass_25_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_0_stall_29 <= io_in_r_bypass_25_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_1_data_29 <= io_in_r_bypass_25_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_1_load_store_29 <= io_in_r_bypass_25_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_1_df_is_ws_29 <= io_in_r_bypass_25_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_1_stall_29 <= io_in_r_bypass_25_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_2_data_29 <= io_in_r_bypass_25_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_2_load_store_29 <= io_in_r_bypass_25_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_2_df_is_ws_29 <= io_in_r_bypass_25_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_2_stall_29 <= io_in_r_bypass_25_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_3_data_29 <= io_in_r_bypass_25_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_3_load_store_29 <= io_in_r_bypass_25_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_3_df_is_ws_29 <= io_in_r_bypass_25_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_3_stall_29 <= io_in_r_bypass_25_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_0_data_29 <= io_in_r_bypass_26_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_0_load_store_29 <= io_in_r_bypass_26_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_0_df_is_ws_29 <= io_in_r_bypass_26_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_0_stall_29 <= io_in_r_bypass_26_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_1_data_29 <= io_in_r_bypass_26_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_1_load_store_29 <= io_in_r_bypass_26_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_1_df_is_ws_29 <= io_in_r_bypass_26_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_1_stall_29 <= io_in_r_bypass_26_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_2_data_29 <= io_in_r_bypass_26_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_2_load_store_29 <= io_in_r_bypass_26_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_2_df_is_ws_29 <= io_in_r_bypass_26_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_2_stall_29 <= io_in_r_bypass_26_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_3_data_29 <= io_in_r_bypass_26_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_3_load_store_29 <= io_in_r_bypass_26_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_3_df_is_ws_29 <= io_in_r_bypass_26_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_3_stall_29 <= io_in_r_bypass_26_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_0_data_29 <= io_in_r_bypass_27_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_0_load_store_29 <= io_in_r_bypass_27_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_0_df_is_ws_29 <= io_in_r_bypass_27_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_0_stall_29 <= io_in_r_bypass_27_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_1_data_29 <= io_in_r_bypass_27_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_1_load_store_29 <= io_in_r_bypass_27_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_1_df_is_ws_29 <= io_in_r_bypass_27_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_1_stall_29 <= io_in_r_bypass_27_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_2_data_29 <= io_in_r_bypass_27_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_2_load_store_29 <= io_in_r_bypass_27_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_2_df_is_ws_29 <= io_in_r_bypass_27_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_2_stall_29 <= io_in_r_bypass_27_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_3_data_29 <= io_in_r_bypass_27_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_3_load_store_29 <= io_in_r_bypass_27_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_3_df_is_ws_29 <= io_in_r_bypass_27_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_3_stall_29 <= io_in_r_bypass_27_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_0_data_29 <= io_in_r_bypass_28_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_0_load_store_29 <= io_in_r_bypass_28_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_0_df_is_ws_29 <= io_in_r_bypass_28_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_0_stall_29 <= io_in_r_bypass_28_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_1_data_29 <= io_in_r_bypass_28_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_1_load_store_29 <= io_in_r_bypass_28_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_1_df_is_ws_29 <= io_in_r_bypass_28_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_1_stall_29 <= io_in_r_bypass_28_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_2_data_29 <= io_in_r_bypass_28_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_2_load_store_29 <= io_in_r_bypass_28_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_2_df_is_ws_29 <= io_in_r_bypass_28_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_2_stall_29 <= io_in_r_bypass_28_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_3_data_29 <= io_in_r_bypass_28_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_3_load_store_29 <= io_in_r_bypass_28_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_3_df_is_ws_29 <= io_in_r_bypass_28_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_3_stall_29 <= io_in_r_bypass_28_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_0_data_29 <= io_in_r_bypass_29_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_0_load_store_29 <= io_in_r_bypass_29_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_0_df_is_ws_29 <= io_in_r_bypass_29_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_0_stall_29 <= io_in_r_bypass_29_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_1_data_29 <= io_in_r_bypass_29_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_1_load_store_29 <= io_in_r_bypass_29_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_1_df_is_ws_29 <= io_in_r_bypass_29_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_1_stall_29 <= io_in_r_bypass_29_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_2_data_29 <= io_in_r_bypass_29_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_2_load_store_29 <= io_in_r_bypass_29_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_2_df_is_ws_29 <= io_in_r_bypass_29_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_2_stall_29 <= io_in_r_bypass_29_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_3_data_29 <= io_in_r_bypass_29_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_3_load_store_29 <= io_in_r_bypass_29_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_3_df_is_ws_29 <= io_in_r_bypass_29_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_3_stall_29 <= io_in_r_bypass_29_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_0_data_29 <= io_in_r_bypass_30_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_0_load_store_29 <= io_in_r_bypass_30_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_0_df_is_ws_29 <= io_in_r_bypass_30_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_0_stall_29 <= io_in_r_bypass_30_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_1_data_29 <= io_in_r_bypass_30_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_1_load_store_29 <= io_in_r_bypass_30_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_1_df_is_ws_29 <= io_in_r_bypass_30_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_1_stall_29 <= io_in_r_bypass_30_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_2_data_29 <= io_in_r_bypass_30_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_2_load_store_29 <= io_in_r_bypass_30_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_2_df_is_ws_29 <= io_in_r_bypass_30_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_2_stall_29 <= io_in_r_bypass_30_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_3_data_29 <= io_in_r_bypass_30_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_3_load_store_29 <= io_in_r_bypass_30_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_3_df_is_ws_29 <= io_in_r_bypass_30_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_3_stall_29 <= io_in_r_bypass_30_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_0_data_29 <= io_in_r_bypass_31_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_0_load_store_29 <= io_in_r_bypass_31_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_0_df_is_ws_29 <= io_in_r_bypass_31_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_0_stall_29 <= io_in_r_bypass_31_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_1_data_29 <= io_in_r_bypass_31_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_1_load_store_29 <= io_in_r_bypass_31_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_1_df_is_ws_29 <= io_in_r_bypass_31_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_1_stall_29 <= io_in_r_bypass_31_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_2_data_29 <= io_in_r_bypass_31_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_2_load_store_29 <= io_in_r_bypass_31_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_2_df_is_ws_29 <= io_in_r_bypass_31_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_2_stall_29 <= io_in_r_bypass_31_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_3_data_29 <= io_in_r_bypass_31_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_3_load_store_29 <= io_in_r_bypass_31_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_3_df_is_ws_29 <= io_in_r_bypass_31_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_3_stall_29 <= io_in_r_bypass_31_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_0_data_30 <= io_in_r_bypass_0_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_0_load_store_30 <= io_in_r_bypass_0_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_0_df_is_ws_30 <= io_in_r_bypass_0_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_0_stall_30 <= io_in_r_bypass_0_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_1_data_30 <= io_in_r_bypass_0_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_1_load_store_30 <= io_in_r_bypass_0_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_1_df_is_ws_30 <= io_in_r_bypass_0_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_1_stall_30 <= io_in_r_bypass_0_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_2_data_30 <= io_in_r_bypass_0_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_2_load_store_30 <= io_in_r_bypass_0_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_2_df_is_ws_30 <= io_in_r_bypass_0_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_2_stall_30 <= io_in_r_bypass_0_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_3_data_30 <= io_in_r_bypass_0_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_3_load_store_30 <= io_in_r_bypass_0_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_3_df_is_ws_30 <= io_in_r_bypass_0_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_3_stall_30 <= io_in_r_bypass_0_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_0_data_30 <= io_in_r_bypass_1_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_0_load_store_30 <= io_in_r_bypass_1_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_0_df_is_ws_30 <= io_in_r_bypass_1_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_0_stall_30 <= io_in_r_bypass_1_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_1_data_30 <= io_in_r_bypass_1_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_1_load_store_30 <= io_in_r_bypass_1_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_1_df_is_ws_30 <= io_in_r_bypass_1_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_1_stall_30 <= io_in_r_bypass_1_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_2_data_30 <= io_in_r_bypass_1_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_2_load_store_30 <= io_in_r_bypass_1_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_2_df_is_ws_30 <= io_in_r_bypass_1_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_2_stall_30 <= io_in_r_bypass_1_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_3_data_30 <= io_in_r_bypass_1_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_3_load_store_30 <= io_in_r_bypass_1_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_3_df_is_ws_30 <= io_in_r_bypass_1_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_3_stall_30 <= io_in_r_bypass_1_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_0_data_30 <= io_in_r_bypass_2_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_0_load_store_30 <= io_in_r_bypass_2_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_0_df_is_ws_30 <= io_in_r_bypass_2_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_0_stall_30 <= io_in_r_bypass_2_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_1_data_30 <= io_in_r_bypass_2_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_1_load_store_30 <= io_in_r_bypass_2_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_1_df_is_ws_30 <= io_in_r_bypass_2_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_1_stall_30 <= io_in_r_bypass_2_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_2_data_30 <= io_in_r_bypass_2_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_2_load_store_30 <= io_in_r_bypass_2_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_2_df_is_ws_30 <= io_in_r_bypass_2_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_2_stall_30 <= io_in_r_bypass_2_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_3_data_30 <= io_in_r_bypass_2_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_3_load_store_30 <= io_in_r_bypass_2_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_3_df_is_ws_30 <= io_in_r_bypass_2_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_2_3_stall_30 <= io_in_r_bypass_2_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_0_data_30 <= io_in_r_bypass_3_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_0_load_store_30 <= io_in_r_bypass_3_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_0_df_is_ws_30 <= io_in_r_bypass_3_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_0_stall_30 <= io_in_r_bypass_3_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_1_data_30 <= io_in_r_bypass_3_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_1_load_store_30 <= io_in_r_bypass_3_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_1_df_is_ws_30 <= io_in_r_bypass_3_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_1_stall_30 <= io_in_r_bypass_3_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_2_data_30 <= io_in_r_bypass_3_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_2_load_store_30 <= io_in_r_bypass_3_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_2_df_is_ws_30 <= io_in_r_bypass_3_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_2_stall_30 <= io_in_r_bypass_3_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_3_data_30 <= io_in_r_bypass_3_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_3_load_store_30 <= io_in_r_bypass_3_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_3_df_is_ws_30 <= io_in_r_bypass_3_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_3_3_stall_30 <= io_in_r_bypass_3_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_0_data_30 <= io_in_r_bypass_4_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_0_load_store_30 <= io_in_r_bypass_4_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_0_df_is_ws_30 <= io_in_r_bypass_4_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_0_stall_30 <= io_in_r_bypass_4_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_1_data_30 <= io_in_r_bypass_4_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_1_load_store_30 <= io_in_r_bypass_4_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_1_df_is_ws_30 <= io_in_r_bypass_4_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_1_stall_30 <= io_in_r_bypass_4_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_2_data_30 <= io_in_r_bypass_4_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_2_load_store_30 <= io_in_r_bypass_4_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_2_df_is_ws_30 <= io_in_r_bypass_4_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_2_stall_30 <= io_in_r_bypass_4_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_3_data_30 <= io_in_r_bypass_4_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_3_load_store_30 <= io_in_r_bypass_4_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_3_df_is_ws_30 <= io_in_r_bypass_4_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_4_3_stall_30 <= io_in_r_bypass_4_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_0_data_30 <= io_in_r_bypass_5_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_0_load_store_30 <= io_in_r_bypass_5_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_0_df_is_ws_30 <= io_in_r_bypass_5_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_0_stall_30 <= io_in_r_bypass_5_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_1_data_30 <= io_in_r_bypass_5_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_1_load_store_30 <= io_in_r_bypass_5_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_1_df_is_ws_30 <= io_in_r_bypass_5_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_1_stall_30 <= io_in_r_bypass_5_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_2_data_30 <= io_in_r_bypass_5_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_2_load_store_30 <= io_in_r_bypass_5_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_2_df_is_ws_30 <= io_in_r_bypass_5_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_2_stall_30 <= io_in_r_bypass_5_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_3_data_30 <= io_in_r_bypass_5_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_3_load_store_30 <= io_in_r_bypass_5_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_3_df_is_ws_30 <= io_in_r_bypass_5_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_5_3_stall_30 <= io_in_r_bypass_5_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_0_data_30 <= io_in_r_bypass_6_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_0_load_store_30 <= io_in_r_bypass_6_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_0_df_is_ws_30 <= io_in_r_bypass_6_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_0_stall_30 <= io_in_r_bypass_6_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_1_data_30 <= io_in_r_bypass_6_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_1_load_store_30 <= io_in_r_bypass_6_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_1_df_is_ws_30 <= io_in_r_bypass_6_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_1_stall_30 <= io_in_r_bypass_6_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_2_data_30 <= io_in_r_bypass_6_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_2_load_store_30 <= io_in_r_bypass_6_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_2_df_is_ws_30 <= io_in_r_bypass_6_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_2_stall_30 <= io_in_r_bypass_6_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_3_data_30 <= io_in_r_bypass_6_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_3_load_store_30 <= io_in_r_bypass_6_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_3_df_is_ws_30 <= io_in_r_bypass_6_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_6_3_stall_30 <= io_in_r_bypass_6_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_0_data_30 <= io_in_r_bypass_7_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_0_load_store_30 <= io_in_r_bypass_7_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_0_df_is_ws_30 <= io_in_r_bypass_7_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_0_stall_30 <= io_in_r_bypass_7_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_1_data_30 <= io_in_r_bypass_7_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_1_load_store_30 <= io_in_r_bypass_7_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_1_df_is_ws_30 <= io_in_r_bypass_7_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_1_stall_30 <= io_in_r_bypass_7_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_2_data_30 <= io_in_r_bypass_7_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_2_load_store_30 <= io_in_r_bypass_7_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_2_df_is_ws_30 <= io_in_r_bypass_7_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_2_stall_30 <= io_in_r_bypass_7_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_3_data_30 <= io_in_r_bypass_7_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_3_load_store_30 <= io_in_r_bypass_7_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_3_df_is_ws_30 <= io_in_r_bypass_7_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_7_3_stall_30 <= io_in_r_bypass_7_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_0_data_30 <= io_in_r_bypass_8_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_0_load_store_30 <= io_in_r_bypass_8_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_0_df_is_ws_30 <= io_in_r_bypass_8_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_0_stall_30 <= io_in_r_bypass_8_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_1_data_30 <= io_in_r_bypass_8_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_1_load_store_30 <= io_in_r_bypass_8_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_1_df_is_ws_30 <= io_in_r_bypass_8_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_1_stall_30 <= io_in_r_bypass_8_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_2_data_30 <= io_in_r_bypass_8_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_2_load_store_30 <= io_in_r_bypass_8_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_2_df_is_ws_30 <= io_in_r_bypass_8_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_2_stall_30 <= io_in_r_bypass_8_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_3_data_30 <= io_in_r_bypass_8_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_3_load_store_30 <= io_in_r_bypass_8_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_3_df_is_ws_30 <= io_in_r_bypass_8_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_8_3_stall_30 <= io_in_r_bypass_8_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_0_data_30 <= io_in_r_bypass_9_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_0_load_store_30 <= io_in_r_bypass_9_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_0_df_is_ws_30 <= io_in_r_bypass_9_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_0_stall_30 <= io_in_r_bypass_9_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_1_data_30 <= io_in_r_bypass_9_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_1_load_store_30 <= io_in_r_bypass_9_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_1_df_is_ws_30 <= io_in_r_bypass_9_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_1_stall_30 <= io_in_r_bypass_9_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_2_data_30 <= io_in_r_bypass_9_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_2_load_store_30 <= io_in_r_bypass_9_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_2_df_is_ws_30 <= io_in_r_bypass_9_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_2_stall_30 <= io_in_r_bypass_9_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_3_data_30 <= io_in_r_bypass_9_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_3_load_store_30 <= io_in_r_bypass_9_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_3_df_is_ws_30 <= io_in_r_bypass_9_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_9_3_stall_30 <= io_in_r_bypass_9_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_0_data_30 <= io_in_r_bypass_10_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_0_load_store_30 <= io_in_r_bypass_10_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_0_df_is_ws_30 <= io_in_r_bypass_10_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_0_stall_30 <= io_in_r_bypass_10_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_1_data_30 <= io_in_r_bypass_10_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_1_load_store_30 <= io_in_r_bypass_10_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_1_df_is_ws_30 <= io_in_r_bypass_10_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_1_stall_30 <= io_in_r_bypass_10_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_2_data_30 <= io_in_r_bypass_10_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_2_load_store_30 <= io_in_r_bypass_10_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_2_df_is_ws_30 <= io_in_r_bypass_10_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_2_stall_30 <= io_in_r_bypass_10_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_3_data_30 <= io_in_r_bypass_10_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_3_load_store_30 <= io_in_r_bypass_10_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_3_df_is_ws_30 <= io_in_r_bypass_10_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_10_3_stall_30 <= io_in_r_bypass_10_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_0_data_30 <= io_in_r_bypass_11_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_0_load_store_30 <= io_in_r_bypass_11_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_0_df_is_ws_30 <= io_in_r_bypass_11_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_0_stall_30 <= io_in_r_bypass_11_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_1_data_30 <= io_in_r_bypass_11_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_1_load_store_30 <= io_in_r_bypass_11_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_1_df_is_ws_30 <= io_in_r_bypass_11_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_1_stall_30 <= io_in_r_bypass_11_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_2_data_30 <= io_in_r_bypass_11_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_2_load_store_30 <= io_in_r_bypass_11_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_2_df_is_ws_30 <= io_in_r_bypass_11_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_2_stall_30 <= io_in_r_bypass_11_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_3_data_30 <= io_in_r_bypass_11_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_3_load_store_30 <= io_in_r_bypass_11_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_3_df_is_ws_30 <= io_in_r_bypass_11_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_11_3_stall_30 <= io_in_r_bypass_11_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_0_data_30 <= io_in_r_bypass_12_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_0_load_store_30 <= io_in_r_bypass_12_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_0_df_is_ws_30 <= io_in_r_bypass_12_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_0_stall_30 <= io_in_r_bypass_12_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_1_data_30 <= io_in_r_bypass_12_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_1_load_store_30 <= io_in_r_bypass_12_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_1_df_is_ws_30 <= io_in_r_bypass_12_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_1_stall_30 <= io_in_r_bypass_12_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_2_data_30 <= io_in_r_bypass_12_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_2_load_store_30 <= io_in_r_bypass_12_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_2_df_is_ws_30 <= io_in_r_bypass_12_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_2_stall_30 <= io_in_r_bypass_12_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_3_data_30 <= io_in_r_bypass_12_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_3_load_store_30 <= io_in_r_bypass_12_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_3_df_is_ws_30 <= io_in_r_bypass_12_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_12_3_stall_30 <= io_in_r_bypass_12_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_0_data_30 <= io_in_r_bypass_13_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_0_load_store_30 <= io_in_r_bypass_13_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_0_df_is_ws_30 <= io_in_r_bypass_13_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_0_stall_30 <= io_in_r_bypass_13_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_1_data_30 <= io_in_r_bypass_13_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_1_load_store_30 <= io_in_r_bypass_13_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_1_df_is_ws_30 <= io_in_r_bypass_13_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_1_stall_30 <= io_in_r_bypass_13_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_2_data_30 <= io_in_r_bypass_13_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_2_load_store_30 <= io_in_r_bypass_13_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_2_df_is_ws_30 <= io_in_r_bypass_13_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_2_stall_30 <= io_in_r_bypass_13_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_3_data_30 <= io_in_r_bypass_13_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_3_load_store_30 <= io_in_r_bypass_13_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_3_df_is_ws_30 <= io_in_r_bypass_13_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_13_3_stall_30 <= io_in_r_bypass_13_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_0_data_30 <= io_in_r_bypass_14_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_0_load_store_30 <= io_in_r_bypass_14_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_0_df_is_ws_30 <= io_in_r_bypass_14_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_0_stall_30 <= io_in_r_bypass_14_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_1_data_30 <= io_in_r_bypass_14_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_1_load_store_30 <= io_in_r_bypass_14_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_1_df_is_ws_30 <= io_in_r_bypass_14_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_1_stall_30 <= io_in_r_bypass_14_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_2_data_30 <= io_in_r_bypass_14_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_2_load_store_30 <= io_in_r_bypass_14_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_2_df_is_ws_30 <= io_in_r_bypass_14_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_2_stall_30 <= io_in_r_bypass_14_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_3_data_30 <= io_in_r_bypass_14_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_3_load_store_30 <= io_in_r_bypass_14_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_3_df_is_ws_30 <= io_in_r_bypass_14_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_14_3_stall_30 <= io_in_r_bypass_14_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_0_data_30 <= io_in_r_bypass_15_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_0_load_store_30 <= io_in_r_bypass_15_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_0_df_is_ws_30 <= io_in_r_bypass_15_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_0_stall_30 <= io_in_r_bypass_15_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_1_data_30 <= io_in_r_bypass_15_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_1_load_store_30 <= io_in_r_bypass_15_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_1_df_is_ws_30 <= io_in_r_bypass_15_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_1_stall_30 <= io_in_r_bypass_15_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_2_data_30 <= io_in_r_bypass_15_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_2_load_store_30 <= io_in_r_bypass_15_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_2_df_is_ws_30 <= io_in_r_bypass_15_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_2_stall_30 <= io_in_r_bypass_15_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_3_data_30 <= io_in_r_bypass_15_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_3_load_store_30 <= io_in_r_bypass_15_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_3_df_is_ws_30 <= io_in_r_bypass_15_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_15_3_stall_30 <= io_in_r_bypass_15_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_0_data_30 <= io_in_r_bypass_16_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_0_load_store_30 <= io_in_r_bypass_16_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_0_df_is_ws_30 <= io_in_r_bypass_16_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_0_stall_30 <= io_in_r_bypass_16_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_1_data_30 <= io_in_r_bypass_16_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_1_load_store_30 <= io_in_r_bypass_16_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_1_df_is_ws_30 <= io_in_r_bypass_16_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_1_stall_30 <= io_in_r_bypass_16_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_2_data_30 <= io_in_r_bypass_16_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_2_load_store_30 <= io_in_r_bypass_16_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_2_df_is_ws_30 <= io_in_r_bypass_16_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_2_stall_30 <= io_in_r_bypass_16_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_3_data_30 <= io_in_r_bypass_16_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_3_load_store_30 <= io_in_r_bypass_16_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_3_df_is_ws_30 <= io_in_r_bypass_16_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_16_3_stall_30 <= io_in_r_bypass_16_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_0_data_30 <= io_in_r_bypass_17_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_0_load_store_30 <= io_in_r_bypass_17_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_0_df_is_ws_30 <= io_in_r_bypass_17_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_0_stall_30 <= io_in_r_bypass_17_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_1_data_30 <= io_in_r_bypass_17_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_1_load_store_30 <= io_in_r_bypass_17_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_1_df_is_ws_30 <= io_in_r_bypass_17_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_1_stall_30 <= io_in_r_bypass_17_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_2_data_30 <= io_in_r_bypass_17_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_2_load_store_30 <= io_in_r_bypass_17_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_2_df_is_ws_30 <= io_in_r_bypass_17_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_2_stall_30 <= io_in_r_bypass_17_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_3_data_30 <= io_in_r_bypass_17_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_3_load_store_30 <= io_in_r_bypass_17_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_3_df_is_ws_30 <= io_in_r_bypass_17_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_17_3_stall_30 <= io_in_r_bypass_17_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_0_data_30 <= io_in_r_bypass_18_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_0_load_store_30 <= io_in_r_bypass_18_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_0_df_is_ws_30 <= io_in_r_bypass_18_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_0_stall_30 <= io_in_r_bypass_18_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_1_data_30 <= io_in_r_bypass_18_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_1_load_store_30 <= io_in_r_bypass_18_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_1_df_is_ws_30 <= io_in_r_bypass_18_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_1_stall_30 <= io_in_r_bypass_18_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_2_data_30 <= io_in_r_bypass_18_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_2_load_store_30 <= io_in_r_bypass_18_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_2_df_is_ws_30 <= io_in_r_bypass_18_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_2_stall_30 <= io_in_r_bypass_18_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_3_data_30 <= io_in_r_bypass_18_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_3_load_store_30 <= io_in_r_bypass_18_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_3_df_is_ws_30 <= io_in_r_bypass_18_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_18_3_stall_30 <= io_in_r_bypass_18_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_0_data_30 <= io_in_r_bypass_19_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_0_load_store_30 <= io_in_r_bypass_19_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_0_df_is_ws_30 <= io_in_r_bypass_19_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_0_stall_30 <= io_in_r_bypass_19_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_1_data_30 <= io_in_r_bypass_19_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_1_load_store_30 <= io_in_r_bypass_19_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_1_df_is_ws_30 <= io_in_r_bypass_19_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_1_stall_30 <= io_in_r_bypass_19_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_2_data_30 <= io_in_r_bypass_19_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_2_load_store_30 <= io_in_r_bypass_19_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_2_df_is_ws_30 <= io_in_r_bypass_19_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_2_stall_30 <= io_in_r_bypass_19_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_3_data_30 <= io_in_r_bypass_19_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_3_load_store_30 <= io_in_r_bypass_19_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_3_df_is_ws_30 <= io_in_r_bypass_19_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_19_3_stall_30 <= io_in_r_bypass_19_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_0_data_30 <= io_in_r_bypass_20_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_0_load_store_30 <= io_in_r_bypass_20_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_0_df_is_ws_30 <= io_in_r_bypass_20_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_0_stall_30 <= io_in_r_bypass_20_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_1_data_30 <= io_in_r_bypass_20_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_1_load_store_30 <= io_in_r_bypass_20_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_1_df_is_ws_30 <= io_in_r_bypass_20_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_1_stall_30 <= io_in_r_bypass_20_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_2_data_30 <= io_in_r_bypass_20_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_2_load_store_30 <= io_in_r_bypass_20_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_2_df_is_ws_30 <= io_in_r_bypass_20_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_2_stall_30 <= io_in_r_bypass_20_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_3_data_30 <= io_in_r_bypass_20_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_3_load_store_30 <= io_in_r_bypass_20_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_3_df_is_ws_30 <= io_in_r_bypass_20_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_20_3_stall_30 <= io_in_r_bypass_20_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_0_data_30 <= io_in_r_bypass_21_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_0_load_store_30 <= io_in_r_bypass_21_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_0_df_is_ws_30 <= io_in_r_bypass_21_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_0_stall_30 <= io_in_r_bypass_21_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_1_data_30 <= io_in_r_bypass_21_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_1_load_store_30 <= io_in_r_bypass_21_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_1_df_is_ws_30 <= io_in_r_bypass_21_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_1_stall_30 <= io_in_r_bypass_21_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_2_data_30 <= io_in_r_bypass_21_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_2_load_store_30 <= io_in_r_bypass_21_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_2_df_is_ws_30 <= io_in_r_bypass_21_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_2_stall_30 <= io_in_r_bypass_21_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_3_data_30 <= io_in_r_bypass_21_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_3_load_store_30 <= io_in_r_bypass_21_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_3_df_is_ws_30 <= io_in_r_bypass_21_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_21_3_stall_30 <= io_in_r_bypass_21_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_0_data_30 <= io_in_r_bypass_22_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_0_load_store_30 <= io_in_r_bypass_22_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_0_df_is_ws_30 <= io_in_r_bypass_22_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_0_stall_30 <= io_in_r_bypass_22_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_1_data_30 <= io_in_r_bypass_22_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_1_load_store_30 <= io_in_r_bypass_22_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_1_df_is_ws_30 <= io_in_r_bypass_22_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_1_stall_30 <= io_in_r_bypass_22_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_2_data_30 <= io_in_r_bypass_22_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_2_load_store_30 <= io_in_r_bypass_22_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_2_df_is_ws_30 <= io_in_r_bypass_22_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_2_stall_30 <= io_in_r_bypass_22_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_3_data_30 <= io_in_r_bypass_22_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_3_load_store_30 <= io_in_r_bypass_22_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_3_df_is_ws_30 <= io_in_r_bypass_22_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_22_3_stall_30 <= io_in_r_bypass_22_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_0_data_30 <= io_in_r_bypass_23_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_0_load_store_30 <= io_in_r_bypass_23_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_0_df_is_ws_30 <= io_in_r_bypass_23_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_0_stall_30 <= io_in_r_bypass_23_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_1_data_30 <= io_in_r_bypass_23_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_1_load_store_30 <= io_in_r_bypass_23_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_1_df_is_ws_30 <= io_in_r_bypass_23_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_1_stall_30 <= io_in_r_bypass_23_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_2_data_30 <= io_in_r_bypass_23_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_2_load_store_30 <= io_in_r_bypass_23_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_2_df_is_ws_30 <= io_in_r_bypass_23_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_2_stall_30 <= io_in_r_bypass_23_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_3_data_30 <= io_in_r_bypass_23_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_3_load_store_30 <= io_in_r_bypass_23_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_3_df_is_ws_30 <= io_in_r_bypass_23_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_23_3_stall_30 <= io_in_r_bypass_23_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_0_data_30 <= io_in_r_bypass_24_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_0_load_store_30 <= io_in_r_bypass_24_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_0_df_is_ws_30 <= io_in_r_bypass_24_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_0_stall_30 <= io_in_r_bypass_24_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_1_data_30 <= io_in_r_bypass_24_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_1_load_store_30 <= io_in_r_bypass_24_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_1_df_is_ws_30 <= io_in_r_bypass_24_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_1_stall_30 <= io_in_r_bypass_24_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_2_data_30 <= io_in_r_bypass_24_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_2_load_store_30 <= io_in_r_bypass_24_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_2_df_is_ws_30 <= io_in_r_bypass_24_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_2_stall_30 <= io_in_r_bypass_24_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_3_data_30 <= io_in_r_bypass_24_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_3_load_store_30 <= io_in_r_bypass_24_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_3_df_is_ws_30 <= io_in_r_bypass_24_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_24_3_stall_30 <= io_in_r_bypass_24_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_0_data_30 <= io_in_r_bypass_25_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_0_load_store_30 <= io_in_r_bypass_25_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_0_df_is_ws_30 <= io_in_r_bypass_25_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_0_stall_30 <= io_in_r_bypass_25_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_1_data_30 <= io_in_r_bypass_25_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_1_load_store_30 <= io_in_r_bypass_25_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_1_df_is_ws_30 <= io_in_r_bypass_25_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_1_stall_30 <= io_in_r_bypass_25_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_2_data_30 <= io_in_r_bypass_25_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_2_load_store_30 <= io_in_r_bypass_25_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_2_df_is_ws_30 <= io_in_r_bypass_25_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_2_stall_30 <= io_in_r_bypass_25_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_3_data_30 <= io_in_r_bypass_25_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_3_load_store_30 <= io_in_r_bypass_25_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_3_df_is_ws_30 <= io_in_r_bypass_25_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_25_3_stall_30 <= io_in_r_bypass_25_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_0_data_30 <= io_in_r_bypass_26_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_0_load_store_30 <= io_in_r_bypass_26_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_0_df_is_ws_30 <= io_in_r_bypass_26_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_0_stall_30 <= io_in_r_bypass_26_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_1_data_30 <= io_in_r_bypass_26_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_1_load_store_30 <= io_in_r_bypass_26_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_1_df_is_ws_30 <= io_in_r_bypass_26_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_1_stall_30 <= io_in_r_bypass_26_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_2_data_30 <= io_in_r_bypass_26_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_2_load_store_30 <= io_in_r_bypass_26_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_2_df_is_ws_30 <= io_in_r_bypass_26_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_2_stall_30 <= io_in_r_bypass_26_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_3_data_30 <= io_in_r_bypass_26_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_3_load_store_30 <= io_in_r_bypass_26_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_3_df_is_ws_30 <= io_in_r_bypass_26_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_26_3_stall_30 <= io_in_r_bypass_26_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_0_data_30 <= io_in_r_bypass_27_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_0_load_store_30 <= io_in_r_bypass_27_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_0_df_is_ws_30 <= io_in_r_bypass_27_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_0_stall_30 <= io_in_r_bypass_27_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_1_data_30 <= io_in_r_bypass_27_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_1_load_store_30 <= io_in_r_bypass_27_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_1_df_is_ws_30 <= io_in_r_bypass_27_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_1_stall_30 <= io_in_r_bypass_27_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_2_data_30 <= io_in_r_bypass_27_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_2_load_store_30 <= io_in_r_bypass_27_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_2_df_is_ws_30 <= io_in_r_bypass_27_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_2_stall_30 <= io_in_r_bypass_27_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_3_data_30 <= io_in_r_bypass_27_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_3_load_store_30 <= io_in_r_bypass_27_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_3_df_is_ws_30 <= io_in_r_bypass_27_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_27_3_stall_30 <= io_in_r_bypass_27_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_0_data_30 <= io_in_r_bypass_28_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_0_load_store_30 <= io_in_r_bypass_28_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_0_df_is_ws_30 <= io_in_r_bypass_28_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_0_stall_30 <= io_in_r_bypass_28_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_1_data_30 <= io_in_r_bypass_28_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_1_load_store_30 <= io_in_r_bypass_28_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_1_df_is_ws_30 <= io_in_r_bypass_28_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_1_stall_30 <= io_in_r_bypass_28_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_2_data_30 <= io_in_r_bypass_28_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_2_load_store_30 <= io_in_r_bypass_28_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_2_df_is_ws_30 <= io_in_r_bypass_28_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_2_stall_30 <= io_in_r_bypass_28_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_3_data_30 <= io_in_r_bypass_28_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_3_load_store_30 <= io_in_r_bypass_28_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_3_df_is_ws_30 <= io_in_r_bypass_28_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_28_3_stall_30 <= io_in_r_bypass_28_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_0_data_30 <= io_in_r_bypass_29_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_0_load_store_30 <= io_in_r_bypass_29_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_0_df_is_ws_30 <= io_in_r_bypass_29_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_0_stall_30 <= io_in_r_bypass_29_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_1_data_30 <= io_in_r_bypass_29_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_1_load_store_30 <= io_in_r_bypass_29_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_1_df_is_ws_30 <= io_in_r_bypass_29_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_1_stall_30 <= io_in_r_bypass_29_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_2_data_30 <= io_in_r_bypass_29_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_2_load_store_30 <= io_in_r_bypass_29_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_2_df_is_ws_30 <= io_in_r_bypass_29_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_2_stall_30 <= io_in_r_bypass_29_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_3_data_30 <= io_in_r_bypass_29_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_3_load_store_30 <= io_in_r_bypass_29_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_3_df_is_ws_30 <= io_in_r_bypass_29_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_29_3_stall_30 <= io_in_r_bypass_29_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_0_data_30 <= io_in_r_bypass_30_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_0_load_store_30 <= io_in_r_bypass_30_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_0_df_is_ws_30 <= io_in_r_bypass_30_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_0_stall_30 <= io_in_r_bypass_30_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_1_data_30 <= io_in_r_bypass_30_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_1_load_store_30 <= io_in_r_bypass_30_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_1_df_is_ws_30 <= io_in_r_bypass_30_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_1_stall_30 <= io_in_r_bypass_30_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_2_data_30 <= io_in_r_bypass_30_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_2_load_store_30 <= io_in_r_bypass_30_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_2_df_is_ws_30 <= io_in_r_bypass_30_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_2_stall_30 <= io_in_r_bypass_30_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_3_data_30 <= io_in_r_bypass_30_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_3_load_store_30 <= io_in_r_bypass_30_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_3_df_is_ws_30 <= io_in_r_bypass_30_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_30_3_stall_30 <= io_in_r_bypass_30_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_0_data_30 <= io_in_r_bypass_31_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_0_load_store_30 <= io_in_r_bypass_31_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_0_df_is_ws_30 <= io_in_r_bypass_31_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_0_stall_30 <= io_in_r_bypass_31_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_1_data_30 <= io_in_r_bypass_31_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_1_load_store_30 <= io_in_r_bypass_31_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_1_df_is_ws_30 <= io_in_r_bypass_31_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_1_stall_30 <= io_in_r_bypass_31_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_2_data_30 <= io_in_r_bypass_31_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_2_load_store_30 <= io_in_r_bypass_31_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_2_df_is_ws_30 <= io_in_r_bypass_31_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_2_stall_30 <= io_in_r_bypass_31_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_3_data_30 <= io_in_r_bypass_31_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_3_load_store_30 <= io_in_r_bypass_31_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_3_df_is_ws_30 <= io_in_r_bypass_31_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_31_3_stall_30 <= io_in_r_bypass_31_3_stall; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_0_data <= io_in_c_bypass_0_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_0_is_stationary <= io_in_c_bypass_0_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_1_data <= io_in_c_bypass_0_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_1_is_stationary <= io_in_c_bypass_0_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_2_data <= io_in_c_bypass_0_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_2_is_stationary <= io_in_c_bypass_0_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_3_data <= io_in_c_bypass_0_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_3_is_stationary <= io_in_c_bypass_0_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_0_data <= io_in_c_bypass_1_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_0_is_stationary <= io_in_c_bypass_1_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_1_data <= io_in_c_bypass_1_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_1_is_stationary <= io_in_c_bypass_1_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_2_data <= io_in_c_bypass_1_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_2_is_stationary <= io_in_c_bypass_1_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_3_data <= io_in_c_bypass_1_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_3_is_stationary <= io_in_c_bypass_1_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_0_data <= io_in_c_bypass_2_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_0_is_stationary <= io_in_c_bypass_2_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_1_data <= io_in_c_bypass_2_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_1_is_stationary <= io_in_c_bypass_2_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_2_data <= io_in_c_bypass_2_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_2_is_stationary <= io_in_c_bypass_2_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_3_data <= io_in_c_bypass_2_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_3_is_stationary <= io_in_c_bypass_2_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_0_data <= io_in_c_bypass_3_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_0_is_stationary <= io_in_c_bypass_3_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_1_data <= io_in_c_bypass_3_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_1_is_stationary <= io_in_c_bypass_3_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_2_data <= io_in_c_bypass_3_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_2_is_stationary <= io_in_c_bypass_3_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_3_data <= io_in_c_bypass_3_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_3_is_stationary <= io_in_c_bypass_3_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_0_data <= io_in_c_bypass_4_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_0_is_stationary <= io_in_c_bypass_4_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_1_data <= io_in_c_bypass_4_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_1_is_stationary <= io_in_c_bypass_4_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_2_data <= io_in_c_bypass_4_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_2_is_stationary <= io_in_c_bypass_4_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_3_data <= io_in_c_bypass_4_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_3_is_stationary <= io_in_c_bypass_4_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_0_data <= io_in_c_bypass_5_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_0_is_stationary <= io_in_c_bypass_5_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_1_data <= io_in_c_bypass_5_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_1_is_stationary <= io_in_c_bypass_5_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_2_data <= io_in_c_bypass_5_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_2_is_stationary <= io_in_c_bypass_5_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_3_data <= io_in_c_bypass_5_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_3_is_stationary <= io_in_c_bypass_5_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_0_data <= io_in_c_bypass_6_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_0_is_stationary <= io_in_c_bypass_6_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_1_data <= io_in_c_bypass_6_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_1_is_stationary <= io_in_c_bypass_6_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_2_data <= io_in_c_bypass_6_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_2_is_stationary <= io_in_c_bypass_6_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_3_data <= io_in_c_bypass_6_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_3_is_stationary <= io_in_c_bypass_6_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_0_data <= io_in_c_bypass_7_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_0_is_stationary <= io_in_c_bypass_7_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_1_data <= io_in_c_bypass_7_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_1_is_stationary <= io_in_c_bypass_7_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_2_data <= io_in_c_bypass_7_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_2_is_stationary <= io_in_c_bypass_7_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_3_data <= io_in_c_bypass_7_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_3_is_stationary <= io_in_c_bypass_7_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_0_data <= io_in_c_bypass_8_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_0_is_stationary <= io_in_c_bypass_8_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_1_data <= io_in_c_bypass_8_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_1_is_stationary <= io_in_c_bypass_8_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_2_data <= io_in_c_bypass_8_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_2_is_stationary <= io_in_c_bypass_8_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_3_data <= io_in_c_bypass_8_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_3_is_stationary <= io_in_c_bypass_8_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_0_data <= io_in_c_bypass_9_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_0_is_stationary <= io_in_c_bypass_9_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_1_data <= io_in_c_bypass_9_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_1_is_stationary <= io_in_c_bypass_9_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_2_data <= io_in_c_bypass_9_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_2_is_stationary <= io_in_c_bypass_9_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_3_data <= io_in_c_bypass_9_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_3_is_stationary <= io_in_c_bypass_9_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_0_data <= io_in_c_bypass_10_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_0_is_stationary <= io_in_c_bypass_10_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_1_data <= io_in_c_bypass_10_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_1_is_stationary <= io_in_c_bypass_10_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_2_data <= io_in_c_bypass_10_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_2_is_stationary <= io_in_c_bypass_10_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_3_data <= io_in_c_bypass_10_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_3_is_stationary <= io_in_c_bypass_10_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_0_data <= io_in_c_bypass_11_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_0_is_stationary <= io_in_c_bypass_11_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_1_data <= io_in_c_bypass_11_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_1_is_stationary <= io_in_c_bypass_11_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_2_data <= io_in_c_bypass_11_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_2_is_stationary <= io_in_c_bypass_11_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_3_data <= io_in_c_bypass_11_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_3_is_stationary <= io_in_c_bypass_11_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_0_data <= io_in_c_bypass_12_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_0_is_stationary <= io_in_c_bypass_12_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_1_data <= io_in_c_bypass_12_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_1_is_stationary <= io_in_c_bypass_12_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_2_data <= io_in_c_bypass_12_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_2_is_stationary <= io_in_c_bypass_12_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_3_data <= io_in_c_bypass_12_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_3_is_stationary <= io_in_c_bypass_12_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_0_data <= io_in_c_bypass_13_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_0_is_stationary <= io_in_c_bypass_13_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_1_data <= io_in_c_bypass_13_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_1_is_stationary <= io_in_c_bypass_13_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_2_data <= io_in_c_bypass_13_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_2_is_stationary <= io_in_c_bypass_13_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_3_data <= io_in_c_bypass_13_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_3_is_stationary <= io_in_c_bypass_13_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_0_data <= io_in_c_bypass_14_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_0_is_stationary <= io_in_c_bypass_14_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_1_data <= io_in_c_bypass_14_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_1_is_stationary <= io_in_c_bypass_14_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_2_data <= io_in_c_bypass_14_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_2_is_stationary <= io_in_c_bypass_14_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_3_data <= io_in_c_bypass_14_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_3_is_stationary <= io_in_c_bypass_14_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_0_data <= io_in_c_bypass_15_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_0_is_stationary <= io_in_c_bypass_15_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_1_data <= io_in_c_bypass_15_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_1_is_stationary <= io_in_c_bypass_15_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_2_data <= io_in_c_bypass_15_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_2_is_stationary <= io_in_c_bypass_15_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_3_data <= io_in_c_bypass_15_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_3_is_stationary <= io_in_c_bypass_15_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_0_data <= io_in_c_bypass_16_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_0_is_stationary <= io_in_c_bypass_16_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_1_data <= io_in_c_bypass_16_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_1_is_stationary <= io_in_c_bypass_16_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_2_data <= io_in_c_bypass_16_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_2_is_stationary <= io_in_c_bypass_16_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_3_data <= io_in_c_bypass_16_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_3_is_stationary <= io_in_c_bypass_16_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_0_data <= io_in_c_bypass_17_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_0_is_stationary <= io_in_c_bypass_17_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_1_data <= io_in_c_bypass_17_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_1_is_stationary <= io_in_c_bypass_17_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_2_data <= io_in_c_bypass_17_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_2_is_stationary <= io_in_c_bypass_17_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_3_data <= io_in_c_bypass_17_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_3_is_stationary <= io_in_c_bypass_17_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_0_data <= io_in_c_bypass_18_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_0_is_stationary <= io_in_c_bypass_18_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_1_data <= io_in_c_bypass_18_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_1_is_stationary <= io_in_c_bypass_18_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_2_data <= io_in_c_bypass_18_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_2_is_stationary <= io_in_c_bypass_18_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_3_data <= io_in_c_bypass_18_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_3_is_stationary <= io_in_c_bypass_18_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_0_data <= io_in_c_bypass_19_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_0_is_stationary <= io_in_c_bypass_19_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_1_data <= io_in_c_bypass_19_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_1_is_stationary <= io_in_c_bypass_19_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_2_data <= io_in_c_bypass_19_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_2_is_stationary <= io_in_c_bypass_19_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_3_data <= io_in_c_bypass_19_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_3_is_stationary <= io_in_c_bypass_19_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_0_data <= io_in_c_bypass_20_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_0_is_stationary <= io_in_c_bypass_20_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_1_data <= io_in_c_bypass_20_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_1_is_stationary <= io_in_c_bypass_20_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_2_data <= io_in_c_bypass_20_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_2_is_stationary <= io_in_c_bypass_20_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_3_data <= io_in_c_bypass_20_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_3_is_stationary <= io_in_c_bypass_20_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_0_data <= io_in_c_bypass_21_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_0_is_stationary <= io_in_c_bypass_21_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_1_data <= io_in_c_bypass_21_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_1_is_stationary <= io_in_c_bypass_21_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_2_data <= io_in_c_bypass_21_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_2_is_stationary <= io_in_c_bypass_21_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_3_data <= io_in_c_bypass_21_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_3_is_stationary <= io_in_c_bypass_21_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_0_data <= io_in_c_bypass_22_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_0_is_stationary <= io_in_c_bypass_22_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_1_data <= io_in_c_bypass_22_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_1_is_stationary <= io_in_c_bypass_22_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_2_data <= io_in_c_bypass_22_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_2_is_stationary <= io_in_c_bypass_22_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_3_data <= io_in_c_bypass_22_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_3_is_stationary <= io_in_c_bypass_22_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_0_data <= io_in_c_bypass_23_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_0_is_stationary <= io_in_c_bypass_23_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_1_data <= io_in_c_bypass_23_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_1_is_stationary <= io_in_c_bypass_23_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_2_data <= io_in_c_bypass_23_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_2_is_stationary <= io_in_c_bypass_23_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_3_data <= io_in_c_bypass_23_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_3_is_stationary <= io_in_c_bypass_23_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_0_data <= io_in_c_bypass_24_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_0_is_stationary <= io_in_c_bypass_24_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_1_data <= io_in_c_bypass_24_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_1_is_stationary <= io_in_c_bypass_24_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_2_data <= io_in_c_bypass_24_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_2_is_stationary <= io_in_c_bypass_24_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_3_data <= io_in_c_bypass_24_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_3_is_stationary <= io_in_c_bypass_24_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_0_data <= io_in_c_bypass_25_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_0_is_stationary <= io_in_c_bypass_25_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_1_data <= io_in_c_bypass_25_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_1_is_stationary <= io_in_c_bypass_25_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_2_data <= io_in_c_bypass_25_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_2_is_stationary <= io_in_c_bypass_25_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_3_data <= io_in_c_bypass_25_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_3_is_stationary <= io_in_c_bypass_25_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_0_data <= io_in_c_bypass_26_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_0_is_stationary <= io_in_c_bypass_26_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_1_data <= io_in_c_bypass_26_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_1_is_stationary <= io_in_c_bypass_26_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_2_data <= io_in_c_bypass_26_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_2_is_stationary <= io_in_c_bypass_26_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_3_data <= io_in_c_bypass_26_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_3_is_stationary <= io_in_c_bypass_26_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_0_data <= io_in_c_bypass_27_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_0_is_stationary <= io_in_c_bypass_27_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_1_data <= io_in_c_bypass_27_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_1_is_stationary <= io_in_c_bypass_27_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_2_data <= io_in_c_bypass_27_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_2_is_stationary <= io_in_c_bypass_27_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_3_data <= io_in_c_bypass_27_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_3_is_stationary <= io_in_c_bypass_27_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_0_data <= io_in_c_bypass_28_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_0_is_stationary <= io_in_c_bypass_28_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_1_data <= io_in_c_bypass_28_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_1_is_stationary <= io_in_c_bypass_28_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_2_data <= io_in_c_bypass_28_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_2_is_stationary <= io_in_c_bypass_28_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_3_data <= io_in_c_bypass_28_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_3_is_stationary <= io_in_c_bypass_28_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_0_data <= io_in_c_bypass_29_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_0_is_stationary <= io_in_c_bypass_29_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_1_data <= io_in_c_bypass_29_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_1_is_stationary <= io_in_c_bypass_29_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_2_data <= io_in_c_bypass_29_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_2_is_stationary <= io_in_c_bypass_29_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_3_data <= io_in_c_bypass_29_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_3_is_stationary <= io_in_c_bypass_29_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_0_data <= io_in_c_bypass_30_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_0_is_stationary <= io_in_c_bypass_30_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_1_data <= io_in_c_bypass_30_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_1_is_stationary <= io_in_c_bypass_30_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_2_data <= io_in_c_bypass_30_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_2_is_stationary <= io_in_c_bypass_30_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_3_data <= io_in_c_bypass_30_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_3_is_stationary <= io_in_c_bypass_30_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_0_data <= io_in_c_bypass_31_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_0_is_stationary <= io_in_c_bypass_31_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_1_data <= io_in_c_bypass_31_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_1_is_stationary <= io_in_c_bypass_31_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_2_data <= io_in_c_bypass_31_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_2_is_stationary <= io_in_c_bypass_31_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_3_data <= io_in_c_bypass_31_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_3_is_stationary <= io_in_c_bypass_31_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_0_data_1 <= io_in_c_bypass_0_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_0_is_stationary_1 <= io_in_c_bypass_0_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_1_data_1 <= io_in_c_bypass_0_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_1_is_stationary_1 <= io_in_c_bypass_0_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_2_data_1 <= io_in_c_bypass_0_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_2_is_stationary_1 <= io_in_c_bypass_0_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_3_data_1 <= io_in_c_bypass_0_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_3_is_stationary_1 <= io_in_c_bypass_0_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_0_data_1 <= io_in_c_bypass_1_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_0_is_stationary_1 <= io_in_c_bypass_1_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_1_data_1 <= io_in_c_bypass_1_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_1_is_stationary_1 <= io_in_c_bypass_1_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_2_data_1 <= io_in_c_bypass_1_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_2_is_stationary_1 <= io_in_c_bypass_1_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_3_data_1 <= io_in_c_bypass_1_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_3_is_stationary_1 <= io_in_c_bypass_1_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_0_data_1 <= io_in_c_bypass_2_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_0_is_stationary_1 <= io_in_c_bypass_2_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_1_data_1 <= io_in_c_bypass_2_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_1_is_stationary_1 <= io_in_c_bypass_2_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_2_data_1 <= io_in_c_bypass_2_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_2_is_stationary_1 <= io_in_c_bypass_2_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_3_data_1 <= io_in_c_bypass_2_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_3_is_stationary_1 <= io_in_c_bypass_2_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_0_data_1 <= io_in_c_bypass_3_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_0_is_stationary_1 <= io_in_c_bypass_3_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_1_data_1 <= io_in_c_bypass_3_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_1_is_stationary_1 <= io_in_c_bypass_3_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_2_data_1 <= io_in_c_bypass_3_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_2_is_stationary_1 <= io_in_c_bypass_3_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_3_data_1 <= io_in_c_bypass_3_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_3_is_stationary_1 <= io_in_c_bypass_3_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_0_data_1 <= io_in_c_bypass_4_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_0_is_stationary_1 <= io_in_c_bypass_4_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_1_data_1 <= io_in_c_bypass_4_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_1_is_stationary_1 <= io_in_c_bypass_4_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_2_data_1 <= io_in_c_bypass_4_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_2_is_stationary_1 <= io_in_c_bypass_4_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_3_data_1 <= io_in_c_bypass_4_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_3_is_stationary_1 <= io_in_c_bypass_4_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_0_data_1 <= io_in_c_bypass_5_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_0_is_stationary_1 <= io_in_c_bypass_5_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_1_data_1 <= io_in_c_bypass_5_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_1_is_stationary_1 <= io_in_c_bypass_5_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_2_data_1 <= io_in_c_bypass_5_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_2_is_stationary_1 <= io_in_c_bypass_5_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_3_data_1 <= io_in_c_bypass_5_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_3_is_stationary_1 <= io_in_c_bypass_5_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_0_data_1 <= io_in_c_bypass_6_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_0_is_stationary_1 <= io_in_c_bypass_6_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_1_data_1 <= io_in_c_bypass_6_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_1_is_stationary_1 <= io_in_c_bypass_6_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_2_data_1 <= io_in_c_bypass_6_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_2_is_stationary_1 <= io_in_c_bypass_6_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_3_data_1 <= io_in_c_bypass_6_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_3_is_stationary_1 <= io_in_c_bypass_6_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_0_data_1 <= io_in_c_bypass_7_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_0_is_stationary_1 <= io_in_c_bypass_7_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_1_data_1 <= io_in_c_bypass_7_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_1_is_stationary_1 <= io_in_c_bypass_7_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_2_data_1 <= io_in_c_bypass_7_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_2_is_stationary_1 <= io_in_c_bypass_7_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_3_data_1 <= io_in_c_bypass_7_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_3_is_stationary_1 <= io_in_c_bypass_7_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_0_data_1 <= io_in_c_bypass_8_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_0_is_stationary_1 <= io_in_c_bypass_8_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_1_data_1 <= io_in_c_bypass_8_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_1_is_stationary_1 <= io_in_c_bypass_8_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_2_data_1 <= io_in_c_bypass_8_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_2_is_stationary_1 <= io_in_c_bypass_8_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_3_data_1 <= io_in_c_bypass_8_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_3_is_stationary_1 <= io_in_c_bypass_8_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_0_data_1 <= io_in_c_bypass_9_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_0_is_stationary_1 <= io_in_c_bypass_9_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_1_data_1 <= io_in_c_bypass_9_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_1_is_stationary_1 <= io_in_c_bypass_9_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_2_data_1 <= io_in_c_bypass_9_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_2_is_stationary_1 <= io_in_c_bypass_9_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_3_data_1 <= io_in_c_bypass_9_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_3_is_stationary_1 <= io_in_c_bypass_9_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_0_data_1 <= io_in_c_bypass_10_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_0_is_stationary_1 <= io_in_c_bypass_10_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_1_data_1 <= io_in_c_bypass_10_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_1_is_stationary_1 <= io_in_c_bypass_10_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_2_data_1 <= io_in_c_bypass_10_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_2_is_stationary_1 <= io_in_c_bypass_10_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_3_data_1 <= io_in_c_bypass_10_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_3_is_stationary_1 <= io_in_c_bypass_10_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_0_data_1 <= io_in_c_bypass_11_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_0_is_stationary_1 <= io_in_c_bypass_11_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_1_data_1 <= io_in_c_bypass_11_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_1_is_stationary_1 <= io_in_c_bypass_11_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_2_data_1 <= io_in_c_bypass_11_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_2_is_stationary_1 <= io_in_c_bypass_11_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_3_data_1 <= io_in_c_bypass_11_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_3_is_stationary_1 <= io_in_c_bypass_11_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_0_data_1 <= io_in_c_bypass_12_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_0_is_stationary_1 <= io_in_c_bypass_12_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_1_data_1 <= io_in_c_bypass_12_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_1_is_stationary_1 <= io_in_c_bypass_12_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_2_data_1 <= io_in_c_bypass_12_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_2_is_stationary_1 <= io_in_c_bypass_12_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_3_data_1 <= io_in_c_bypass_12_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_3_is_stationary_1 <= io_in_c_bypass_12_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_0_data_1 <= io_in_c_bypass_13_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_0_is_stationary_1 <= io_in_c_bypass_13_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_1_data_1 <= io_in_c_bypass_13_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_1_is_stationary_1 <= io_in_c_bypass_13_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_2_data_1 <= io_in_c_bypass_13_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_2_is_stationary_1 <= io_in_c_bypass_13_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_3_data_1 <= io_in_c_bypass_13_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_3_is_stationary_1 <= io_in_c_bypass_13_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_0_data_1 <= io_in_c_bypass_14_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_0_is_stationary_1 <= io_in_c_bypass_14_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_1_data_1 <= io_in_c_bypass_14_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_1_is_stationary_1 <= io_in_c_bypass_14_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_2_data_1 <= io_in_c_bypass_14_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_2_is_stationary_1 <= io_in_c_bypass_14_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_3_data_1 <= io_in_c_bypass_14_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_3_is_stationary_1 <= io_in_c_bypass_14_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_0_data_1 <= io_in_c_bypass_15_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_0_is_stationary_1 <= io_in_c_bypass_15_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_1_data_1 <= io_in_c_bypass_15_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_1_is_stationary_1 <= io_in_c_bypass_15_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_2_data_1 <= io_in_c_bypass_15_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_2_is_stationary_1 <= io_in_c_bypass_15_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_3_data_1 <= io_in_c_bypass_15_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_3_is_stationary_1 <= io_in_c_bypass_15_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_0_data_1 <= io_in_c_bypass_16_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_0_is_stationary_1 <= io_in_c_bypass_16_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_1_data_1 <= io_in_c_bypass_16_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_1_is_stationary_1 <= io_in_c_bypass_16_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_2_data_1 <= io_in_c_bypass_16_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_2_is_stationary_1 <= io_in_c_bypass_16_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_3_data_1 <= io_in_c_bypass_16_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_3_is_stationary_1 <= io_in_c_bypass_16_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_0_data_1 <= io_in_c_bypass_17_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_0_is_stationary_1 <= io_in_c_bypass_17_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_1_data_1 <= io_in_c_bypass_17_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_1_is_stationary_1 <= io_in_c_bypass_17_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_2_data_1 <= io_in_c_bypass_17_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_2_is_stationary_1 <= io_in_c_bypass_17_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_3_data_1 <= io_in_c_bypass_17_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_3_is_stationary_1 <= io_in_c_bypass_17_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_0_data_1 <= io_in_c_bypass_18_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_0_is_stationary_1 <= io_in_c_bypass_18_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_1_data_1 <= io_in_c_bypass_18_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_1_is_stationary_1 <= io_in_c_bypass_18_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_2_data_1 <= io_in_c_bypass_18_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_2_is_stationary_1 <= io_in_c_bypass_18_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_3_data_1 <= io_in_c_bypass_18_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_3_is_stationary_1 <= io_in_c_bypass_18_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_0_data_1 <= io_in_c_bypass_19_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_0_is_stationary_1 <= io_in_c_bypass_19_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_1_data_1 <= io_in_c_bypass_19_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_1_is_stationary_1 <= io_in_c_bypass_19_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_2_data_1 <= io_in_c_bypass_19_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_2_is_stationary_1 <= io_in_c_bypass_19_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_3_data_1 <= io_in_c_bypass_19_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_3_is_stationary_1 <= io_in_c_bypass_19_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_0_data_1 <= io_in_c_bypass_20_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_0_is_stationary_1 <= io_in_c_bypass_20_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_1_data_1 <= io_in_c_bypass_20_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_1_is_stationary_1 <= io_in_c_bypass_20_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_2_data_1 <= io_in_c_bypass_20_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_2_is_stationary_1 <= io_in_c_bypass_20_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_3_data_1 <= io_in_c_bypass_20_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_3_is_stationary_1 <= io_in_c_bypass_20_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_0_data_1 <= io_in_c_bypass_21_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_0_is_stationary_1 <= io_in_c_bypass_21_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_1_data_1 <= io_in_c_bypass_21_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_1_is_stationary_1 <= io_in_c_bypass_21_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_2_data_1 <= io_in_c_bypass_21_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_2_is_stationary_1 <= io_in_c_bypass_21_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_3_data_1 <= io_in_c_bypass_21_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_3_is_stationary_1 <= io_in_c_bypass_21_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_0_data_1 <= io_in_c_bypass_22_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_0_is_stationary_1 <= io_in_c_bypass_22_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_1_data_1 <= io_in_c_bypass_22_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_1_is_stationary_1 <= io_in_c_bypass_22_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_2_data_1 <= io_in_c_bypass_22_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_2_is_stationary_1 <= io_in_c_bypass_22_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_3_data_1 <= io_in_c_bypass_22_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_3_is_stationary_1 <= io_in_c_bypass_22_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_0_data_1 <= io_in_c_bypass_23_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_0_is_stationary_1 <= io_in_c_bypass_23_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_1_data_1 <= io_in_c_bypass_23_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_1_is_stationary_1 <= io_in_c_bypass_23_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_2_data_1 <= io_in_c_bypass_23_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_2_is_stationary_1 <= io_in_c_bypass_23_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_3_data_1 <= io_in_c_bypass_23_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_3_is_stationary_1 <= io_in_c_bypass_23_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_0_data_1 <= io_in_c_bypass_24_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_0_is_stationary_1 <= io_in_c_bypass_24_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_1_data_1 <= io_in_c_bypass_24_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_1_is_stationary_1 <= io_in_c_bypass_24_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_2_data_1 <= io_in_c_bypass_24_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_2_is_stationary_1 <= io_in_c_bypass_24_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_3_data_1 <= io_in_c_bypass_24_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_3_is_stationary_1 <= io_in_c_bypass_24_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_0_data_1 <= io_in_c_bypass_25_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_0_is_stationary_1 <= io_in_c_bypass_25_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_1_data_1 <= io_in_c_bypass_25_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_1_is_stationary_1 <= io_in_c_bypass_25_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_2_data_1 <= io_in_c_bypass_25_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_2_is_stationary_1 <= io_in_c_bypass_25_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_3_data_1 <= io_in_c_bypass_25_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_3_is_stationary_1 <= io_in_c_bypass_25_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_0_data_1 <= io_in_c_bypass_26_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_0_is_stationary_1 <= io_in_c_bypass_26_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_1_data_1 <= io_in_c_bypass_26_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_1_is_stationary_1 <= io_in_c_bypass_26_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_2_data_1 <= io_in_c_bypass_26_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_2_is_stationary_1 <= io_in_c_bypass_26_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_3_data_1 <= io_in_c_bypass_26_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_3_is_stationary_1 <= io_in_c_bypass_26_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_0_data_1 <= io_in_c_bypass_27_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_0_is_stationary_1 <= io_in_c_bypass_27_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_1_data_1 <= io_in_c_bypass_27_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_1_is_stationary_1 <= io_in_c_bypass_27_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_2_data_1 <= io_in_c_bypass_27_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_2_is_stationary_1 <= io_in_c_bypass_27_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_3_data_1 <= io_in_c_bypass_27_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_3_is_stationary_1 <= io_in_c_bypass_27_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_0_data_1 <= io_in_c_bypass_28_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_0_is_stationary_1 <= io_in_c_bypass_28_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_1_data_1 <= io_in_c_bypass_28_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_1_is_stationary_1 <= io_in_c_bypass_28_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_2_data_1 <= io_in_c_bypass_28_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_2_is_stationary_1 <= io_in_c_bypass_28_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_3_data_1 <= io_in_c_bypass_28_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_3_is_stationary_1 <= io_in_c_bypass_28_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_0_data_1 <= io_in_c_bypass_29_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_0_is_stationary_1 <= io_in_c_bypass_29_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_1_data_1 <= io_in_c_bypass_29_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_1_is_stationary_1 <= io_in_c_bypass_29_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_2_data_1 <= io_in_c_bypass_29_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_2_is_stationary_1 <= io_in_c_bypass_29_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_3_data_1 <= io_in_c_bypass_29_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_3_is_stationary_1 <= io_in_c_bypass_29_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_0_data_1 <= io_in_c_bypass_30_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_0_is_stationary_1 <= io_in_c_bypass_30_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_1_data_1 <= io_in_c_bypass_30_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_1_is_stationary_1 <= io_in_c_bypass_30_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_2_data_1 <= io_in_c_bypass_30_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_2_is_stationary_1 <= io_in_c_bypass_30_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_3_data_1 <= io_in_c_bypass_30_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_3_is_stationary_1 <= io_in_c_bypass_30_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_0_data_1 <= io_in_c_bypass_31_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_0_is_stationary_1 <= io_in_c_bypass_31_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_1_data_1 <= io_in_c_bypass_31_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_1_is_stationary_1 <= io_in_c_bypass_31_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_2_data_1 <= io_in_c_bypass_31_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_2_is_stationary_1 <= io_in_c_bypass_31_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_3_data_1 <= io_in_c_bypass_31_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_3_is_stationary_1 <= io_in_c_bypass_31_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_0_data_2 <= io_in_c_bypass_0_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_0_is_stationary_2 <= io_in_c_bypass_0_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_1_data_2 <= io_in_c_bypass_0_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_1_is_stationary_2 <= io_in_c_bypass_0_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_2_data_2 <= io_in_c_bypass_0_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_2_is_stationary_2 <= io_in_c_bypass_0_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_3_data_2 <= io_in_c_bypass_0_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_3_is_stationary_2 <= io_in_c_bypass_0_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_0_data_2 <= io_in_c_bypass_1_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_0_is_stationary_2 <= io_in_c_bypass_1_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_1_data_2 <= io_in_c_bypass_1_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_1_is_stationary_2 <= io_in_c_bypass_1_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_2_data_2 <= io_in_c_bypass_1_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_2_is_stationary_2 <= io_in_c_bypass_1_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_3_data_2 <= io_in_c_bypass_1_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_3_is_stationary_2 <= io_in_c_bypass_1_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_0_data_2 <= io_in_c_bypass_2_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_0_is_stationary_2 <= io_in_c_bypass_2_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_1_data_2 <= io_in_c_bypass_2_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_1_is_stationary_2 <= io_in_c_bypass_2_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_2_data_2 <= io_in_c_bypass_2_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_2_is_stationary_2 <= io_in_c_bypass_2_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_3_data_2 <= io_in_c_bypass_2_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_3_is_stationary_2 <= io_in_c_bypass_2_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_0_data_2 <= io_in_c_bypass_3_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_0_is_stationary_2 <= io_in_c_bypass_3_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_1_data_2 <= io_in_c_bypass_3_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_1_is_stationary_2 <= io_in_c_bypass_3_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_2_data_2 <= io_in_c_bypass_3_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_2_is_stationary_2 <= io_in_c_bypass_3_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_3_data_2 <= io_in_c_bypass_3_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_3_is_stationary_2 <= io_in_c_bypass_3_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_0_data_2 <= io_in_c_bypass_4_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_0_is_stationary_2 <= io_in_c_bypass_4_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_1_data_2 <= io_in_c_bypass_4_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_1_is_stationary_2 <= io_in_c_bypass_4_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_2_data_2 <= io_in_c_bypass_4_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_2_is_stationary_2 <= io_in_c_bypass_4_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_3_data_2 <= io_in_c_bypass_4_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_3_is_stationary_2 <= io_in_c_bypass_4_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_0_data_2 <= io_in_c_bypass_5_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_0_is_stationary_2 <= io_in_c_bypass_5_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_1_data_2 <= io_in_c_bypass_5_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_1_is_stationary_2 <= io_in_c_bypass_5_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_2_data_2 <= io_in_c_bypass_5_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_2_is_stationary_2 <= io_in_c_bypass_5_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_3_data_2 <= io_in_c_bypass_5_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_3_is_stationary_2 <= io_in_c_bypass_5_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_0_data_2 <= io_in_c_bypass_6_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_0_is_stationary_2 <= io_in_c_bypass_6_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_1_data_2 <= io_in_c_bypass_6_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_1_is_stationary_2 <= io_in_c_bypass_6_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_2_data_2 <= io_in_c_bypass_6_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_2_is_stationary_2 <= io_in_c_bypass_6_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_3_data_2 <= io_in_c_bypass_6_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_3_is_stationary_2 <= io_in_c_bypass_6_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_0_data_2 <= io_in_c_bypass_7_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_0_is_stationary_2 <= io_in_c_bypass_7_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_1_data_2 <= io_in_c_bypass_7_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_1_is_stationary_2 <= io_in_c_bypass_7_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_2_data_2 <= io_in_c_bypass_7_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_2_is_stationary_2 <= io_in_c_bypass_7_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_3_data_2 <= io_in_c_bypass_7_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_3_is_stationary_2 <= io_in_c_bypass_7_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_0_data_2 <= io_in_c_bypass_8_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_0_is_stationary_2 <= io_in_c_bypass_8_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_1_data_2 <= io_in_c_bypass_8_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_1_is_stationary_2 <= io_in_c_bypass_8_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_2_data_2 <= io_in_c_bypass_8_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_2_is_stationary_2 <= io_in_c_bypass_8_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_3_data_2 <= io_in_c_bypass_8_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_3_is_stationary_2 <= io_in_c_bypass_8_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_0_data_2 <= io_in_c_bypass_9_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_0_is_stationary_2 <= io_in_c_bypass_9_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_1_data_2 <= io_in_c_bypass_9_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_1_is_stationary_2 <= io_in_c_bypass_9_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_2_data_2 <= io_in_c_bypass_9_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_2_is_stationary_2 <= io_in_c_bypass_9_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_3_data_2 <= io_in_c_bypass_9_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_3_is_stationary_2 <= io_in_c_bypass_9_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_0_data_2 <= io_in_c_bypass_10_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_0_is_stationary_2 <= io_in_c_bypass_10_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_1_data_2 <= io_in_c_bypass_10_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_1_is_stationary_2 <= io_in_c_bypass_10_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_2_data_2 <= io_in_c_bypass_10_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_2_is_stationary_2 <= io_in_c_bypass_10_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_3_data_2 <= io_in_c_bypass_10_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_3_is_stationary_2 <= io_in_c_bypass_10_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_0_data_2 <= io_in_c_bypass_11_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_0_is_stationary_2 <= io_in_c_bypass_11_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_1_data_2 <= io_in_c_bypass_11_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_1_is_stationary_2 <= io_in_c_bypass_11_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_2_data_2 <= io_in_c_bypass_11_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_2_is_stationary_2 <= io_in_c_bypass_11_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_3_data_2 <= io_in_c_bypass_11_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_3_is_stationary_2 <= io_in_c_bypass_11_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_0_data_2 <= io_in_c_bypass_12_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_0_is_stationary_2 <= io_in_c_bypass_12_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_1_data_2 <= io_in_c_bypass_12_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_1_is_stationary_2 <= io_in_c_bypass_12_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_2_data_2 <= io_in_c_bypass_12_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_2_is_stationary_2 <= io_in_c_bypass_12_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_3_data_2 <= io_in_c_bypass_12_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_3_is_stationary_2 <= io_in_c_bypass_12_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_0_data_2 <= io_in_c_bypass_13_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_0_is_stationary_2 <= io_in_c_bypass_13_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_1_data_2 <= io_in_c_bypass_13_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_1_is_stationary_2 <= io_in_c_bypass_13_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_2_data_2 <= io_in_c_bypass_13_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_2_is_stationary_2 <= io_in_c_bypass_13_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_3_data_2 <= io_in_c_bypass_13_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_3_is_stationary_2 <= io_in_c_bypass_13_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_0_data_2 <= io_in_c_bypass_14_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_0_is_stationary_2 <= io_in_c_bypass_14_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_1_data_2 <= io_in_c_bypass_14_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_1_is_stationary_2 <= io_in_c_bypass_14_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_2_data_2 <= io_in_c_bypass_14_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_2_is_stationary_2 <= io_in_c_bypass_14_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_3_data_2 <= io_in_c_bypass_14_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_3_is_stationary_2 <= io_in_c_bypass_14_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_0_data_2 <= io_in_c_bypass_15_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_0_is_stationary_2 <= io_in_c_bypass_15_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_1_data_2 <= io_in_c_bypass_15_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_1_is_stationary_2 <= io_in_c_bypass_15_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_2_data_2 <= io_in_c_bypass_15_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_2_is_stationary_2 <= io_in_c_bypass_15_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_3_data_2 <= io_in_c_bypass_15_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_3_is_stationary_2 <= io_in_c_bypass_15_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_0_data_2 <= io_in_c_bypass_16_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_0_is_stationary_2 <= io_in_c_bypass_16_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_1_data_2 <= io_in_c_bypass_16_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_1_is_stationary_2 <= io_in_c_bypass_16_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_2_data_2 <= io_in_c_bypass_16_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_2_is_stationary_2 <= io_in_c_bypass_16_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_3_data_2 <= io_in_c_bypass_16_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_3_is_stationary_2 <= io_in_c_bypass_16_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_0_data_2 <= io_in_c_bypass_17_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_0_is_stationary_2 <= io_in_c_bypass_17_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_1_data_2 <= io_in_c_bypass_17_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_1_is_stationary_2 <= io_in_c_bypass_17_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_2_data_2 <= io_in_c_bypass_17_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_2_is_stationary_2 <= io_in_c_bypass_17_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_3_data_2 <= io_in_c_bypass_17_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_3_is_stationary_2 <= io_in_c_bypass_17_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_0_data_2 <= io_in_c_bypass_18_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_0_is_stationary_2 <= io_in_c_bypass_18_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_1_data_2 <= io_in_c_bypass_18_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_1_is_stationary_2 <= io_in_c_bypass_18_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_2_data_2 <= io_in_c_bypass_18_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_2_is_stationary_2 <= io_in_c_bypass_18_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_3_data_2 <= io_in_c_bypass_18_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_3_is_stationary_2 <= io_in_c_bypass_18_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_0_data_2 <= io_in_c_bypass_19_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_0_is_stationary_2 <= io_in_c_bypass_19_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_1_data_2 <= io_in_c_bypass_19_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_1_is_stationary_2 <= io_in_c_bypass_19_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_2_data_2 <= io_in_c_bypass_19_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_2_is_stationary_2 <= io_in_c_bypass_19_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_3_data_2 <= io_in_c_bypass_19_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_3_is_stationary_2 <= io_in_c_bypass_19_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_0_data_2 <= io_in_c_bypass_20_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_0_is_stationary_2 <= io_in_c_bypass_20_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_1_data_2 <= io_in_c_bypass_20_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_1_is_stationary_2 <= io_in_c_bypass_20_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_2_data_2 <= io_in_c_bypass_20_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_2_is_stationary_2 <= io_in_c_bypass_20_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_3_data_2 <= io_in_c_bypass_20_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_3_is_stationary_2 <= io_in_c_bypass_20_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_0_data_2 <= io_in_c_bypass_21_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_0_is_stationary_2 <= io_in_c_bypass_21_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_1_data_2 <= io_in_c_bypass_21_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_1_is_stationary_2 <= io_in_c_bypass_21_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_2_data_2 <= io_in_c_bypass_21_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_2_is_stationary_2 <= io_in_c_bypass_21_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_3_data_2 <= io_in_c_bypass_21_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_3_is_stationary_2 <= io_in_c_bypass_21_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_0_data_2 <= io_in_c_bypass_22_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_0_is_stationary_2 <= io_in_c_bypass_22_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_1_data_2 <= io_in_c_bypass_22_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_1_is_stationary_2 <= io_in_c_bypass_22_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_2_data_2 <= io_in_c_bypass_22_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_2_is_stationary_2 <= io_in_c_bypass_22_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_3_data_2 <= io_in_c_bypass_22_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_3_is_stationary_2 <= io_in_c_bypass_22_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_0_data_2 <= io_in_c_bypass_23_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_0_is_stationary_2 <= io_in_c_bypass_23_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_1_data_2 <= io_in_c_bypass_23_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_1_is_stationary_2 <= io_in_c_bypass_23_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_2_data_2 <= io_in_c_bypass_23_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_2_is_stationary_2 <= io_in_c_bypass_23_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_3_data_2 <= io_in_c_bypass_23_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_3_is_stationary_2 <= io_in_c_bypass_23_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_0_data_2 <= io_in_c_bypass_24_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_0_is_stationary_2 <= io_in_c_bypass_24_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_1_data_2 <= io_in_c_bypass_24_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_1_is_stationary_2 <= io_in_c_bypass_24_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_2_data_2 <= io_in_c_bypass_24_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_2_is_stationary_2 <= io_in_c_bypass_24_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_3_data_2 <= io_in_c_bypass_24_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_3_is_stationary_2 <= io_in_c_bypass_24_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_0_data_2 <= io_in_c_bypass_25_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_0_is_stationary_2 <= io_in_c_bypass_25_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_1_data_2 <= io_in_c_bypass_25_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_1_is_stationary_2 <= io_in_c_bypass_25_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_2_data_2 <= io_in_c_bypass_25_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_2_is_stationary_2 <= io_in_c_bypass_25_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_3_data_2 <= io_in_c_bypass_25_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_3_is_stationary_2 <= io_in_c_bypass_25_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_0_data_2 <= io_in_c_bypass_26_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_0_is_stationary_2 <= io_in_c_bypass_26_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_1_data_2 <= io_in_c_bypass_26_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_1_is_stationary_2 <= io_in_c_bypass_26_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_2_data_2 <= io_in_c_bypass_26_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_2_is_stationary_2 <= io_in_c_bypass_26_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_3_data_2 <= io_in_c_bypass_26_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_3_is_stationary_2 <= io_in_c_bypass_26_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_0_data_2 <= io_in_c_bypass_27_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_0_is_stationary_2 <= io_in_c_bypass_27_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_1_data_2 <= io_in_c_bypass_27_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_1_is_stationary_2 <= io_in_c_bypass_27_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_2_data_2 <= io_in_c_bypass_27_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_2_is_stationary_2 <= io_in_c_bypass_27_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_3_data_2 <= io_in_c_bypass_27_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_3_is_stationary_2 <= io_in_c_bypass_27_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_0_data_2 <= io_in_c_bypass_28_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_0_is_stationary_2 <= io_in_c_bypass_28_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_1_data_2 <= io_in_c_bypass_28_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_1_is_stationary_2 <= io_in_c_bypass_28_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_2_data_2 <= io_in_c_bypass_28_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_2_is_stationary_2 <= io_in_c_bypass_28_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_3_data_2 <= io_in_c_bypass_28_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_3_is_stationary_2 <= io_in_c_bypass_28_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_0_data_2 <= io_in_c_bypass_29_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_0_is_stationary_2 <= io_in_c_bypass_29_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_1_data_2 <= io_in_c_bypass_29_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_1_is_stationary_2 <= io_in_c_bypass_29_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_2_data_2 <= io_in_c_bypass_29_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_2_is_stationary_2 <= io_in_c_bypass_29_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_3_data_2 <= io_in_c_bypass_29_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_3_is_stationary_2 <= io_in_c_bypass_29_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_0_data_2 <= io_in_c_bypass_30_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_0_is_stationary_2 <= io_in_c_bypass_30_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_1_data_2 <= io_in_c_bypass_30_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_1_is_stationary_2 <= io_in_c_bypass_30_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_2_data_2 <= io_in_c_bypass_30_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_2_is_stationary_2 <= io_in_c_bypass_30_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_3_data_2 <= io_in_c_bypass_30_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_3_is_stationary_2 <= io_in_c_bypass_30_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_0_data_2 <= io_in_c_bypass_31_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_0_is_stationary_2 <= io_in_c_bypass_31_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_1_data_2 <= io_in_c_bypass_31_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_1_is_stationary_2 <= io_in_c_bypass_31_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_2_data_2 <= io_in_c_bypass_31_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_2_is_stationary_2 <= io_in_c_bypass_31_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_3_data_2 <= io_in_c_bypass_31_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_3_is_stationary_2 <= io_in_c_bypass_31_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_0_data_3 <= io_in_c_bypass_0_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_0_is_stationary_3 <= io_in_c_bypass_0_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_1_data_3 <= io_in_c_bypass_0_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_1_is_stationary_3 <= io_in_c_bypass_0_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_2_data_3 <= io_in_c_bypass_0_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_2_is_stationary_3 <= io_in_c_bypass_0_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_3_data_3 <= io_in_c_bypass_0_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_3_is_stationary_3 <= io_in_c_bypass_0_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_0_data_3 <= io_in_c_bypass_1_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_0_is_stationary_3 <= io_in_c_bypass_1_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_1_data_3 <= io_in_c_bypass_1_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_1_is_stationary_3 <= io_in_c_bypass_1_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_2_data_3 <= io_in_c_bypass_1_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_2_is_stationary_3 <= io_in_c_bypass_1_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_3_data_3 <= io_in_c_bypass_1_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_3_is_stationary_3 <= io_in_c_bypass_1_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_0_data_3 <= io_in_c_bypass_2_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_0_is_stationary_3 <= io_in_c_bypass_2_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_1_data_3 <= io_in_c_bypass_2_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_1_is_stationary_3 <= io_in_c_bypass_2_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_2_data_3 <= io_in_c_bypass_2_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_2_is_stationary_3 <= io_in_c_bypass_2_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_3_data_3 <= io_in_c_bypass_2_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_3_is_stationary_3 <= io_in_c_bypass_2_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_0_data_3 <= io_in_c_bypass_3_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_0_is_stationary_3 <= io_in_c_bypass_3_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_1_data_3 <= io_in_c_bypass_3_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_1_is_stationary_3 <= io_in_c_bypass_3_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_2_data_3 <= io_in_c_bypass_3_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_2_is_stationary_3 <= io_in_c_bypass_3_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_3_data_3 <= io_in_c_bypass_3_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_3_is_stationary_3 <= io_in_c_bypass_3_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_0_data_3 <= io_in_c_bypass_4_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_0_is_stationary_3 <= io_in_c_bypass_4_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_1_data_3 <= io_in_c_bypass_4_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_1_is_stationary_3 <= io_in_c_bypass_4_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_2_data_3 <= io_in_c_bypass_4_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_2_is_stationary_3 <= io_in_c_bypass_4_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_3_data_3 <= io_in_c_bypass_4_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_3_is_stationary_3 <= io_in_c_bypass_4_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_0_data_3 <= io_in_c_bypass_5_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_0_is_stationary_3 <= io_in_c_bypass_5_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_1_data_3 <= io_in_c_bypass_5_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_1_is_stationary_3 <= io_in_c_bypass_5_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_2_data_3 <= io_in_c_bypass_5_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_2_is_stationary_3 <= io_in_c_bypass_5_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_3_data_3 <= io_in_c_bypass_5_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_3_is_stationary_3 <= io_in_c_bypass_5_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_0_data_3 <= io_in_c_bypass_6_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_0_is_stationary_3 <= io_in_c_bypass_6_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_1_data_3 <= io_in_c_bypass_6_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_1_is_stationary_3 <= io_in_c_bypass_6_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_2_data_3 <= io_in_c_bypass_6_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_2_is_stationary_3 <= io_in_c_bypass_6_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_3_data_3 <= io_in_c_bypass_6_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_3_is_stationary_3 <= io_in_c_bypass_6_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_0_data_3 <= io_in_c_bypass_7_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_0_is_stationary_3 <= io_in_c_bypass_7_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_1_data_3 <= io_in_c_bypass_7_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_1_is_stationary_3 <= io_in_c_bypass_7_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_2_data_3 <= io_in_c_bypass_7_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_2_is_stationary_3 <= io_in_c_bypass_7_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_3_data_3 <= io_in_c_bypass_7_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_3_is_stationary_3 <= io_in_c_bypass_7_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_0_data_3 <= io_in_c_bypass_8_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_0_is_stationary_3 <= io_in_c_bypass_8_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_1_data_3 <= io_in_c_bypass_8_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_1_is_stationary_3 <= io_in_c_bypass_8_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_2_data_3 <= io_in_c_bypass_8_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_2_is_stationary_3 <= io_in_c_bypass_8_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_3_data_3 <= io_in_c_bypass_8_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_3_is_stationary_3 <= io_in_c_bypass_8_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_0_data_3 <= io_in_c_bypass_9_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_0_is_stationary_3 <= io_in_c_bypass_9_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_1_data_3 <= io_in_c_bypass_9_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_1_is_stationary_3 <= io_in_c_bypass_9_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_2_data_3 <= io_in_c_bypass_9_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_2_is_stationary_3 <= io_in_c_bypass_9_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_3_data_3 <= io_in_c_bypass_9_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_3_is_stationary_3 <= io_in_c_bypass_9_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_0_data_3 <= io_in_c_bypass_10_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_0_is_stationary_3 <= io_in_c_bypass_10_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_1_data_3 <= io_in_c_bypass_10_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_1_is_stationary_3 <= io_in_c_bypass_10_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_2_data_3 <= io_in_c_bypass_10_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_2_is_stationary_3 <= io_in_c_bypass_10_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_3_data_3 <= io_in_c_bypass_10_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_3_is_stationary_3 <= io_in_c_bypass_10_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_0_data_3 <= io_in_c_bypass_11_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_0_is_stationary_3 <= io_in_c_bypass_11_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_1_data_3 <= io_in_c_bypass_11_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_1_is_stationary_3 <= io_in_c_bypass_11_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_2_data_3 <= io_in_c_bypass_11_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_2_is_stationary_3 <= io_in_c_bypass_11_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_3_data_3 <= io_in_c_bypass_11_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_3_is_stationary_3 <= io_in_c_bypass_11_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_0_data_3 <= io_in_c_bypass_12_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_0_is_stationary_3 <= io_in_c_bypass_12_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_1_data_3 <= io_in_c_bypass_12_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_1_is_stationary_3 <= io_in_c_bypass_12_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_2_data_3 <= io_in_c_bypass_12_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_2_is_stationary_3 <= io_in_c_bypass_12_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_3_data_3 <= io_in_c_bypass_12_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_3_is_stationary_3 <= io_in_c_bypass_12_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_0_data_3 <= io_in_c_bypass_13_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_0_is_stationary_3 <= io_in_c_bypass_13_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_1_data_3 <= io_in_c_bypass_13_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_1_is_stationary_3 <= io_in_c_bypass_13_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_2_data_3 <= io_in_c_bypass_13_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_2_is_stationary_3 <= io_in_c_bypass_13_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_3_data_3 <= io_in_c_bypass_13_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_3_is_stationary_3 <= io_in_c_bypass_13_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_0_data_3 <= io_in_c_bypass_14_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_0_is_stationary_3 <= io_in_c_bypass_14_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_1_data_3 <= io_in_c_bypass_14_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_1_is_stationary_3 <= io_in_c_bypass_14_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_2_data_3 <= io_in_c_bypass_14_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_2_is_stationary_3 <= io_in_c_bypass_14_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_3_data_3 <= io_in_c_bypass_14_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_3_is_stationary_3 <= io_in_c_bypass_14_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_0_data_3 <= io_in_c_bypass_15_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_0_is_stationary_3 <= io_in_c_bypass_15_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_1_data_3 <= io_in_c_bypass_15_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_1_is_stationary_3 <= io_in_c_bypass_15_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_2_data_3 <= io_in_c_bypass_15_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_2_is_stationary_3 <= io_in_c_bypass_15_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_3_data_3 <= io_in_c_bypass_15_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_3_is_stationary_3 <= io_in_c_bypass_15_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_0_data_3 <= io_in_c_bypass_16_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_0_is_stationary_3 <= io_in_c_bypass_16_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_1_data_3 <= io_in_c_bypass_16_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_1_is_stationary_3 <= io_in_c_bypass_16_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_2_data_3 <= io_in_c_bypass_16_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_2_is_stationary_3 <= io_in_c_bypass_16_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_3_data_3 <= io_in_c_bypass_16_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_3_is_stationary_3 <= io_in_c_bypass_16_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_0_data_3 <= io_in_c_bypass_17_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_0_is_stationary_3 <= io_in_c_bypass_17_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_1_data_3 <= io_in_c_bypass_17_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_1_is_stationary_3 <= io_in_c_bypass_17_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_2_data_3 <= io_in_c_bypass_17_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_2_is_stationary_3 <= io_in_c_bypass_17_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_3_data_3 <= io_in_c_bypass_17_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_3_is_stationary_3 <= io_in_c_bypass_17_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_0_data_3 <= io_in_c_bypass_18_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_0_is_stationary_3 <= io_in_c_bypass_18_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_1_data_3 <= io_in_c_bypass_18_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_1_is_stationary_3 <= io_in_c_bypass_18_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_2_data_3 <= io_in_c_bypass_18_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_2_is_stationary_3 <= io_in_c_bypass_18_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_3_data_3 <= io_in_c_bypass_18_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_3_is_stationary_3 <= io_in_c_bypass_18_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_0_data_3 <= io_in_c_bypass_19_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_0_is_stationary_3 <= io_in_c_bypass_19_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_1_data_3 <= io_in_c_bypass_19_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_1_is_stationary_3 <= io_in_c_bypass_19_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_2_data_3 <= io_in_c_bypass_19_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_2_is_stationary_3 <= io_in_c_bypass_19_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_3_data_3 <= io_in_c_bypass_19_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_3_is_stationary_3 <= io_in_c_bypass_19_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_0_data_3 <= io_in_c_bypass_20_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_0_is_stationary_3 <= io_in_c_bypass_20_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_1_data_3 <= io_in_c_bypass_20_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_1_is_stationary_3 <= io_in_c_bypass_20_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_2_data_3 <= io_in_c_bypass_20_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_2_is_stationary_3 <= io_in_c_bypass_20_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_3_data_3 <= io_in_c_bypass_20_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_3_is_stationary_3 <= io_in_c_bypass_20_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_0_data_3 <= io_in_c_bypass_21_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_0_is_stationary_3 <= io_in_c_bypass_21_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_1_data_3 <= io_in_c_bypass_21_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_1_is_stationary_3 <= io_in_c_bypass_21_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_2_data_3 <= io_in_c_bypass_21_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_2_is_stationary_3 <= io_in_c_bypass_21_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_3_data_3 <= io_in_c_bypass_21_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_3_is_stationary_3 <= io_in_c_bypass_21_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_0_data_3 <= io_in_c_bypass_22_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_0_is_stationary_3 <= io_in_c_bypass_22_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_1_data_3 <= io_in_c_bypass_22_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_1_is_stationary_3 <= io_in_c_bypass_22_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_2_data_3 <= io_in_c_bypass_22_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_2_is_stationary_3 <= io_in_c_bypass_22_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_3_data_3 <= io_in_c_bypass_22_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_3_is_stationary_3 <= io_in_c_bypass_22_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_0_data_3 <= io_in_c_bypass_23_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_0_is_stationary_3 <= io_in_c_bypass_23_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_1_data_3 <= io_in_c_bypass_23_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_1_is_stationary_3 <= io_in_c_bypass_23_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_2_data_3 <= io_in_c_bypass_23_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_2_is_stationary_3 <= io_in_c_bypass_23_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_3_data_3 <= io_in_c_bypass_23_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_3_is_stationary_3 <= io_in_c_bypass_23_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_0_data_3 <= io_in_c_bypass_24_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_0_is_stationary_3 <= io_in_c_bypass_24_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_1_data_3 <= io_in_c_bypass_24_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_1_is_stationary_3 <= io_in_c_bypass_24_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_2_data_3 <= io_in_c_bypass_24_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_2_is_stationary_3 <= io_in_c_bypass_24_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_3_data_3 <= io_in_c_bypass_24_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_3_is_stationary_3 <= io_in_c_bypass_24_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_0_data_3 <= io_in_c_bypass_25_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_0_is_stationary_3 <= io_in_c_bypass_25_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_1_data_3 <= io_in_c_bypass_25_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_1_is_stationary_3 <= io_in_c_bypass_25_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_2_data_3 <= io_in_c_bypass_25_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_2_is_stationary_3 <= io_in_c_bypass_25_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_3_data_3 <= io_in_c_bypass_25_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_3_is_stationary_3 <= io_in_c_bypass_25_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_0_data_3 <= io_in_c_bypass_26_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_0_is_stationary_3 <= io_in_c_bypass_26_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_1_data_3 <= io_in_c_bypass_26_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_1_is_stationary_3 <= io_in_c_bypass_26_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_2_data_3 <= io_in_c_bypass_26_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_2_is_stationary_3 <= io_in_c_bypass_26_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_3_data_3 <= io_in_c_bypass_26_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_3_is_stationary_3 <= io_in_c_bypass_26_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_0_data_3 <= io_in_c_bypass_27_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_0_is_stationary_3 <= io_in_c_bypass_27_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_1_data_3 <= io_in_c_bypass_27_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_1_is_stationary_3 <= io_in_c_bypass_27_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_2_data_3 <= io_in_c_bypass_27_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_2_is_stationary_3 <= io_in_c_bypass_27_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_3_data_3 <= io_in_c_bypass_27_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_3_is_stationary_3 <= io_in_c_bypass_27_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_0_data_3 <= io_in_c_bypass_28_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_0_is_stationary_3 <= io_in_c_bypass_28_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_1_data_3 <= io_in_c_bypass_28_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_1_is_stationary_3 <= io_in_c_bypass_28_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_2_data_3 <= io_in_c_bypass_28_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_2_is_stationary_3 <= io_in_c_bypass_28_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_3_data_3 <= io_in_c_bypass_28_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_3_is_stationary_3 <= io_in_c_bypass_28_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_0_data_3 <= io_in_c_bypass_29_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_0_is_stationary_3 <= io_in_c_bypass_29_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_1_data_3 <= io_in_c_bypass_29_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_1_is_stationary_3 <= io_in_c_bypass_29_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_2_data_3 <= io_in_c_bypass_29_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_2_is_stationary_3 <= io_in_c_bypass_29_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_3_data_3 <= io_in_c_bypass_29_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_3_is_stationary_3 <= io_in_c_bypass_29_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_0_data_3 <= io_in_c_bypass_30_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_0_is_stationary_3 <= io_in_c_bypass_30_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_1_data_3 <= io_in_c_bypass_30_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_1_is_stationary_3 <= io_in_c_bypass_30_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_2_data_3 <= io_in_c_bypass_30_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_2_is_stationary_3 <= io_in_c_bypass_30_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_3_data_3 <= io_in_c_bypass_30_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_3_is_stationary_3 <= io_in_c_bypass_30_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_0_data_3 <= io_in_c_bypass_31_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_0_is_stationary_3 <= io_in_c_bypass_31_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_1_data_3 <= io_in_c_bypass_31_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_1_is_stationary_3 <= io_in_c_bypass_31_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_2_data_3 <= io_in_c_bypass_31_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_2_is_stationary_3 <= io_in_c_bypass_31_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_3_data_3 <= io_in_c_bypass_31_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_3_is_stationary_3 <= io_in_c_bypass_31_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_0_data_4 <= io_in_c_bypass_0_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_0_is_stationary_4 <= io_in_c_bypass_0_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_1_data_4 <= io_in_c_bypass_0_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_1_is_stationary_4 <= io_in_c_bypass_0_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_2_data_4 <= io_in_c_bypass_0_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_2_is_stationary_4 <= io_in_c_bypass_0_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_3_data_4 <= io_in_c_bypass_0_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_3_is_stationary_4 <= io_in_c_bypass_0_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_0_data_4 <= io_in_c_bypass_1_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_0_is_stationary_4 <= io_in_c_bypass_1_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_1_data_4 <= io_in_c_bypass_1_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_1_is_stationary_4 <= io_in_c_bypass_1_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_2_data_4 <= io_in_c_bypass_1_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_2_is_stationary_4 <= io_in_c_bypass_1_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_3_data_4 <= io_in_c_bypass_1_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_3_is_stationary_4 <= io_in_c_bypass_1_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_0_data_4 <= io_in_c_bypass_2_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_0_is_stationary_4 <= io_in_c_bypass_2_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_1_data_4 <= io_in_c_bypass_2_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_1_is_stationary_4 <= io_in_c_bypass_2_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_2_data_4 <= io_in_c_bypass_2_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_2_is_stationary_4 <= io_in_c_bypass_2_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_3_data_4 <= io_in_c_bypass_2_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_3_is_stationary_4 <= io_in_c_bypass_2_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_0_data_4 <= io_in_c_bypass_3_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_0_is_stationary_4 <= io_in_c_bypass_3_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_1_data_4 <= io_in_c_bypass_3_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_1_is_stationary_4 <= io_in_c_bypass_3_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_2_data_4 <= io_in_c_bypass_3_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_2_is_stationary_4 <= io_in_c_bypass_3_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_3_data_4 <= io_in_c_bypass_3_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_3_is_stationary_4 <= io_in_c_bypass_3_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_0_data_4 <= io_in_c_bypass_4_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_0_is_stationary_4 <= io_in_c_bypass_4_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_1_data_4 <= io_in_c_bypass_4_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_1_is_stationary_4 <= io_in_c_bypass_4_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_2_data_4 <= io_in_c_bypass_4_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_2_is_stationary_4 <= io_in_c_bypass_4_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_3_data_4 <= io_in_c_bypass_4_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_3_is_stationary_4 <= io_in_c_bypass_4_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_0_data_4 <= io_in_c_bypass_5_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_0_is_stationary_4 <= io_in_c_bypass_5_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_1_data_4 <= io_in_c_bypass_5_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_1_is_stationary_4 <= io_in_c_bypass_5_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_2_data_4 <= io_in_c_bypass_5_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_2_is_stationary_4 <= io_in_c_bypass_5_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_3_data_4 <= io_in_c_bypass_5_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_3_is_stationary_4 <= io_in_c_bypass_5_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_0_data_4 <= io_in_c_bypass_6_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_0_is_stationary_4 <= io_in_c_bypass_6_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_1_data_4 <= io_in_c_bypass_6_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_1_is_stationary_4 <= io_in_c_bypass_6_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_2_data_4 <= io_in_c_bypass_6_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_2_is_stationary_4 <= io_in_c_bypass_6_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_3_data_4 <= io_in_c_bypass_6_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_3_is_stationary_4 <= io_in_c_bypass_6_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_0_data_4 <= io_in_c_bypass_7_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_0_is_stationary_4 <= io_in_c_bypass_7_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_1_data_4 <= io_in_c_bypass_7_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_1_is_stationary_4 <= io_in_c_bypass_7_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_2_data_4 <= io_in_c_bypass_7_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_2_is_stationary_4 <= io_in_c_bypass_7_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_3_data_4 <= io_in_c_bypass_7_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_3_is_stationary_4 <= io_in_c_bypass_7_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_0_data_4 <= io_in_c_bypass_8_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_0_is_stationary_4 <= io_in_c_bypass_8_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_1_data_4 <= io_in_c_bypass_8_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_1_is_stationary_4 <= io_in_c_bypass_8_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_2_data_4 <= io_in_c_bypass_8_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_2_is_stationary_4 <= io_in_c_bypass_8_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_3_data_4 <= io_in_c_bypass_8_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_3_is_stationary_4 <= io_in_c_bypass_8_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_0_data_4 <= io_in_c_bypass_9_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_0_is_stationary_4 <= io_in_c_bypass_9_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_1_data_4 <= io_in_c_bypass_9_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_1_is_stationary_4 <= io_in_c_bypass_9_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_2_data_4 <= io_in_c_bypass_9_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_2_is_stationary_4 <= io_in_c_bypass_9_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_3_data_4 <= io_in_c_bypass_9_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_3_is_stationary_4 <= io_in_c_bypass_9_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_0_data_4 <= io_in_c_bypass_10_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_0_is_stationary_4 <= io_in_c_bypass_10_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_1_data_4 <= io_in_c_bypass_10_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_1_is_stationary_4 <= io_in_c_bypass_10_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_2_data_4 <= io_in_c_bypass_10_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_2_is_stationary_4 <= io_in_c_bypass_10_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_3_data_4 <= io_in_c_bypass_10_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_3_is_stationary_4 <= io_in_c_bypass_10_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_0_data_4 <= io_in_c_bypass_11_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_0_is_stationary_4 <= io_in_c_bypass_11_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_1_data_4 <= io_in_c_bypass_11_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_1_is_stationary_4 <= io_in_c_bypass_11_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_2_data_4 <= io_in_c_bypass_11_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_2_is_stationary_4 <= io_in_c_bypass_11_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_3_data_4 <= io_in_c_bypass_11_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_3_is_stationary_4 <= io_in_c_bypass_11_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_0_data_4 <= io_in_c_bypass_12_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_0_is_stationary_4 <= io_in_c_bypass_12_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_1_data_4 <= io_in_c_bypass_12_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_1_is_stationary_4 <= io_in_c_bypass_12_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_2_data_4 <= io_in_c_bypass_12_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_2_is_stationary_4 <= io_in_c_bypass_12_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_3_data_4 <= io_in_c_bypass_12_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_3_is_stationary_4 <= io_in_c_bypass_12_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_0_data_4 <= io_in_c_bypass_13_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_0_is_stationary_4 <= io_in_c_bypass_13_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_1_data_4 <= io_in_c_bypass_13_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_1_is_stationary_4 <= io_in_c_bypass_13_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_2_data_4 <= io_in_c_bypass_13_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_2_is_stationary_4 <= io_in_c_bypass_13_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_3_data_4 <= io_in_c_bypass_13_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_3_is_stationary_4 <= io_in_c_bypass_13_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_0_data_4 <= io_in_c_bypass_14_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_0_is_stationary_4 <= io_in_c_bypass_14_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_1_data_4 <= io_in_c_bypass_14_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_1_is_stationary_4 <= io_in_c_bypass_14_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_2_data_4 <= io_in_c_bypass_14_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_2_is_stationary_4 <= io_in_c_bypass_14_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_3_data_4 <= io_in_c_bypass_14_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_3_is_stationary_4 <= io_in_c_bypass_14_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_0_data_4 <= io_in_c_bypass_15_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_0_is_stationary_4 <= io_in_c_bypass_15_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_1_data_4 <= io_in_c_bypass_15_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_1_is_stationary_4 <= io_in_c_bypass_15_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_2_data_4 <= io_in_c_bypass_15_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_2_is_stationary_4 <= io_in_c_bypass_15_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_3_data_4 <= io_in_c_bypass_15_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_3_is_stationary_4 <= io_in_c_bypass_15_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_0_data_4 <= io_in_c_bypass_16_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_0_is_stationary_4 <= io_in_c_bypass_16_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_1_data_4 <= io_in_c_bypass_16_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_1_is_stationary_4 <= io_in_c_bypass_16_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_2_data_4 <= io_in_c_bypass_16_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_2_is_stationary_4 <= io_in_c_bypass_16_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_3_data_4 <= io_in_c_bypass_16_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_3_is_stationary_4 <= io_in_c_bypass_16_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_0_data_4 <= io_in_c_bypass_17_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_0_is_stationary_4 <= io_in_c_bypass_17_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_1_data_4 <= io_in_c_bypass_17_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_1_is_stationary_4 <= io_in_c_bypass_17_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_2_data_4 <= io_in_c_bypass_17_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_2_is_stationary_4 <= io_in_c_bypass_17_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_3_data_4 <= io_in_c_bypass_17_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_3_is_stationary_4 <= io_in_c_bypass_17_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_0_data_4 <= io_in_c_bypass_18_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_0_is_stationary_4 <= io_in_c_bypass_18_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_1_data_4 <= io_in_c_bypass_18_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_1_is_stationary_4 <= io_in_c_bypass_18_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_2_data_4 <= io_in_c_bypass_18_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_2_is_stationary_4 <= io_in_c_bypass_18_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_3_data_4 <= io_in_c_bypass_18_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_3_is_stationary_4 <= io_in_c_bypass_18_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_0_data_4 <= io_in_c_bypass_19_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_0_is_stationary_4 <= io_in_c_bypass_19_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_1_data_4 <= io_in_c_bypass_19_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_1_is_stationary_4 <= io_in_c_bypass_19_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_2_data_4 <= io_in_c_bypass_19_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_2_is_stationary_4 <= io_in_c_bypass_19_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_3_data_4 <= io_in_c_bypass_19_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_3_is_stationary_4 <= io_in_c_bypass_19_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_0_data_4 <= io_in_c_bypass_20_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_0_is_stationary_4 <= io_in_c_bypass_20_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_1_data_4 <= io_in_c_bypass_20_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_1_is_stationary_4 <= io_in_c_bypass_20_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_2_data_4 <= io_in_c_bypass_20_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_2_is_stationary_4 <= io_in_c_bypass_20_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_3_data_4 <= io_in_c_bypass_20_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_3_is_stationary_4 <= io_in_c_bypass_20_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_0_data_4 <= io_in_c_bypass_21_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_0_is_stationary_4 <= io_in_c_bypass_21_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_1_data_4 <= io_in_c_bypass_21_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_1_is_stationary_4 <= io_in_c_bypass_21_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_2_data_4 <= io_in_c_bypass_21_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_2_is_stationary_4 <= io_in_c_bypass_21_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_3_data_4 <= io_in_c_bypass_21_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_3_is_stationary_4 <= io_in_c_bypass_21_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_0_data_4 <= io_in_c_bypass_22_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_0_is_stationary_4 <= io_in_c_bypass_22_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_1_data_4 <= io_in_c_bypass_22_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_1_is_stationary_4 <= io_in_c_bypass_22_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_2_data_4 <= io_in_c_bypass_22_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_2_is_stationary_4 <= io_in_c_bypass_22_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_3_data_4 <= io_in_c_bypass_22_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_3_is_stationary_4 <= io_in_c_bypass_22_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_0_data_4 <= io_in_c_bypass_23_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_0_is_stationary_4 <= io_in_c_bypass_23_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_1_data_4 <= io_in_c_bypass_23_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_1_is_stationary_4 <= io_in_c_bypass_23_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_2_data_4 <= io_in_c_bypass_23_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_2_is_stationary_4 <= io_in_c_bypass_23_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_3_data_4 <= io_in_c_bypass_23_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_3_is_stationary_4 <= io_in_c_bypass_23_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_0_data_4 <= io_in_c_bypass_24_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_0_is_stationary_4 <= io_in_c_bypass_24_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_1_data_4 <= io_in_c_bypass_24_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_1_is_stationary_4 <= io_in_c_bypass_24_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_2_data_4 <= io_in_c_bypass_24_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_2_is_stationary_4 <= io_in_c_bypass_24_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_3_data_4 <= io_in_c_bypass_24_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_3_is_stationary_4 <= io_in_c_bypass_24_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_0_data_4 <= io_in_c_bypass_25_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_0_is_stationary_4 <= io_in_c_bypass_25_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_1_data_4 <= io_in_c_bypass_25_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_1_is_stationary_4 <= io_in_c_bypass_25_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_2_data_4 <= io_in_c_bypass_25_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_2_is_stationary_4 <= io_in_c_bypass_25_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_3_data_4 <= io_in_c_bypass_25_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_3_is_stationary_4 <= io_in_c_bypass_25_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_0_data_4 <= io_in_c_bypass_26_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_0_is_stationary_4 <= io_in_c_bypass_26_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_1_data_4 <= io_in_c_bypass_26_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_1_is_stationary_4 <= io_in_c_bypass_26_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_2_data_4 <= io_in_c_bypass_26_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_2_is_stationary_4 <= io_in_c_bypass_26_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_3_data_4 <= io_in_c_bypass_26_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_3_is_stationary_4 <= io_in_c_bypass_26_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_0_data_4 <= io_in_c_bypass_27_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_0_is_stationary_4 <= io_in_c_bypass_27_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_1_data_4 <= io_in_c_bypass_27_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_1_is_stationary_4 <= io_in_c_bypass_27_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_2_data_4 <= io_in_c_bypass_27_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_2_is_stationary_4 <= io_in_c_bypass_27_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_3_data_4 <= io_in_c_bypass_27_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_3_is_stationary_4 <= io_in_c_bypass_27_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_0_data_4 <= io_in_c_bypass_28_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_0_is_stationary_4 <= io_in_c_bypass_28_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_1_data_4 <= io_in_c_bypass_28_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_1_is_stationary_4 <= io_in_c_bypass_28_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_2_data_4 <= io_in_c_bypass_28_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_2_is_stationary_4 <= io_in_c_bypass_28_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_3_data_4 <= io_in_c_bypass_28_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_3_is_stationary_4 <= io_in_c_bypass_28_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_0_data_4 <= io_in_c_bypass_29_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_0_is_stationary_4 <= io_in_c_bypass_29_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_1_data_4 <= io_in_c_bypass_29_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_1_is_stationary_4 <= io_in_c_bypass_29_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_2_data_4 <= io_in_c_bypass_29_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_2_is_stationary_4 <= io_in_c_bypass_29_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_3_data_4 <= io_in_c_bypass_29_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_3_is_stationary_4 <= io_in_c_bypass_29_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_0_data_4 <= io_in_c_bypass_30_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_0_is_stationary_4 <= io_in_c_bypass_30_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_1_data_4 <= io_in_c_bypass_30_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_1_is_stationary_4 <= io_in_c_bypass_30_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_2_data_4 <= io_in_c_bypass_30_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_2_is_stationary_4 <= io_in_c_bypass_30_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_3_data_4 <= io_in_c_bypass_30_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_3_is_stationary_4 <= io_in_c_bypass_30_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_0_data_4 <= io_in_c_bypass_31_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_0_is_stationary_4 <= io_in_c_bypass_31_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_1_data_4 <= io_in_c_bypass_31_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_1_is_stationary_4 <= io_in_c_bypass_31_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_2_data_4 <= io_in_c_bypass_31_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_2_is_stationary_4 <= io_in_c_bypass_31_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_3_data_4 <= io_in_c_bypass_31_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_3_is_stationary_4 <= io_in_c_bypass_31_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_0_data_5 <= io_in_c_bypass_0_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_0_is_stationary_5 <= io_in_c_bypass_0_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_1_data_5 <= io_in_c_bypass_0_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_1_is_stationary_5 <= io_in_c_bypass_0_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_2_data_5 <= io_in_c_bypass_0_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_2_is_stationary_5 <= io_in_c_bypass_0_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_3_data_5 <= io_in_c_bypass_0_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_3_is_stationary_5 <= io_in_c_bypass_0_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_0_data_5 <= io_in_c_bypass_1_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_0_is_stationary_5 <= io_in_c_bypass_1_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_1_data_5 <= io_in_c_bypass_1_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_1_is_stationary_5 <= io_in_c_bypass_1_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_2_data_5 <= io_in_c_bypass_1_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_2_is_stationary_5 <= io_in_c_bypass_1_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_3_data_5 <= io_in_c_bypass_1_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_3_is_stationary_5 <= io_in_c_bypass_1_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_0_data_5 <= io_in_c_bypass_2_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_0_is_stationary_5 <= io_in_c_bypass_2_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_1_data_5 <= io_in_c_bypass_2_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_1_is_stationary_5 <= io_in_c_bypass_2_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_2_data_5 <= io_in_c_bypass_2_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_2_is_stationary_5 <= io_in_c_bypass_2_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_3_data_5 <= io_in_c_bypass_2_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_3_is_stationary_5 <= io_in_c_bypass_2_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_0_data_5 <= io_in_c_bypass_3_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_0_is_stationary_5 <= io_in_c_bypass_3_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_1_data_5 <= io_in_c_bypass_3_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_1_is_stationary_5 <= io_in_c_bypass_3_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_2_data_5 <= io_in_c_bypass_3_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_2_is_stationary_5 <= io_in_c_bypass_3_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_3_data_5 <= io_in_c_bypass_3_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_3_is_stationary_5 <= io_in_c_bypass_3_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_0_data_5 <= io_in_c_bypass_4_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_0_is_stationary_5 <= io_in_c_bypass_4_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_1_data_5 <= io_in_c_bypass_4_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_1_is_stationary_5 <= io_in_c_bypass_4_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_2_data_5 <= io_in_c_bypass_4_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_2_is_stationary_5 <= io_in_c_bypass_4_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_3_data_5 <= io_in_c_bypass_4_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_3_is_stationary_5 <= io_in_c_bypass_4_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_0_data_5 <= io_in_c_bypass_5_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_0_is_stationary_5 <= io_in_c_bypass_5_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_1_data_5 <= io_in_c_bypass_5_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_1_is_stationary_5 <= io_in_c_bypass_5_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_2_data_5 <= io_in_c_bypass_5_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_2_is_stationary_5 <= io_in_c_bypass_5_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_3_data_5 <= io_in_c_bypass_5_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_3_is_stationary_5 <= io_in_c_bypass_5_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_0_data_5 <= io_in_c_bypass_6_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_0_is_stationary_5 <= io_in_c_bypass_6_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_1_data_5 <= io_in_c_bypass_6_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_1_is_stationary_5 <= io_in_c_bypass_6_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_2_data_5 <= io_in_c_bypass_6_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_2_is_stationary_5 <= io_in_c_bypass_6_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_3_data_5 <= io_in_c_bypass_6_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_3_is_stationary_5 <= io_in_c_bypass_6_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_0_data_5 <= io_in_c_bypass_7_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_0_is_stationary_5 <= io_in_c_bypass_7_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_1_data_5 <= io_in_c_bypass_7_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_1_is_stationary_5 <= io_in_c_bypass_7_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_2_data_5 <= io_in_c_bypass_7_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_2_is_stationary_5 <= io_in_c_bypass_7_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_3_data_5 <= io_in_c_bypass_7_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_3_is_stationary_5 <= io_in_c_bypass_7_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_0_data_5 <= io_in_c_bypass_8_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_0_is_stationary_5 <= io_in_c_bypass_8_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_1_data_5 <= io_in_c_bypass_8_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_1_is_stationary_5 <= io_in_c_bypass_8_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_2_data_5 <= io_in_c_bypass_8_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_2_is_stationary_5 <= io_in_c_bypass_8_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_3_data_5 <= io_in_c_bypass_8_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_3_is_stationary_5 <= io_in_c_bypass_8_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_0_data_5 <= io_in_c_bypass_9_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_0_is_stationary_5 <= io_in_c_bypass_9_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_1_data_5 <= io_in_c_bypass_9_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_1_is_stationary_5 <= io_in_c_bypass_9_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_2_data_5 <= io_in_c_bypass_9_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_2_is_stationary_5 <= io_in_c_bypass_9_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_3_data_5 <= io_in_c_bypass_9_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_3_is_stationary_5 <= io_in_c_bypass_9_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_0_data_5 <= io_in_c_bypass_10_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_0_is_stationary_5 <= io_in_c_bypass_10_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_1_data_5 <= io_in_c_bypass_10_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_1_is_stationary_5 <= io_in_c_bypass_10_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_2_data_5 <= io_in_c_bypass_10_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_2_is_stationary_5 <= io_in_c_bypass_10_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_3_data_5 <= io_in_c_bypass_10_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_3_is_stationary_5 <= io_in_c_bypass_10_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_0_data_5 <= io_in_c_bypass_11_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_0_is_stationary_5 <= io_in_c_bypass_11_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_1_data_5 <= io_in_c_bypass_11_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_1_is_stationary_5 <= io_in_c_bypass_11_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_2_data_5 <= io_in_c_bypass_11_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_2_is_stationary_5 <= io_in_c_bypass_11_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_3_data_5 <= io_in_c_bypass_11_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_3_is_stationary_5 <= io_in_c_bypass_11_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_0_data_5 <= io_in_c_bypass_12_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_0_is_stationary_5 <= io_in_c_bypass_12_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_1_data_5 <= io_in_c_bypass_12_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_1_is_stationary_5 <= io_in_c_bypass_12_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_2_data_5 <= io_in_c_bypass_12_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_2_is_stationary_5 <= io_in_c_bypass_12_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_3_data_5 <= io_in_c_bypass_12_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_3_is_stationary_5 <= io_in_c_bypass_12_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_0_data_5 <= io_in_c_bypass_13_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_0_is_stationary_5 <= io_in_c_bypass_13_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_1_data_5 <= io_in_c_bypass_13_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_1_is_stationary_5 <= io_in_c_bypass_13_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_2_data_5 <= io_in_c_bypass_13_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_2_is_stationary_5 <= io_in_c_bypass_13_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_3_data_5 <= io_in_c_bypass_13_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_3_is_stationary_5 <= io_in_c_bypass_13_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_0_data_5 <= io_in_c_bypass_14_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_0_is_stationary_5 <= io_in_c_bypass_14_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_1_data_5 <= io_in_c_bypass_14_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_1_is_stationary_5 <= io_in_c_bypass_14_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_2_data_5 <= io_in_c_bypass_14_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_2_is_stationary_5 <= io_in_c_bypass_14_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_3_data_5 <= io_in_c_bypass_14_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_3_is_stationary_5 <= io_in_c_bypass_14_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_0_data_5 <= io_in_c_bypass_15_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_0_is_stationary_5 <= io_in_c_bypass_15_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_1_data_5 <= io_in_c_bypass_15_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_1_is_stationary_5 <= io_in_c_bypass_15_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_2_data_5 <= io_in_c_bypass_15_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_2_is_stationary_5 <= io_in_c_bypass_15_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_3_data_5 <= io_in_c_bypass_15_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_3_is_stationary_5 <= io_in_c_bypass_15_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_0_data_5 <= io_in_c_bypass_16_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_0_is_stationary_5 <= io_in_c_bypass_16_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_1_data_5 <= io_in_c_bypass_16_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_1_is_stationary_5 <= io_in_c_bypass_16_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_2_data_5 <= io_in_c_bypass_16_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_2_is_stationary_5 <= io_in_c_bypass_16_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_3_data_5 <= io_in_c_bypass_16_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_3_is_stationary_5 <= io_in_c_bypass_16_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_0_data_5 <= io_in_c_bypass_17_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_0_is_stationary_5 <= io_in_c_bypass_17_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_1_data_5 <= io_in_c_bypass_17_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_1_is_stationary_5 <= io_in_c_bypass_17_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_2_data_5 <= io_in_c_bypass_17_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_2_is_stationary_5 <= io_in_c_bypass_17_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_3_data_5 <= io_in_c_bypass_17_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_3_is_stationary_5 <= io_in_c_bypass_17_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_0_data_5 <= io_in_c_bypass_18_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_0_is_stationary_5 <= io_in_c_bypass_18_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_1_data_5 <= io_in_c_bypass_18_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_1_is_stationary_5 <= io_in_c_bypass_18_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_2_data_5 <= io_in_c_bypass_18_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_2_is_stationary_5 <= io_in_c_bypass_18_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_3_data_5 <= io_in_c_bypass_18_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_3_is_stationary_5 <= io_in_c_bypass_18_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_0_data_5 <= io_in_c_bypass_19_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_0_is_stationary_5 <= io_in_c_bypass_19_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_1_data_5 <= io_in_c_bypass_19_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_1_is_stationary_5 <= io_in_c_bypass_19_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_2_data_5 <= io_in_c_bypass_19_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_2_is_stationary_5 <= io_in_c_bypass_19_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_3_data_5 <= io_in_c_bypass_19_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_3_is_stationary_5 <= io_in_c_bypass_19_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_0_data_5 <= io_in_c_bypass_20_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_0_is_stationary_5 <= io_in_c_bypass_20_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_1_data_5 <= io_in_c_bypass_20_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_1_is_stationary_5 <= io_in_c_bypass_20_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_2_data_5 <= io_in_c_bypass_20_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_2_is_stationary_5 <= io_in_c_bypass_20_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_3_data_5 <= io_in_c_bypass_20_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_3_is_stationary_5 <= io_in_c_bypass_20_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_0_data_5 <= io_in_c_bypass_21_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_0_is_stationary_5 <= io_in_c_bypass_21_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_1_data_5 <= io_in_c_bypass_21_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_1_is_stationary_5 <= io_in_c_bypass_21_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_2_data_5 <= io_in_c_bypass_21_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_2_is_stationary_5 <= io_in_c_bypass_21_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_3_data_5 <= io_in_c_bypass_21_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_3_is_stationary_5 <= io_in_c_bypass_21_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_0_data_5 <= io_in_c_bypass_22_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_0_is_stationary_5 <= io_in_c_bypass_22_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_1_data_5 <= io_in_c_bypass_22_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_1_is_stationary_5 <= io_in_c_bypass_22_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_2_data_5 <= io_in_c_bypass_22_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_2_is_stationary_5 <= io_in_c_bypass_22_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_3_data_5 <= io_in_c_bypass_22_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_3_is_stationary_5 <= io_in_c_bypass_22_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_0_data_5 <= io_in_c_bypass_23_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_0_is_stationary_5 <= io_in_c_bypass_23_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_1_data_5 <= io_in_c_bypass_23_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_1_is_stationary_5 <= io_in_c_bypass_23_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_2_data_5 <= io_in_c_bypass_23_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_2_is_stationary_5 <= io_in_c_bypass_23_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_3_data_5 <= io_in_c_bypass_23_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_3_is_stationary_5 <= io_in_c_bypass_23_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_0_data_5 <= io_in_c_bypass_24_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_0_is_stationary_5 <= io_in_c_bypass_24_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_1_data_5 <= io_in_c_bypass_24_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_1_is_stationary_5 <= io_in_c_bypass_24_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_2_data_5 <= io_in_c_bypass_24_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_2_is_stationary_5 <= io_in_c_bypass_24_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_3_data_5 <= io_in_c_bypass_24_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_3_is_stationary_5 <= io_in_c_bypass_24_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_0_data_5 <= io_in_c_bypass_25_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_0_is_stationary_5 <= io_in_c_bypass_25_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_1_data_5 <= io_in_c_bypass_25_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_1_is_stationary_5 <= io_in_c_bypass_25_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_2_data_5 <= io_in_c_bypass_25_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_2_is_stationary_5 <= io_in_c_bypass_25_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_3_data_5 <= io_in_c_bypass_25_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_3_is_stationary_5 <= io_in_c_bypass_25_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_0_data_5 <= io_in_c_bypass_26_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_0_is_stationary_5 <= io_in_c_bypass_26_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_1_data_5 <= io_in_c_bypass_26_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_1_is_stationary_5 <= io_in_c_bypass_26_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_2_data_5 <= io_in_c_bypass_26_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_2_is_stationary_5 <= io_in_c_bypass_26_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_3_data_5 <= io_in_c_bypass_26_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_3_is_stationary_5 <= io_in_c_bypass_26_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_0_data_5 <= io_in_c_bypass_27_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_0_is_stationary_5 <= io_in_c_bypass_27_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_1_data_5 <= io_in_c_bypass_27_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_1_is_stationary_5 <= io_in_c_bypass_27_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_2_data_5 <= io_in_c_bypass_27_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_2_is_stationary_5 <= io_in_c_bypass_27_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_3_data_5 <= io_in_c_bypass_27_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_3_is_stationary_5 <= io_in_c_bypass_27_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_0_data_5 <= io_in_c_bypass_28_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_0_is_stationary_5 <= io_in_c_bypass_28_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_1_data_5 <= io_in_c_bypass_28_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_1_is_stationary_5 <= io_in_c_bypass_28_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_2_data_5 <= io_in_c_bypass_28_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_2_is_stationary_5 <= io_in_c_bypass_28_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_3_data_5 <= io_in_c_bypass_28_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_3_is_stationary_5 <= io_in_c_bypass_28_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_0_data_5 <= io_in_c_bypass_29_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_0_is_stationary_5 <= io_in_c_bypass_29_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_1_data_5 <= io_in_c_bypass_29_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_1_is_stationary_5 <= io_in_c_bypass_29_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_2_data_5 <= io_in_c_bypass_29_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_2_is_stationary_5 <= io_in_c_bypass_29_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_3_data_5 <= io_in_c_bypass_29_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_3_is_stationary_5 <= io_in_c_bypass_29_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_0_data_5 <= io_in_c_bypass_30_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_0_is_stationary_5 <= io_in_c_bypass_30_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_1_data_5 <= io_in_c_bypass_30_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_1_is_stationary_5 <= io_in_c_bypass_30_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_2_data_5 <= io_in_c_bypass_30_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_2_is_stationary_5 <= io_in_c_bypass_30_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_3_data_5 <= io_in_c_bypass_30_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_3_is_stationary_5 <= io_in_c_bypass_30_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_0_data_5 <= io_in_c_bypass_31_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_0_is_stationary_5 <= io_in_c_bypass_31_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_1_data_5 <= io_in_c_bypass_31_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_1_is_stationary_5 <= io_in_c_bypass_31_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_2_data_5 <= io_in_c_bypass_31_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_2_is_stationary_5 <= io_in_c_bypass_31_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_3_data_5 <= io_in_c_bypass_31_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_3_is_stationary_5 <= io_in_c_bypass_31_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_0_data_6 <= io_in_c_bypass_0_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_0_is_stationary_6 <= io_in_c_bypass_0_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_1_data_6 <= io_in_c_bypass_0_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_1_is_stationary_6 <= io_in_c_bypass_0_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_2_data_6 <= io_in_c_bypass_0_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_2_is_stationary_6 <= io_in_c_bypass_0_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_3_data_6 <= io_in_c_bypass_0_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_3_is_stationary_6 <= io_in_c_bypass_0_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_0_data_6 <= io_in_c_bypass_1_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_0_is_stationary_6 <= io_in_c_bypass_1_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_1_data_6 <= io_in_c_bypass_1_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_1_is_stationary_6 <= io_in_c_bypass_1_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_2_data_6 <= io_in_c_bypass_1_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_2_is_stationary_6 <= io_in_c_bypass_1_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_3_data_6 <= io_in_c_bypass_1_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_3_is_stationary_6 <= io_in_c_bypass_1_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_0_data_6 <= io_in_c_bypass_2_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_0_is_stationary_6 <= io_in_c_bypass_2_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_1_data_6 <= io_in_c_bypass_2_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_1_is_stationary_6 <= io_in_c_bypass_2_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_2_data_6 <= io_in_c_bypass_2_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_2_is_stationary_6 <= io_in_c_bypass_2_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_3_data_6 <= io_in_c_bypass_2_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_3_is_stationary_6 <= io_in_c_bypass_2_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_0_data_6 <= io_in_c_bypass_3_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_0_is_stationary_6 <= io_in_c_bypass_3_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_1_data_6 <= io_in_c_bypass_3_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_1_is_stationary_6 <= io_in_c_bypass_3_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_2_data_6 <= io_in_c_bypass_3_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_2_is_stationary_6 <= io_in_c_bypass_3_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_3_data_6 <= io_in_c_bypass_3_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_3_is_stationary_6 <= io_in_c_bypass_3_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_0_data_6 <= io_in_c_bypass_4_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_0_is_stationary_6 <= io_in_c_bypass_4_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_1_data_6 <= io_in_c_bypass_4_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_1_is_stationary_6 <= io_in_c_bypass_4_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_2_data_6 <= io_in_c_bypass_4_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_2_is_stationary_6 <= io_in_c_bypass_4_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_3_data_6 <= io_in_c_bypass_4_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_3_is_stationary_6 <= io_in_c_bypass_4_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_0_data_6 <= io_in_c_bypass_5_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_0_is_stationary_6 <= io_in_c_bypass_5_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_1_data_6 <= io_in_c_bypass_5_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_1_is_stationary_6 <= io_in_c_bypass_5_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_2_data_6 <= io_in_c_bypass_5_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_2_is_stationary_6 <= io_in_c_bypass_5_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_3_data_6 <= io_in_c_bypass_5_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_3_is_stationary_6 <= io_in_c_bypass_5_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_0_data_6 <= io_in_c_bypass_6_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_0_is_stationary_6 <= io_in_c_bypass_6_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_1_data_6 <= io_in_c_bypass_6_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_1_is_stationary_6 <= io_in_c_bypass_6_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_2_data_6 <= io_in_c_bypass_6_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_2_is_stationary_6 <= io_in_c_bypass_6_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_3_data_6 <= io_in_c_bypass_6_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_3_is_stationary_6 <= io_in_c_bypass_6_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_0_data_6 <= io_in_c_bypass_7_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_0_is_stationary_6 <= io_in_c_bypass_7_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_1_data_6 <= io_in_c_bypass_7_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_1_is_stationary_6 <= io_in_c_bypass_7_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_2_data_6 <= io_in_c_bypass_7_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_2_is_stationary_6 <= io_in_c_bypass_7_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_3_data_6 <= io_in_c_bypass_7_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_3_is_stationary_6 <= io_in_c_bypass_7_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_0_data_6 <= io_in_c_bypass_8_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_0_is_stationary_6 <= io_in_c_bypass_8_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_1_data_6 <= io_in_c_bypass_8_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_1_is_stationary_6 <= io_in_c_bypass_8_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_2_data_6 <= io_in_c_bypass_8_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_2_is_stationary_6 <= io_in_c_bypass_8_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_3_data_6 <= io_in_c_bypass_8_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_3_is_stationary_6 <= io_in_c_bypass_8_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_0_data_6 <= io_in_c_bypass_9_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_0_is_stationary_6 <= io_in_c_bypass_9_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_1_data_6 <= io_in_c_bypass_9_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_1_is_stationary_6 <= io_in_c_bypass_9_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_2_data_6 <= io_in_c_bypass_9_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_2_is_stationary_6 <= io_in_c_bypass_9_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_3_data_6 <= io_in_c_bypass_9_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_3_is_stationary_6 <= io_in_c_bypass_9_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_0_data_6 <= io_in_c_bypass_10_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_0_is_stationary_6 <= io_in_c_bypass_10_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_1_data_6 <= io_in_c_bypass_10_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_1_is_stationary_6 <= io_in_c_bypass_10_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_2_data_6 <= io_in_c_bypass_10_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_2_is_stationary_6 <= io_in_c_bypass_10_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_3_data_6 <= io_in_c_bypass_10_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_3_is_stationary_6 <= io_in_c_bypass_10_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_0_data_6 <= io_in_c_bypass_11_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_0_is_stationary_6 <= io_in_c_bypass_11_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_1_data_6 <= io_in_c_bypass_11_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_1_is_stationary_6 <= io_in_c_bypass_11_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_2_data_6 <= io_in_c_bypass_11_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_2_is_stationary_6 <= io_in_c_bypass_11_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_3_data_6 <= io_in_c_bypass_11_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_3_is_stationary_6 <= io_in_c_bypass_11_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_0_data_6 <= io_in_c_bypass_12_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_0_is_stationary_6 <= io_in_c_bypass_12_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_1_data_6 <= io_in_c_bypass_12_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_1_is_stationary_6 <= io_in_c_bypass_12_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_2_data_6 <= io_in_c_bypass_12_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_2_is_stationary_6 <= io_in_c_bypass_12_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_3_data_6 <= io_in_c_bypass_12_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_3_is_stationary_6 <= io_in_c_bypass_12_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_0_data_6 <= io_in_c_bypass_13_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_0_is_stationary_6 <= io_in_c_bypass_13_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_1_data_6 <= io_in_c_bypass_13_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_1_is_stationary_6 <= io_in_c_bypass_13_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_2_data_6 <= io_in_c_bypass_13_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_2_is_stationary_6 <= io_in_c_bypass_13_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_3_data_6 <= io_in_c_bypass_13_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_3_is_stationary_6 <= io_in_c_bypass_13_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_0_data_6 <= io_in_c_bypass_14_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_0_is_stationary_6 <= io_in_c_bypass_14_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_1_data_6 <= io_in_c_bypass_14_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_1_is_stationary_6 <= io_in_c_bypass_14_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_2_data_6 <= io_in_c_bypass_14_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_2_is_stationary_6 <= io_in_c_bypass_14_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_3_data_6 <= io_in_c_bypass_14_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_3_is_stationary_6 <= io_in_c_bypass_14_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_0_data_6 <= io_in_c_bypass_15_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_0_is_stationary_6 <= io_in_c_bypass_15_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_1_data_6 <= io_in_c_bypass_15_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_1_is_stationary_6 <= io_in_c_bypass_15_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_2_data_6 <= io_in_c_bypass_15_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_2_is_stationary_6 <= io_in_c_bypass_15_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_3_data_6 <= io_in_c_bypass_15_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_3_is_stationary_6 <= io_in_c_bypass_15_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_0_data_6 <= io_in_c_bypass_16_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_0_is_stationary_6 <= io_in_c_bypass_16_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_1_data_6 <= io_in_c_bypass_16_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_1_is_stationary_6 <= io_in_c_bypass_16_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_2_data_6 <= io_in_c_bypass_16_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_2_is_stationary_6 <= io_in_c_bypass_16_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_3_data_6 <= io_in_c_bypass_16_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_3_is_stationary_6 <= io_in_c_bypass_16_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_0_data_6 <= io_in_c_bypass_17_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_0_is_stationary_6 <= io_in_c_bypass_17_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_1_data_6 <= io_in_c_bypass_17_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_1_is_stationary_6 <= io_in_c_bypass_17_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_2_data_6 <= io_in_c_bypass_17_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_2_is_stationary_6 <= io_in_c_bypass_17_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_3_data_6 <= io_in_c_bypass_17_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_3_is_stationary_6 <= io_in_c_bypass_17_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_0_data_6 <= io_in_c_bypass_18_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_0_is_stationary_6 <= io_in_c_bypass_18_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_1_data_6 <= io_in_c_bypass_18_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_1_is_stationary_6 <= io_in_c_bypass_18_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_2_data_6 <= io_in_c_bypass_18_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_2_is_stationary_6 <= io_in_c_bypass_18_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_3_data_6 <= io_in_c_bypass_18_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_3_is_stationary_6 <= io_in_c_bypass_18_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_0_data_6 <= io_in_c_bypass_19_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_0_is_stationary_6 <= io_in_c_bypass_19_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_1_data_6 <= io_in_c_bypass_19_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_1_is_stationary_6 <= io_in_c_bypass_19_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_2_data_6 <= io_in_c_bypass_19_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_2_is_stationary_6 <= io_in_c_bypass_19_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_3_data_6 <= io_in_c_bypass_19_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_3_is_stationary_6 <= io_in_c_bypass_19_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_0_data_6 <= io_in_c_bypass_20_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_0_is_stationary_6 <= io_in_c_bypass_20_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_1_data_6 <= io_in_c_bypass_20_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_1_is_stationary_6 <= io_in_c_bypass_20_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_2_data_6 <= io_in_c_bypass_20_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_2_is_stationary_6 <= io_in_c_bypass_20_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_3_data_6 <= io_in_c_bypass_20_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_3_is_stationary_6 <= io_in_c_bypass_20_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_0_data_6 <= io_in_c_bypass_21_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_0_is_stationary_6 <= io_in_c_bypass_21_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_1_data_6 <= io_in_c_bypass_21_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_1_is_stationary_6 <= io_in_c_bypass_21_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_2_data_6 <= io_in_c_bypass_21_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_2_is_stationary_6 <= io_in_c_bypass_21_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_3_data_6 <= io_in_c_bypass_21_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_3_is_stationary_6 <= io_in_c_bypass_21_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_0_data_6 <= io_in_c_bypass_22_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_0_is_stationary_6 <= io_in_c_bypass_22_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_1_data_6 <= io_in_c_bypass_22_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_1_is_stationary_6 <= io_in_c_bypass_22_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_2_data_6 <= io_in_c_bypass_22_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_2_is_stationary_6 <= io_in_c_bypass_22_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_3_data_6 <= io_in_c_bypass_22_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_3_is_stationary_6 <= io_in_c_bypass_22_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_0_data_6 <= io_in_c_bypass_23_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_0_is_stationary_6 <= io_in_c_bypass_23_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_1_data_6 <= io_in_c_bypass_23_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_1_is_stationary_6 <= io_in_c_bypass_23_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_2_data_6 <= io_in_c_bypass_23_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_2_is_stationary_6 <= io_in_c_bypass_23_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_3_data_6 <= io_in_c_bypass_23_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_3_is_stationary_6 <= io_in_c_bypass_23_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_0_data_6 <= io_in_c_bypass_24_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_0_is_stationary_6 <= io_in_c_bypass_24_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_1_data_6 <= io_in_c_bypass_24_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_1_is_stationary_6 <= io_in_c_bypass_24_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_2_data_6 <= io_in_c_bypass_24_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_2_is_stationary_6 <= io_in_c_bypass_24_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_3_data_6 <= io_in_c_bypass_24_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_3_is_stationary_6 <= io_in_c_bypass_24_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_0_data_6 <= io_in_c_bypass_25_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_0_is_stationary_6 <= io_in_c_bypass_25_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_1_data_6 <= io_in_c_bypass_25_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_1_is_stationary_6 <= io_in_c_bypass_25_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_2_data_6 <= io_in_c_bypass_25_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_2_is_stationary_6 <= io_in_c_bypass_25_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_3_data_6 <= io_in_c_bypass_25_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_3_is_stationary_6 <= io_in_c_bypass_25_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_0_data_6 <= io_in_c_bypass_26_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_0_is_stationary_6 <= io_in_c_bypass_26_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_1_data_6 <= io_in_c_bypass_26_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_1_is_stationary_6 <= io_in_c_bypass_26_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_2_data_6 <= io_in_c_bypass_26_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_2_is_stationary_6 <= io_in_c_bypass_26_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_3_data_6 <= io_in_c_bypass_26_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_3_is_stationary_6 <= io_in_c_bypass_26_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_0_data_6 <= io_in_c_bypass_27_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_0_is_stationary_6 <= io_in_c_bypass_27_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_1_data_6 <= io_in_c_bypass_27_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_1_is_stationary_6 <= io_in_c_bypass_27_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_2_data_6 <= io_in_c_bypass_27_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_2_is_stationary_6 <= io_in_c_bypass_27_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_3_data_6 <= io_in_c_bypass_27_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_3_is_stationary_6 <= io_in_c_bypass_27_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_0_data_6 <= io_in_c_bypass_28_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_0_is_stationary_6 <= io_in_c_bypass_28_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_1_data_6 <= io_in_c_bypass_28_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_1_is_stationary_6 <= io_in_c_bypass_28_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_2_data_6 <= io_in_c_bypass_28_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_2_is_stationary_6 <= io_in_c_bypass_28_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_3_data_6 <= io_in_c_bypass_28_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_3_is_stationary_6 <= io_in_c_bypass_28_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_0_data_6 <= io_in_c_bypass_29_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_0_is_stationary_6 <= io_in_c_bypass_29_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_1_data_6 <= io_in_c_bypass_29_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_1_is_stationary_6 <= io_in_c_bypass_29_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_2_data_6 <= io_in_c_bypass_29_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_2_is_stationary_6 <= io_in_c_bypass_29_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_3_data_6 <= io_in_c_bypass_29_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_3_is_stationary_6 <= io_in_c_bypass_29_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_0_data_6 <= io_in_c_bypass_30_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_0_is_stationary_6 <= io_in_c_bypass_30_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_1_data_6 <= io_in_c_bypass_30_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_1_is_stationary_6 <= io_in_c_bypass_30_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_2_data_6 <= io_in_c_bypass_30_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_2_is_stationary_6 <= io_in_c_bypass_30_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_3_data_6 <= io_in_c_bypass_30_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_3_is_stationary_6 <= io_in_c_bypass_30_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_0_data_6 <= io_in_c_bypass_31_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_0_is_stationary_6 <= io_in_c_bypass_31_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_1_data_6 <= io_in_c_bypass_31_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_1_is_stationary_6 <= io_in_c_bypass_31_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_2_data_6 <= io_in_c_bypass_31_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_2_is_stationary_6 <= io_in_c_bypass_31_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_3_data_6 <= io_in_c_bypass_31_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_3_is_stationary_6 <= io_in_c_bypass_31_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_0_data_7 <= io_in_c_bypass_0_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_0_is_stationary_7 <= io_in_c_bypass_0_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_1_data_7 <= io_in_c_bypass_0_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_1_is_stationary_7 <= io_in_c_bypass_0_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_2_data_7 <= io_in_c_bypass_0_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_2_is_stationary_7 <= io_in_c_bypass_0_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_3_data_7 <= io_in_c_bypass_0_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_3_is_stationary_7 <= io_in_c_bypass_0_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_0_data_7 <= io_in_c_bypass_1_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_0_is_stationary_7 <= io_in_c_bypass_1_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_1_data_7 <= io_in_c_bypass_1_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_1_is_stationary_7 <= io_in_c_bypass_1_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_2_data_7 <= io_in_c_bypass_1_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_2_is_stationary_7 <= io_in_c_bypass_1_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_3_data_7 <= io_in_c_bypass_1_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_3_is_stationary_7 <= io_in_c_bypass_1_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_0_data_7 <= io_in_c_bypass_2_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_0_is_stationary_7 <= io_in_c_bypass_2_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_1_data_7 <= io_in_c_bypass_2_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_1_is_stationary_7 <= io_in_c_bypass_2_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_2_data_7 <= io_in_c_bypass_2_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_2_is_stationary_7 <= io_in_c_bypass_2_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_3_data_7 <= io_in_c_bypass_2_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_3_is_stationary_7 <= io_in_c_bypass_2_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_0_data_7 <= io_in_c_bypass_3_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_0_is_stationary_7 <= io_in_c_bypass_3_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_1_data_7 <= io_in_c_bypass_3_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_1_is_stationary_7 <= io_in_c_bypass_3_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_2_data_7 <= io_in_c_bypass_3_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_2_is_stationary_7 <= io_in_c_bypass_3_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_3_data_7 <= io_in_c_bypass_3_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_3_is_stationary_7 <= io_in_c_bypass_3_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_0_data_7 <= io_in_c_bypass_4_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_0_is_stationary_7 <= io_in_c_bypass_4_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_1_data_7 <= io_in_c_bypass_4_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_1_is_stationary_7 <= io_in_c_bypass_4_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_2_data_7 <= io_in_c_bypass_4_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_2_is_stationary_7 <= io_in_c_bypass_4_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_3_data_7 <= io_in_c_bypass_4_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_3_is_stationary_7 <= io_in_c_bypass_4_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_0_data_7 <= io_in_c_bypass_5_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_0_is_stationary_7 <= io_in_c_bypass_5_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_1_data_7 <= io_in_c_bypass_5_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_1_is_stationary_7 <= io_in_c_bypass_5_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_2_data_7 <= io_in_c_bypass_5_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_2_is_stationary_7 <= io_in_c_bypass_5_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_3_data_7 <= io_in_c_bypass_5_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_3_is_stationary_7 <= io_in_c_bypass_5_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_0_data_7 <= io_in_c_bypass_6_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_0_is_stationary_7 <= io_in_c_bypass_6_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_1_data_7 <= io_in_c_bypass_6_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_1_is_stationary_7 <= io_in_c_bypass_6_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_2_data_7 <= io_in_c_bypass_6_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_2_is_stationary_7 <= io_in_c_bypass_6_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_3_data_7 <= io_in_c_bypass_6_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_3_is_stationary_7 <= io_in_c_bypass_6_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_0_data_7 <= io_in_c_bypass_7_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_0_is_stationary_7 <= io_in_c_bypass_7_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_1_data_7 <= io_in_c_bypass_7_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_1_is_stationary_7 <= io_in_c_bypass_7_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_2_data_7 <= io_in_c_bypass_7_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_2_is_stationary_7 <= io_in_c_bypass_7_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_3_data_7 <= io_in_c_bypass_7_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_3_is_stationary_7 <= io_in_c_bypass_7_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_0_data_7 <= io_in_c_bypass_8_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_0_is_stationary_7 <= io_in_c_bypass_8_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_1_data_7 <= io_in_c_bypass_8_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_1_is_stationary_7 <= io_in_c_bypass_8_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_2_data_7 <= io_in_c_bypass_8_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_2_is_stationary_7 <= io_in_c_bypass_8_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_3_data_7 <= io_in_c_bypass_8_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_3_is_stationary_7 <= io_in_c_bypass_8_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_0_data_7 <= io_in_c_bypass_9_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_0_is_stationary_7 <= io_in_c_bypass_9_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_1_data_7 <= io_in_c_bypass_9_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_1_is_stationary_7 <= io_in_c_bypass_9_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_2_data_7 <= io_in_c_bypass_9_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_2_is_stationary_7 <= io_in_c_bypass_9_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_3_data_7 <= io_in_c_bypass_9_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_3_is_stationary_7 <= io_in_c_bypass_9_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_0_data_7 <= io_in_c_bypass_10_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_0_is_stationary_7 <= io_in_c_bypass_10_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_1_data_7 <= io_in_c_bypass_10_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_1_is_stationary_7 <= io_in_c_bypass_10_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_2_data_7 <= io_in_c_bypass_10_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_2_is_stationary_7 <= io_in_c_bypass_10_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_3_data_7 <= io_in_c_bypass_10_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_3_is_stationary_7 <= io_in_c_bypass_10_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_0_data_7 <= io_in_c_bypass_11_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_0_is_stationary_7 <= io_in_c_bypass_11_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_1_data_7 <= io_in_c_bypass_11_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_1_is_stationary_7 <= io_in_c_bypass_11_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_2_data_7 <= io_in_c_bypass_11_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_2_is_stationary_7 <= io_in_c_bypass_11_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_3_data_7 <= io_in_c_bypass_11_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_3_is_stationary_7 <= io_in_c_bypass_11_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_0_data_7 <= io_in_c_bypass_12_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_0_is_stationary_7 <= io_in_c_bypass_12_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_1_data_7 <= io_in_c_bypass_12_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_1_is_stationary_7 <= io_in_c_bypass_12_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_2_data_7 <= io_in_c_bypass_12_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_2_is_stationary_7 <= io_in_c_bypass_12_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_3_data_7 <= io_in_c_bypass_12_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_3_is_stationary_7 <= io_in_c_bypass_12_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_0_data_7 <= io_in_c_bypass_13_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_0_is_stationary_7 <= io_in_c_bypass_13_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_1_data_7 <= io_in_c_bypass_13_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_1_is_stationary_7 <= io_in_c_bypass_13_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_2_data_7 <= io_in_c_bypass_13_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_2_is_stationary_7 <= io_in_c_bypass_13_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_3_data_7 <= io_in_c_bypass_13_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_3_is_stationary_7 <= io_in_c_bypass_13_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_0_data_7 <= io_in_c_bypass_14_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_0_is_stationary_7 <= io_in_c_bypass_14_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_1_data_7 <= io_in_c_bypass_14_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_1_is_stationary_7 <= io_in_c_bypass_14_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_2_data_7 <= io_in_c_bypass_14_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_2_is_stationary_7 <= io_in_c_bypass_14_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_3_data_7 <= io_in_c_bypass_14_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_3_is_stationary_7 <= io_in_c_bypass_14_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_0_data_7 <= io_in_c_bypass_15_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_0_is_stationary_7 <= io_in_c_bypass_15_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_1_data_7 <= io_in_c_bypass_15_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_1_is_stationary_7 <= io_in_c_bypass_15_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_2_data_7 <= io_in_c_bypass_15_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_2_is_stationary_7 <= io_in_c_bypass_15_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_3_data_7 <= io_in_c_bypass_15_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_3_is_stationary_7 <= io_in_c_bypass_15_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_0_data_7 <= io_in_c_bypass_16_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_0_is_stationary_7 <= io_in_c_bypass_16_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_1_data_7 <= io_in_c_bypass_16_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_1_is_stationary_7 <= io_in_c_bypass_16_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_2_data_7 <= io_in_c_bypass_16_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_2_is_stationary_7 <= io_in_c_bypass_16_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_3_data_7 <= io_in_c_bypass_16_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_3_is_stationary_7 <= io_in_c_bypass_16_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_0_data_7 <= io_in_c_bypass_17_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_0_is_stationary_7 <= io_in_c_bypass_17_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_1_data_7 <= io_in_c_bypass_17_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_1_is_stationary_7 <= io_in_c_bypass_17_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_2_data_7 <= io_in_c_bypass_17_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_2_is_stationary_7 <= io_in_c_bypass_17_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_3_data_7 <= io_in_c_bypass_17_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_3_is_stationary_7 <= io_in_c_bypass_17_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_0_data_7 <= io_in_c_bypass_18_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_0_is_stationary_7 <= io_in_c_bypass_18_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_1_data_7 <= io_in_c_bypass_18_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_1_is_stationary_7 <= io_in_c_bypass_18_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_2_data_7 <= io_in_c_bypass_18_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_2_is_stationary_7 <= io_in_c_bypass_18_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_3_data_7 <= io_in_c_bypass_18_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_3_is_stationary_7 <= io_in_c_bypass_18_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_0_data_7 <= io_in_c_bypass_19_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_0_is_stationary_7 <= io_in_c_bypass_19_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_1_data_7 <= io_in_c_bypass_19_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_1_is_stationary_7 <= io_in_c_bypass_19_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_2_data_7 <= io_in_c_bypass_19_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_2_is_stationary_7 <= io_in_c_bypass_19_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_3_data_7 <= io_in_c_bypass_19_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_3_is_stationary_7 <= io_in_c_bypass_19_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_0_data_7 <= io_in_c_bypass_20_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_0_is_stationary_7 <= io_in_c_bypass_20_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_1_data_7 <= io_in_c_bypass_20_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_1_is_stationary_7 <= io_in_c_bypass_20_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_2_data_7 <= io_in_c_bypass_20_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_2_is_stationary_7 <= io_in_c_bypass_20_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_3_data_7 <= io_in_c_bypass_20_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_3_is_stationary_7 <= io_in_c_bypass_20_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_0_data_7 <= io_in_c_bypass_21_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_0_is_stationary_7 <= io_in_c_bypass_21_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_1_data_7 <= io_in_c_bypass_21_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_1_is_stationary_7 <= io_in_c_bypass_21_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_2_data_7 <= io_in_c_bypass_21_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_2_is_stationary_7 <= io_in_c_bypass_21_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_3_data_7 <= io_in_c_bypass_21_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_3_is_stationary_7 <= io_in_c_bypass_21_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_0_data_7 <= io_in_c_bypass_22_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_0_is_stationary_7 <= io_in_c_bypass_22_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_1_data_7 <= io_in_c_bypass_22_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_1_is_stationary_7 <= io_in_c_bypass_22_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_2_data_7 <= io_in_c_bypass_22_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_2_is_stationary_7 <= io_in_c_bypass_22_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_3_data_7 <= io_in_c_bypass_22_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_3_is_stationary_7 <= io_in_c_bypass_22_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_0_data_7 <= io_in_c_bypass_23_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_0_is_stationary_7 <= io_in_c_bypass_23_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_1_data_7 <= io_in_c_bypass_23_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_1_is_stationary_7 <= io_in_c_bypass_23_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_2_data_7 <= io_in_c_bypass_23_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_2_is_stationary_7 <= io_in_c_bypass_23_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_3_data_7 <= io_in_c_bypass_23_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_3_is_stationary_7 <= io_in_c_bypass_23_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_0_data_7 <= io_in_c_bypass_24_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_0_is_stationary_7 <= io_in_c_bypass_24_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_1_data_7 <= io_in_c_bypass_24_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_1_is_stationary_7 <= io_in_c_bypass_24_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_2_data_7 <= io_in_c_bypass_24_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_2_is_stationary_7 <= io_in_c_bypass_24_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_3_data_7 <= io_in_c_bypass_24_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_3_is_stationary_7 <= io_in_c_bypass_24_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_0_data_7 <= io_in_c_bypass_25_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_0_is_stationary_7 <= io_in_c_bypass_25_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_1_data_7 <= io_in_c_bypass_25_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_1_is_stationary_7 <= io_in_c_bypass_25_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_2_data_7 <= io_in_c_bypass_25_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_2_is_stationary_7 <= io_in_c_bypass_25_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_3_data_7 <= io_in_c_bypass_25_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_3_is_stationary_7 <= io_in_c_bypass_25_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_0_data_7 <= io_in_c_bypass_26_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_0_is_stationary_7 <= io_in_c_bypass_26_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_1_data_7 <= io_in_c_bypass_26_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_1_is_stationary_7 <= io_in_c_bypass_26_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_2_data_7 <= io_in_c_bypass_26_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_2_is_stationary_7 <= io_in_c_bypass_26_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_3_data_7 <= io_in_c_bypass_26_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_3_is_stationary_7 <= io_in_c_bypass_26_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_0_data_7 <= io_in_c_bypass_27_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_0_is_stationary_7 <= io_in_c_bypass_27_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_1_data_7 <= io_in_c_bypass_27_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_1_is_stationary_7 <= io_in_c_bypass_27_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_2_data_7 <= io_in_c_bypass_27_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_2_is_stationary_7 <= io_in_c_bypass_27_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_3_data_7 <= io_in_c_bypass_27_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_3_is_stationary_7 <= io_in_c_bypass_27_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_0_data_7 <= io_in_c_bypass_28_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_0_is_stationary_7 <= io_in_c_bypass_28_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_1_data_7 <= io_in_c_bypass_28_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_1_is_stationary_7 <= io_in_c_bypass_28_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_2_data_7 <= io_in_c_bypass_28_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_2_is_stationary_7 <= io_in_c_bypass_28_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_3_data_7 <= io_in_c_bypass_28_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_3_is_stationary_7 <= io_in_c_bypass_28_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_0_data_7 <= io_in_c_bypass_29_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_0_is_stationary_7 <= io_in_c_bypass_29_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_1_data_7 <= io_in_c_bypass_29_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_1_is_stationary_7 <= io_in_c_bypass_29_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_2_data_7 <= io_in_c_bypass_29_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_2_is_stationary_7 <= io_in_c_bypass_29_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_3_data_7 <= io_in_c_bypass_29_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_3_is_stationary_7 <= io_in_c_bypass_29_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_0_data_7 <= io_in_c_bypass_30_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_0_is_stationary_7 <= io_in_c_bypass_30_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_1_data_7 <= io_in_c_bypass_30_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_1_is_stationary_7 <= io_in_c_bypass_30_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_2_data_7 <= io_in_c_bypass_30_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_2_is_stationary_7 <= io_in_c_bypass_30_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_3_data_7 <= io_in_c_bypass_30_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_3_is_stationary_7 <= io_in_c_bypass_30_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_0_data_7 <= io_in_c_bypass_31_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_0_is_stationary_7 <= io_in_c_bypass_31_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_1_data_7 <= io_in_c_bypass_31_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_1_is_stationary_7 <= io_in_c_bypass_31_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_2_data_7 <= io_in_c_bypass_31_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_2_is_stationary_7 <= io_in_c_bypass_31_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_3_data_7 <= io_in_c_bypass_31_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_3_is_stationary_7 <= io_in_c_bypass_31_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_0_data_8 <= io_in_c_bypass_0_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_0_is_stationary_8 <= io_in_c_bypass_0_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_1_data_8 <= io_in_c_bypass_0_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_1_is_stationary_8 <= io_in_c_bypass_0_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_2_data_8 <= io_in_c_bypass_0_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_2_is_stationary_8 <= io_in_c_bypass_0_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_3_data_8 <= io_in_c_bypass_0_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_3_is_stationary_8 <= io_in_c_bypass_0_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_0_data_8 <= io_in_c_bypass_1_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_0_is_stationary_8 <= io_in_c_bypass_1_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_1_data_8 <= io_in_c_bypass_1_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_1_is_stationary_8 <= io_in_c_bypass_1_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_2_data_8 <= io_in_c_bypass_1_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_2_is_stationary_8 <= io_in_c_bypass_1_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_3_data_8 <= io_in_c_bypass_1_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_3_is_stationary_8 <= io_in_c_bypass_1_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_0_data_8 <= io_in_c_bypass_2_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_0_is_stationary_8 <= io_in_c_bypass_2_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_1_data_8 <= io_in_c_bypass_2_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_1_is_stationary_8 <= io_in_c_bypass_2_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_2_data_8 <= io_in_c_bypass_2_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_2_is_stationary_8 <= io_in_c_bypass_2_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_3_data_8 <= io_in_c_bypass_2_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_3_is_stationary_8 <= io_in_c_bypass_2_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_0_data_8 <= io_in_c_bypass_3_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_0_is_stationary_8 <= io_in_c_bypass_3_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_1_data_8 <= io_in_c_bypass_3_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_1_is_stationary_8 <= io_in_c_bypass_3_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_2_data_8 <= io_in_c_bypass_3_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_2_is_stationary_8 <= io_in_c_bypass_3_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_3_data_8 <= io_in_c_bypass_3_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_3_is_stationary_8 <= io_in_c_bypass_3_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_0_data_8 <= io_in_c_bypass_4_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_0_is_stationary_8 <= io_in_c_bypass_4_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_1_data_8 <= io_in_c_bypass_4_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_1_is_stationary_8 <= io_in_c_bypass_4_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_2_data_8 <= io_in_c_bypass_4_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_2_is_stationary_8 <= io_in_c_bypass_4_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_3_data_8 <= io_in_c_bypass_4_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_3_is_stationary_8 <= io_in_c_bypass_4_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_0_data_8 <= io_in_c_bypass_5_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_0_is_stationary_8 <= io_in_c_bypass_5_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_1_data_8 <= io_in_c_bypass_5_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_1_is_stationary_8 <= io_in_c_bypass_5_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_2_data_8 <= io_in_c_bypass_5_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_2_is_stationary_8 <= io_in_c_bypass_5_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_3_data_8 <= io_in_c_bypass_5_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_3_is_stationary_8 <= io_in_c_bypass_5_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_0_data_8 <= io_in_c_bypass_6_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_0_is_stationary_8 <= io_in_c_bypass_6_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_1_data_8 <= io_in_c_bypass_6_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_1_is_stationary_8 <= io_in_c_bypass_6_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_2_data_8 <= io_in_c_bypass_6_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_2_is_stationary_8 <= io_in_c_bypass_6_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_3_data_8 <= io_in_c_bypass_6_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_3_is_stationary_8 <= io_in_c_bypass_6_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_0_data_8 <= io_in_c_bypass_7_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_0_is_stationary_8 <= io_in_c_bypass_7_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_1_data_8 <= io_in_c_bypass_7_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_1_is_stationary_8 <= io_in_c_bypass_7_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_2_data_8 <= io_in_c_bypass_7_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_2_is_stationary_8 <= io_in_c_bypass_7_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_3_data_8 <= io_in_c_bypass_7_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_3_is_stationary_8 <= io_in_c_bypass_7_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_0_data_8 <= io_in_c_bypass_8_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_0_is_stationary_8 <= io_in_c_bypass_8_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_1_data_8 <= io_in_c_bypass_8_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_1_is_stationary_8 <= io_in_c_bypass_8_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_2_data_8 <= io_in_c_bypass_8_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_2_is_stationary_8 <= io_in_c_bypass_8_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_3_data_8 <= io_in_c_bypass_8_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_3_is_stationary_8 <= io_in_c_bypass_8_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_0_data_8 <= io_in_c_bypass_9_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_0_is_stationary_8 <= io_in_c_bypass_9_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_1_data_8 <= io_in_c_bypass_9_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_1_is_stationary_8 <= io_in_c_bypass_9_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_2_data_8 <= io_in_c_bypass_9_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_2_is_stationary_8 <= io_in_c_bypass_9_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_3_data_8 <= io_in_c_bypass_9_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_3_is_stationary_8 <= io_in_c_bypass_9_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_0_data_8 <= io_in_c_bypass_10_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_0_is_stationary_8 <= io_in_c_bypass_10_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_1_data_8 <= io_in_c_bypass_10_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_1_is_stationary_8 <= io_in_c_bypass_10_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_2_data_8 <= io_in_c_bypass_10_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_2_is_stationary_8 <= io_in_c_bypass_10_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_3_data_8 <= io_in_c_bypass_10_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_3_is_stationary_8 <= io_in_c_bypass_10_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_0_data_8 <= io_in_c_bypass_11_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_0_is_stationary_8 <= io_in_c_bypass_11_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_1_data_8 <= io_in_c_bypass_11_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_1_is_stationary_8 <= io_in_c_bypass_11_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_2_data_8 <= io_in_c_bypass_11_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_2_is_stationary_8 <= io_in_c_bypass_11_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_3_data_8 <= io_in_c_bypass_11_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_3_is_stationary_8 <= io_in_c_bypass_11_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_0_data_8 <= io_in_c_bypass_12_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_0_is_stationary_8 <= io_in_c_bypass_12_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_1_data_8 <= io_in_c_bypass_12_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_1_is_stationary_8 <= io_in_c_bypass_12_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_2_data_8 <= io_in_c_bypass_12_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_2_is_stationary_8 <= io_in_c_bypass_12_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_3_data_8 <= io_in_c_bypass_12_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_3_is_stationary_8 <= io_in_c_bypass_12_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_0_data_8 <= io_in_c_bypass_13_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_0_is_stationary_8 <= io_in_c_bypass_13_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_1_data_8 <= io_in_c_bypass_13_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_1_is_stationary_8 <= io_in_c_bypass_13_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_2_data_8 <= io_in_c_bypass_13_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_2_is_stationary_8 <= io_in_c_bypass_13_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_3_data_8 <= io_in_c_bypass_13_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_3_is_stationary_8 <= io_in_c_bypass_13_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_0_data_8 <= io_in_c_bypass_14_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_0_is_stationary_8 <= io_in_c_bypass_14_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_1_data_8 <= io_in_c_bypass_14_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_1_is_stationary_8 <= io_in_c_bypass_14_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_2_data_8 <= io_in_c_bypass_14_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_2_is_stationary_8 <= io_in_c_bypass_14_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_3_data_8 <= io_in_c_bypass_14_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_3_is_stationary_8 <= io_in_c_bypass_14_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_0_data_8 <= io_in_c_bypass_15_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_0_is_stationary_8 <= io_in_c_bypass_15_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_1_data_8 <= io_in_c_bypass_15_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_1_is_stationary_8 <= io_in_c_bypass_15_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_2_data_8 <= io_in_c_bypass_15_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_2_is_stationary_8 <= io_in_c_bypass_15_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_3_data_8 <= io_in_c_bypass_15_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_3_is_stationary_8 <= io_in_c_bypass_15_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_0_data_8 <= io_in_c_bypass_16_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_0_is_stationary_8 <= io_in_c_bypass_16_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_1_data_8 <= io_in_c_bypass_16_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_1_is_stationary_8 <= io_in_c_bypass_16_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_2_data_8 <= io_in_c_bypass_16_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_2_is_stationary_8 <= io_in_c_bypass_16_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_3_data_8 <= io_in_c_bypass_16_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_3_is_stationary_8 <= io_in_c_bypass_16_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_0_data_8 <= io_in_c_bypass_17_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_0_is_stationary_8 <= io_in_c_bypass_17_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_1_data_8 <= io_in_c_bypass_17_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_1_is_stationary_8 <= io_in_c_bypass_17_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_2_data_8 <= io_in_c_bypass_17_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_2_is_stationary_8 <= io_in_c_bypass_17_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_3_data_8 <= io_in_c_bypass_17_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_3_is_stationary_8 <= io_in_c_bypass_17_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_0_data_8 <= io_in_c_bypass_18_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_0_is_stationary_8 <= io_in_c_bypass_18_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_1_data_8 <= io_in_c_bypass_18_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_1_is_stationary_8 <= io_in_c_bypass_18_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_2_data_8 <= io_in_c_bypass_18_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_2_is_stationary_8 <= io_in_c_bypass_18_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_3_data_8 <= io_in_c_bypass_18_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_3_is_stationary_8 <= io_in_c_bypass_18_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_0_data_8 <= io_in_c_bypass_19_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_0_is_stationary_8 <= io_in_c_bypass_19_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_1_data_8 <= io_in_c_bypass_19_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_1_is_stationary_8 <= io_in_c_bypass_19_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_2_data_8 <= io_in_c_bypass_19_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_2_is_stationary_8 <= io_in_c_bypass_19_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_3_data_8 <= io_in_c_bypass_19_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_3_is_stationary_8 <= io_in_c_bypass_19_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_0_data_8 <= io_in_c_bypass_20_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_0_is_stationary_8 <= io_in_c_bypass_20_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_1_data_8 <= io_in_c_bypass_20_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_1_is_stationary_8 <= io_in_c_bypass_20_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_2_data_8 <= io_in_c_bypass_20_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_2_is_stationary_8 <= io_in_c_bypass_20_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_3_data_8 <= io_in_c_bypass_20_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_3_is_stationary_8 <= io_in_c_bypass_20_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_0_data_8 <= io_in_c_bypass_21_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_0_is_stationary_8 <= io_in_c_bypass_21_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_1_data_8 <= io_in_c_bypass_21_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_1_is_stationary_8 <= io_in_c_bypass_21_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_2_data_8 <= io_in_c_bypass_21_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_2_is_stationary_8 <= io_in_c_bypass_21_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_3_data_8 <= io_in_c_bypass_21_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_3_is_stationary_8 <= io_in_c_bypass_21_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_0_data_8 <= io_in_c_bypass_22_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_0_is_stationary_8 <= io_in_c_bypass_22_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_1_data_8 <= io_in_c_bypass_22_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_1_is_stationary_8 <= io_in_c_bypass_22_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_2_data_8 <= io_in_c_bypass_22_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_2_is_stationary_8 <= io_in_c_bypass_22_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_3_data_8 <= io_in_c_bypass_22_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_3_is_stationary_8 <= io_in_c_bypass_22_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_0_data_8 <= io_in_c_bypass_23_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_0_is_stationary_8 <= io_in_c_bypass_23_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_1_data_8 <= io_in_c_bypass_23_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_1_is_stationary_8 <= io_in_c_bypass_23_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_2_data_8 <= io_in_c_bypass_23_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_2_is_stationary_8 <= io_in_c_bypass_23_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_3_data_8 <= io_in_c_bypass_23_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_3_is_stationary_8 <= io_in_c_bypass_23_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_0_data_8 <= io_in_c_bypass_24_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_0_is_stationary_8 <= io_in_c_bypass_24_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_1_data_8 <= io_in_c_bypass_24_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_1_is_stationary_8 <= io_in_c_bypass_24_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_2_data_8 <= io_in_c_bypass_24_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_2_is_stationary_8 <= io_in_c_bypass_24_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_3_data_8 <= io_in_c_bypass_24_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_3_is_stationary_8 <= io_in_c_bypass_24_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_0_data_8 <= io_in_c_bypass_25_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_0_is_stationary_8 <= io_in_c_bypass_25_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_1_data_8 <= io_in_c_bypass_25_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_1_is_stationary_8 <= io_in_c_bypass_25_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_2_data_8 <= io_in_c_bypass_25_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_2_is_stationary_8 <= io_in_c_bypass_25_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_3_data_8 <= io_in_c_bypass_25_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_3_is_stationary_8 <= io_in_c_bypass_25_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_0_data_8 <= io_in_c_bypass_26_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_0_is_stationary_8 <= io_in_c_bypass_26_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_1_data_8 <= io_in_c_bypass_26_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_1_is_stationary_8 <= io_in_c_bypass_26_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_2_data_8 <= io_in_c_bypass_26_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_2_is_stationary_8 <= io_in_c_bypass_26_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_3_data_8 <= io_in_c_bypass_26_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_3_is_stationary_8 <= io_in_c_bypass_26_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_0_data_8 <= io_in_c_bypass_27_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_0_is_stationary_8 <= io_in_c_bypass_27_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_1_data_8 <= io_in_c_bypass_27_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_1_is_stationary_8 <= io_in_c_bypass_27_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_2_data_8 <= io_in_c_bypass_27_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_2_is_stationary_8 <= io_in_c_bypass_27_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_3_data_8 <= io_in_c_bypass_27_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_3_is_stationary_8 <= io_in_c_bypass_27_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_0_data_8 <= io_in_c_bypass_28_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_0_is_stationary_8 <= io_in_c_bypass_28_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_1_data_8 <= io_in_c_bypass_28_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_1_is_stationary_8 <= io_in_c_bypass_28_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_2_data_8 <= io_in_c_bypass_28_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_2_is_stationary_8 <= io_in_c_bypass_28_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_3_data_8 <= io_in_c_bypass_28_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_3_is_stationary_8 <= io_in_c_bypass_28_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_0_data_8 <= io_in_c_bypass_29_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_0_is_stationary_8 <= io_in_c_bypass_29_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_1_data_8 <= io_in_c_bypass_29_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_1_is_stationary_8 <= io_in_c_bypass_29_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_2_data_8 <= io_in_c_bypass_29_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_2_is_stationary_8 <= io_in_c_bypass_29_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_3_data_8 <= io_in_c_bypass_29_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_3_is_stationary_8 <= io_in_c_bypass_29_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_0_data_8 <= io_in_c_bypass_30_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_0_is_stationary_8 <= io_in_c_bypass_30_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_1_data_8 <= io_in_c_bypass_30_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_1_is_stationary_8 <= io_in_c_bypass_30_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_2_data_8 <= io_in_c_bypass_30_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_2_is_stationary_8 <= io_in_c_bypass_30_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_3_data_8 <= io_in_c_bypass_30_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_3_is_stationary_8 <= io_in_c_bypass_30_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_0_data_8 <= io_in_c_bypass_31_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_0_is_stationary_8 <= io_in_c_bypass_31_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_1_data_8 <= io_in_c_bypass_31_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_1_is_stationary_8 <= io_in_c_bypass_31_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_2_data_8 <= io_in_c_bypass_31_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_2_is_stationary_8 <= io_in_c_bypass_31_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_3_data_8 <= io_in_c_bypass_31_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_3_is_stationary_8 <= io_in_c_bypass_31_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_0_data_9 <= io_in_c_bypass_0_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_0_is_stationary_9 <= io_in_c_bypass_0_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_1_data_9 <= io_in_c_bypass_0_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_1_is_stationary_9 <= io_in_c_bypass_0_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_2_data_9 <= io_in_c_bypass_0_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_2_is_stationary_9 <= io_in_c_bypass_0_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_3_data_9 <= io_in_c_bypass_0_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_3_is_stationary_9 <= io_in_c_bypass_0_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_0_data_9 <= io_in_c_bypass_1_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_0_is_stationary_9 <= io_in_c_bypass_1_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_1_data_9 <= io_in_c_bypass_1_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_1_is_stationary_9 <= io_in_c_bypass_1_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_2_data_9 <= io_in_c_bypass_1_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_2_is_stationary_9 <= io_in_c_bypass_1_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_3_data_9 <= io_in_c_bypass_1_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_3_is_stationary_9 <= io_in_c_bypass_1_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_0_data_9 <= io_in_c_bypass_2_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_0_is_stationary_9 <= io_in_c_bypass_2_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_1_data_9 <= io_in_c_bypass_2_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_1_is_stationary_9 <= io_in_c_bypass_2_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_2_data_9 <= io_in_c_bypass_2_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_2_is_stationary_9 <= io_in_c_bypass_2_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_3_data_9 <= io_in_c_bypass_2_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_3_is_stationary_9 <= io_in_c_bypass_2_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_0_data_9 <= io_in_c_bypass_3_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_0_is_stationary_9 <= io_in_c_bypass_3_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_1_data_9 <= io_in_c_bypass_3_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_1_is_stationary_9 <= io_in_c_bypass_3_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_2_data_9 <= io_in_c_bypass_3_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_2_is_stationary_9 <= io_in_c_bypass_3_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_3_data_9 <= io_in_c_bypass_3_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_3_is_stationary_9 <= io_in_c_bypass_3_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_0_data_9 <= io_in_c_bypass_4_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_0_is_stationary_9 <= io_in_c_bypass_4_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_1_data_9 <= io_in_c_bypass_4_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_1_is_stationary_9 <= io_in_c_bypass_4_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_2_data_9 <= io_in_c_bypass_4_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_2_is_stationary_9 <= io_in_c_bypass_4_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_3_data_9 <= io_in_c_bypass_4_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_3_is_stationary_9 <= io_in_c_bypass_4_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_0_data_9 <= io_in_c_bypass_5_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_0_is_stationary_9 <= io_in_c_bypass_5_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_1_data_9 <= io_in_c_bypass_5_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_1_is_stationary_9 <= io_in_c_bypass_5_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_2_data_9 <= io_in_c_bypass_5_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_2_is_stationary_9 <= io_in_c_bypass_5_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_3_data_9 <= io_in_c_bypass_5_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_3_is_stationary_9 <= io_in_c_bypass_5_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_0_data_9 <= io_in_c_bypass_6_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_0_is_stationary_9 <= io_in_c_bypass_6_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_1_data_9 <= io_in_c_bypass_6_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_1_is_stationary_9 <= io_in_c_bypass_6_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_2_data_9 <= io_in_c_bypass_6_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_2_is_stationary_9 <= io_in_c_bypass_6_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_3_data_9 <= io_in_c_bypass_6_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_3_is_stationary_9 <= io_in_c_bypass_6_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_0_data_9 <= io_in_c_bypass_7_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_0_is_stationary_9 <= io_in_c_bypass_7_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_1_data_9 <= io_in_c_bypass_7_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_1_is_stationary_9 <= io_in_c_bypass_7_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_2_data_9 <= io_in_c_bypass_7_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_2_is_stationary_9 <= io_in_c_bypass_7_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_3_data_9 <= io_in_c_bypass_7_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_3_is_stationary_9 <= io_in_c_bypass_7_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_0_data_9 <= io_in_c_bypass_8_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_0_is_stationary_9 <= io_in_c_bypass_8_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_1_data_9 <= io_in_c_bypass_8_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_1_is_stationary_9 <= io_in_c_bypass_8_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_2_data_9 <= io_in_c_bypass_8_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_2_is_stationary_9 <= io_in_c_bypass_8_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_3_data_9 <= io_in_c_bypass_8_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_3_is_stationary_9 <= io_in_c_bypass_8_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_0_data_9 <= io_in_c_bypass_9_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_0_is_stationary_9 <= io_in_c_bypass_9_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_1_data_9 <= io_in_c_bypass_9_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_1_is_stationary_9 <= io_in_c_bypass_9_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_2_data_9 <= io_in_c_bypass_9_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_2_is_stationary_9 <= io_in_c_bypass_9_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_3_data_9 <= io_in_c_bypass_9_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_3_is_stationary_9 <= io_in_c_bypass_9_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_0_data_9 <= io_in_c_bypass_10_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_0_is_stationary_9 <= io_in_c_bypass_10_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_1_data_9 <= io_in_c_bypass_10_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_1_is_stationary_9 <= io_in_c_bypass_10_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_2_data_9 <= io_in_c_bypass_10_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_2_is_stationary_9 <= io_in_c_bypass_10_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_3_data_9 <= io_in_c_bypass_10_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_3_is_stationary_9 <= io_in_c_bypass_10_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_0_data_9 <= io_in_c_bypass_11_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_0_is_stationary_9 <= io_in_c_bypass_11_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_1_data_9 <= io_in_c_bypass_11_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_1_is_stationary_9 <= io_in_c_bypass_11_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_2_data_9 <= io_in_c_bypass_11_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_2_is_stationary_9 <= io_in_c_bypass_11_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_3_data_9 <= io_in_c_bypass_11_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_3_is_stationary_9 <= io_in_c_bypass_11_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_0_data_9 <= io_in_c_bypass_12_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_0_is_stationary_9 <= io_in_c_bypass_12_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_1_data_9 <= io_in_c_bypass_12_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_1_is_stationary_9 <= io_in_c_bypass_12_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_2_data_9 <= io_in_c_bypass_12_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_2_is_stationary_9 <= io_in_c_bypass_12_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_3_data_9 <= io_in_c_bypass_12_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_3_is_stationary_9 <= io_in_c_bypass_12_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_0_data_9 <= io_in_c_bypass_13_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_0_is_stationary_9 <= io_in_c_bypass_13_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_1_data_9 <= io_in_c_bypass_13_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_1_is_stationary_9 <= io_in_c_bypass_13_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_2_data_9 <= io_in_c_bypass_13_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_2_is_stationary_9 <= io_in_c_bypass_13_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_3_data_9 <= io_in_c_bypass_13_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_3_is_stationary_9 <= io_in_c_bypass_13_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_0_data_9 <= io_in_c_bypass_14_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_0_is_stationary_9 <= io_in_c_bypass_14_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_1_data_9 <= io_in_c_bypass_14_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_1_is_stationary_9 <= io_in_c_bypass_14_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_2_data_9 <= io_in_c_bypass_14_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_2_is_stationary_9 <= io_in_c_bypass_14_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_3_data_9 <= io_in_c_bypass_14_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_3_is_stationary_9 <= io_in_c_bypass_14_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_0_data_9 <= io_in_c_bypass_15_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_0_is_stationary_9 <= io_in_c_bypass_15_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_1_data_9 <= io_in_c_bypass_15_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_1_is_stationary_9 <= io_in_c_bypass_15_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_2_data_9 <= io_in_c_bypass_15_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_2_is_stationary_9 <= io_in_c_bypass_15_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_3_data_9 <= io_in_c_bypass_15_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_3_is_stationary_9 <= io_in_c_bypass_15_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_0_data_9 <= io_in_c_bypass_16_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_0_is_stationary_9 <= io_in_c_bypass_16_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_1_data_9 <= io_in_c_bypass_16_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_1_is_stationary_9 <= io_in_c_bypass_16_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_2_data_9 <= io_in_c_bypass_16_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_2_is_stationary_9 <= io_in_c_bypass_16_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_3_data_9 <= io_in_c_bypass_16_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_3_is_stationary_9 <= io_in_c_bypass_16_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_0_data_9 <= io_in_c_bypass_17_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_0_is_stationary_9 <= io_in_c_bypass_17_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_1_data_9 <= io_in_c_bypass_17_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_1_is_stationary_9 <= io_in_c_bypass_17_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_2_data_9 <= io_in_c_bypass_17_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_2_is_stationary_9 <= io_in_c_bypass_17_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_3_data_9 <= io_in_c_bypass_17_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_3_is_stationary_9 <= io_in_c_bypass_17_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_0_data_9 <= io_in_c_bypass_18_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_0_is_stationary_9 <= io_in_c_bypass_18_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_1_data_9 <= io_in_c_bypass_18_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_1_is_stationary_9 <= io_in_c_bypass_18_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_2_data_9 <= io_in_c_bypass_18_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_2_is_stationary_9 <= io_in_c_bypass_18_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_3_data_9 <= io_in_c_bypass_18_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_3_is_stationary_9 <= io_in_c_bypass_18_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_0_data_9 <= io_in_c_bypass_19_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_0_is_stationary_9 <= io_in_c_bypass_19_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_1_data_9 <= io_in_c_bypass_19_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_1_is_stationary_9 <= io_in_c_bypass_19_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_2_data_9 <= io_in_c_bypass_19_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_2_is_stationary_9 <= io_in_c_bypass_19_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_3_data_9 <= io_in_c_bypass_19_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_3_is_stationary_9 <= io_in_c_bypass_19_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_0_data_9 <= io_in_c_bypass_20_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_0_is_stationary_9 <= io_in_c_bypass_20_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_1_data_9 <= io_in_c_bypass_20_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_1_is_stationary_9 <= io_in_c_bypass_20_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_2_data_9 <= io_in_c_bypass_20_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_2_is_stationary_9 <= io_in_c_bypass_20_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_3_data_9 <= io_in_c_bypass_20_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_3_is_stationary_9 <= io_in_c_bypass_20_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_0_data_9 <= io_in_c_bypass_21_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_0_is_stationary_9 <= io_in_c_bypass_21_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_1_data_9 <= io_in_c_bypass_21_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_1_is_stationary_9 <= io_in_c_bypass_21_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_2_data_9 <= io_in_c_bypass_21_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_2_is_stationary_9 <= io_in_c_bypass_21_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_3_data_9 <= io_in_c_bypass_21_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_3_is_stationary_9 <= io_in_c_bypass_21_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_0_data_9 <= io_in_c_bypass_22_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_0_is_stationary_9 <= io_in_c_bypass_22_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_1_data_9 <= io_in_c_bypass_22_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_1_is_stationary_9 <= io_in_c_bypass_22_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_2_data_9 <= io_in_c_bypass_22_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_2_is_stationary_9 <= io_in_c_bypass_22_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_3_data_9 <= io_in_c_bypass_22_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_3_is_stationary_9 <= io_in_c_bypass_22_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_0_data_9 <= io_in_c_bypass_23_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_0_is_stationary_9 <= io_in_c_bypass_23_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_1_data_9 <= io_in_c_bypass_23_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_1_is_stationary_9 <= io_in_c_bypass_23_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_2_data_9 <= io_in_c_bypass_23_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_2_is_stationary_9 <= io_in_c_bypass_23_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_3_data_9 <= io_in_c_bypass_23_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_3_is_stationary_9 <= io_in_c_bypass_23_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_0_data_9 <= io_in_c_bypass_24_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_0_is_stationary_9 <= io_in_c_bypass_24_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_1_data_9 <= io_in_c_bypass_24_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_1_is_stationary_9 <= io_in_c_bypass_24_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_2_data_9 <= io_in_c_bypass_24_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_2_is_stationary_9 <= io_in_c_bypass_24_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_3_data_9 <= io_in_c_bypass_24_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_3_is_stationary_9 <= io_in_c_bypass_24_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_0_data_9 <= io_in_c_bypass_25_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_0_is_stationary_9 <= io_in_c_bypass_25_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_1_data_9 <= io_in_c_bypass_25_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_1_is_stationary_9 <= io_in_c_bypass_25_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_2_data_9 <= io_in_c_bypass_25_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_2_is_stationary_9 <= io_in_c_bypass_25_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_3_data_9 <= io_in_c_bypass_25_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_3_is_stationary_9 <= io_in_c_bypass_25_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_0_data_9 <= io_in_c_bypass_26_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_0_is_stationary_9 <= io_in_c_bypass_26_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_1_data_9 <= io_in_c_bypass_26_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_1_is_stationary_9 <= io_in_c_bypass_26_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_2_data_9 <= io_in_c_bypass_26_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_2_is_stationary_9 <= io_in_c_bypass_26_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_3_data_9 <= io_in_c_bypass_26_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_3_is_stationary_9 <= io_in_c_bypass_26_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_0_data_9 <= io_in_c_bypass_27_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_0_is_stationary_9 <= io_in_c_bypass_27_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_1_data_9 <= io_in_c_bypass_27_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_1_is_stationary_9 <= io_in_c_bypass_27_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_2_data_9 <= io_in_c_bypass_27_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_2_is_stationary_9 <= io_in_c_bypass_27_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_3_data_9 <= io_in_c_bypass_27_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_3_is_stationary_9 <= io_in_c_bypass_27_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_0_data_9 <= io_in_c_bypass_28_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_0_is_stationary_9 <= io_in_c_bypass_28_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_1_data_9 <= io_in_c_bypass_28_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_1_is_stationary_9 <= io_in_c_bypass_28_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_2_data_9 <= io_in_c_bypass_28_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_2_is_stationary_9 <= io_in_c_bypass_28_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_3_data_9 <= io_in_c_bypass_28_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_3_is_stationary_9 <= io_in_c_bypass_28_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_0_data_9 <= io_in_c_bypass_29_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_0_is_stationary_9 <= io_in_c_bypass_29_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_1_data_9 <= io_in_c_bypass_29_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_1_is_stationary_9 <= io_in_c_bypass_29_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_2_data_9 <= io_in_c_bypass_29_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_2_is_stationary_9 <= io_in_c_bypass_29_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_3_data_9 <= io_in_c_bypass_29_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_3_is_stationary_9 <= io_in_c_bypass_29_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_0_data_9 <= io_in_c_bypass_30_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_0_is_stationary_9 <= io_in_c_bypass_30_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_1_data_9 <= io_in_c_bypass_30_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_1_is_stationary_9 <= io_in_c_bypass_30_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_2_data_9 <= io_in_c_bypass_30_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_2_is_stationary_9 <= io_in_c_bypass_30_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_3_data_9 <= io_in_c_bypass_30_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_3_is_stationary_9 <= io_in_c_bypass_30_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_0_data_9 <= io_in_c_bypass_31_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_0_is_stationary_9 <= io_in_c_bypass_31_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_1_data_9 <= io_in_c_bypass_31_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_1_is_stationary_9 <= io_in_c_bypass_31_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_2_data_9 <= io_in_c_bypass_31_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_2_is_stationary_9 <= io_in_c_bypass_31_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_3_data_9 <= io_in_c_bypass_31_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_3_is_stationary_9 <= io_in_c_bypass_31_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_0_data_10 <= io_in_c_bypass_0_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_0_is_stationary_10 <= io_in_c_bypass_0_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_1_data_10 <= io_in_c_bypass_0_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_1_is_stationary_10 <= io_in_c_bypass_0_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_2_data_10 <= io_in_c_bypass_0_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_2_is_stationary_10 <= io_in_c_bypass_0_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_3_data_10 <= io_in_c_bypass_0_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_3_is_stationary_10 <= io_in_c_bypass_0_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_0_data_10 <= io_in_c_bypass_1_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_0_is_stationary_10 <= io_in_c_bypass_1_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_1_data_10 <= io_in_c_bypass_1_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_1_is_stationary_10 <= io_in_c_bypass_1_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_2_data_10 <= io_in_c_bypass_1_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_2_is_stationary_10 <= io_in_c_bypass_1_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_3_data_10 <= io_in_c_bypass_1_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_3_is_stationary_10 <= io_in_c_bypass_1_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_0_data_10 <= io_in_c_bypass_2_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_0_is_stationary_10 <= io_in_c_bypass_2_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_1_data_10 <= io_in_c_bypass_2_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_1_is_stationary_10 <= io_in_c_bypass_2_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_2_data_10 <= io_in_c_bypass_2_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_2_is_stationary_10 <= io_in_c_bypass_2_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_3_data_10 <= io_in_c_bypass_2_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_3_is_stationary_10 <= io_in_c_bypass_2_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_0_data_10 <= io_in_c_bypass_3_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_0_is_stationary_10 <= io_in_c_bypass_3_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_1_data_10 <= io_in_c_bypass_3_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_1_is_stationary_10 <= io_in_c_bypass_3_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_2_data_10 <= io_in_c_bypass_3_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_2_is_stationary_10 <= io_in_c_bypass_3_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_3_data_10 <= io_in_c_bypass_3_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_3_is_stationary_10 <= io_in_c_bypass_3_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_0_data_10 <= io_in_c_bypass_4_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_0_is_stationary_10 <= io_in_c_bypass_4_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_1_data_10 <= io_in_c_bypass_4_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_1_is_stationary_10 <= io_in_c_bypass_4_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_2_data_10 <= io_in_c_bypass_4_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_2_is_stationary_10 <= io_in_c_bypass_4_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_3_data_10 <= io_in_c_bypass_4_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_3_is_stationary_10 <= io_in_c_bypass_4_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_0_data_10 <= io_in_c_bypass_5_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_0_is_stationary_10 <= io_in_c_bypass_5_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_1_data_10 <= io_in_c_bypass_5_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_1_is_stationary_10 <= io_in_c_bypass_5_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_2_data_10 <= io_in_c_bypass_5_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_2_is_stationary_10 <= io_in_c_bypass_5_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_3_data_10 <= io_in_c_bypass_5_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_3_is_stationary_10 <= io_in_c_bypass_5_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_0_data_10 <= io_in_c_bypass_6_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_0_is_stationary_10 <= io_in_c_bypass_6_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_1_data_10 <= io_in_c_bypass_6_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_1_is_stationary_10 <= io_in_c_bypass_6_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_2_data_10 <= io_in_c_bypass_6_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_2_is_stationary_10 <= io_in_c_bypass_6_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_3_data_10 <= io_in_c_bypass_6_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_3_is_stationary_10 <= io_in_c_bypass_6_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_0_data_10 <= io_in_c_bypass_7_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_0_is_stationary_10 <= io_in_c_bypass_7_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_1_data_10 <= io_in_c_bypass_7_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_1_is_stationary_10 <= io_in_c_bypass_7_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_2_data_10 <= io_in_c_bypass_7_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_2_is_stationary_10 <= io_in_c_bypass_7_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_3_data_10 <= io_in_c_bypass_7_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_3_is_stationary_10 <= io_in_c_bypass_7_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_0_data_10 <= io_in_c_bypass_8_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_0_is_stationary_10 <= io_in_c_bypass_8_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_1_data_10 <= io_in_c_bypass_8_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_1_is_stationary_10 <= io_in_c_bypass_8_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_2_data_10 <= io_in_c_bypass_8_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_2_is_stationary_10 <= io_in_c_bypass_8_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_3_data_10 <= io_in_c_bypass_8_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_3_is_stationary_10 <= io_in_c_bypass_8_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_0_data_10 <= io_in_c_bypass_9_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_0_is_stationary_10 <= io_in_c_bypass_9_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_1_data_10 <= io_in_c_bypass_9_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_1_is_stationary_10 <= io_in_c_bypass_9_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_2_data_10 <= io_in_c_bypass_9_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_2_is_stationary_10 <= io_in_c_bypass_9_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_3_data_10 <= io_in_c_bypass_9_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_3_is_stationary_10 <= io_in_c_bypass_9_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_0_data_10 <= io_in_c_bypass_10_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_0_is_stationary_10 <= io_in_c_bypass_10_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_1_data_10 <= io_in_c_bypass_10_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_1_is_stationary_10 <= io_in_c_bypass_10_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_2_data_10 <= io_in_c_bypass_10_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_2_is_stationary_10 <= io_in_c_bypass_10_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_3_data_10 <= io_in_c_bypass_10_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_3_is_stationary_10 <= io_in_c_bypass_10_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_0_data_10 <= io_in_c_bypass_11_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_0_is_stationary_10 <= io_in_c_bypass_11_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_1_data_10 <= io_in_c_bypass_11_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_1_is_stationary_10 <= io_in_c_bypass_11_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_2_data_10 <= io_in_c_bypass_11_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_2_is_stationary_10 <= io_in_c_bypass_11_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_3_data_10 <= io_in_c_bypass_11_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_3_is_stationary_10 <= io_in_c_bypass_11_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_0_data_10 <= io_in_c_bypass_12_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_0_is_stationary_10 <= io_in_c_bypass_12_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_1_data_10 <= io_in_c_bypass_12_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_1_is_stationary_10 <= io_in_c_bypass_12_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_2_data_10 <= io_in_c_bypass_12_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_2_is_stationary_10 <= io_in_c_bypass_12_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_3_data_10 <= io_in_c_bypass_12_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_3_is_stationary_10 <= io_in_c_bypass_12_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_0_data_10 <= io_in_c_bypass_13_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_0_is_stationary_10 <= io_in_c_bypass_13_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_1_data_10 <= io_in_c_bypass_13_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_1_is_stationary_10 <= io_in_c_bypass_13_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_2_data_10 <= io_in_c_bypass_13_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_2_is_stationary_10 <= io_in_c_bypass_13_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_3_data_10 <= io_in_c_bypass_13_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_3_is_stationary_10 <= io_in_c_bypass_13_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_0_data_10 <= io_in_c_bypass_14_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_0_is_stationary_10 <= io_in_c_bypass_14_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_1_data_10 <= io_in_c_bypass_14_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_1_is_stationary_10 <= io_in_c_bypass_14_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_2_data_10 <= io_in_c_bypass_14_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_2_is_stationary_10 <= io_in_c_bypass_14_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_3_data_10 <= io_in_c_bypass_14_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_3_is_stationary_10 <= io_in_c_bypass_14_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_0_data_10 <= io_in_c_bypass_15_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_0_is_stationary_10 <= io_in_c_bypass_15_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_1_data_10 <= io_in_c_bypass_15_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_1_is_stationary_10 <= io_in_c_bypass_15_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_2_data_10 <= io_in_c_bypass_15_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_2_is_stationary_10 <= io_in_c_bypass_15_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_3_data_10 <= io_in_c_bypass_15_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_3_is_stationary_10 <= io_in_c_bypass_15_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_0_data_10 <= io_in_c_bypass_16_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_0_is_stationary_10 <= io_in_c_bypass_16_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_1_data_10 <= io_in_c_bypass_16_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_1_is_stationary_10 <= io_in_c_bypass_16_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_2_data_10 <= io_in_c_bypass_16_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_2_is_stationary_10 <= io_in_c_bypass_16_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_3_data_10 <= io_in_c_bypass_16_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_3_is_stationary_10 <= io_in_c_bypass_16_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_0_data_10 <= io_in_c_bypass_17_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_0_is_stationary_10 <= io_in_c_bypass_17_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_1_data_10 <= io_in_c_bypass_17_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_1_is_stationary_10 <= io_in_c_bypass_17_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_2_data_10 <= io_in_c_bypass_17_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_2_is_stationary_10 <= io_in_c_bypass_17_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_3_data_10 <= io_in_c_bypass_17_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_3_is_stationary_10 <= io_in_c_bypass_17_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_0_data_10 <= io_in_c_bypass_18_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_0_is_stationary_10 <= io_in_c_bypass_18_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_1_data_10 <= io_in_c_bypass_18_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_1_is_stationary_10 <= io_in_c_bypass_18_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_2_data_10 <= io_in_c_bypass_18_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_2_is_stationary_10 <= io_in_c_bypass_18_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_3_data_10 <= io_in_c_bypass_18_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_3_is_stationary_10 <= io_in_c_bypass_18_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_0_data_10 <= io_in_c_bypass_19_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_0_is_stationary_10 <= io_in_c_bypass_19_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_1_data_10 <= io_in_c_bypass_19_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_1_is_stationary_10 <= io_in_c_bypass_19_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_2_data_10 <= io_in_c_bypass_19_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_2_is_stationary_10 <= io_in_c_bypass_19_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_3_data_10 <= io_in_c_bypass_19_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_3_is_stationary_10 <= io_in_c_bypass_19_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_0_data_10 <= io_in_c_bypass_20_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_0_is_stationary_10 <= io_in_c_bypass_20_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_1_data_10 <= io_in_c_bypass_20_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_1_is_stationary_10 <= io_in_c_bypass_20_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_2_data_10 <= io_in_c_bypass_20_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_2_is_stationary_10 <= io_in_c_bypass_20_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_3_data_10 <= io_in_c_bypass_20_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_3_is_stationary_10 <= io_in_c_bypass_20_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_0_data_10 <= io_in_c_bypass_21_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_0_is_stationary_10 <= io_in_c_bypass_21_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_1_data_10 <= io_in_c_bypass_21_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_1_is_stationary_10 <= io_in_c_bypass_21_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_2_data_10 <= io_in_c_bypass_21_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_2_is_stationary_10 <= io_in_c_bypass_21_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_3_data_10 <= io_in_c_bypass_21_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_3_is_stationary_10 <= io_in_c_bypass_21_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_0_data_10 <= io_in_c_bypass_22_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_0_is_stationary_10 <= io_in_c_bypass_22_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_1_data_10 <= io_in_c_bypass_22_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_1_is_stationary_10 <= io_in_c_bypass_22_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_2_data_10 <= io_in_c_bypass_22_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_2_is_stationary_10 <= io_in_c_bypass_22_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_3_data_10 <= io_in_c_bypass_22_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_3_is_stationary_10 <= io_in_c_bypass_22_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_0_data_10 <= io_in_c_bypass_23_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_0_is_stationary_10 <= io_in_c_bypass_23_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_1_data_10 <= io_in_c_bypass_23_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_1_is_stationary_10 <= io_in_c_bypass_23_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_2_data_10 <= io_in_c_bypass_23_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_2_is_stationary_10 <= io_in_c_bypass_23_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_3_data_10 <= io_in_c_bypass_23_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_3_is_stationary_10 <= io_in_c_bypass_23_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_0_data_10 <= io_in_c_bypass_24_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_0_is_stationary_10 <= io_in_c_bypass_24_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_1_data_10 <= io_in_c_bypass_24_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_1_is_stationary_10 <= io_in_c_bypass_24_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_2_data_10 <= io_in_c_bypass_24_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_2_is_stationary_10 <= io_in_c_bypass_24_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_3_data_10 <= io_in_c_bypass_24_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_3_is_stationary_10 <= io_in_c_bypass_24_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_0_data_10 <= io_in_c_bypass_25_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_0_is_stationary_10 <= io_in_c_bypass_25_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_1_data_10 <= io_in_c_bypass_25_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_1_is_stationary_10 <= io_in_c_bypass_25_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_2_data_10 <= io_in_c_bypass_25_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_2_is_stationary_10 <= io_in_c_bypass_25_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_3_data_10 <= io_in_c_bypass_25_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_3_is_stationary_10 <= io_in_c_bypass_25_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_0_data_10 <= io_in_c_bypass_26_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_0_is_stationary_10 <= io_in_c_bypass_26_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_1_data_10 <= io_in_c_bypass_26_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_1_is_stationary_10 <= io_in_c_bypass_26_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_2_data_10 <= io_in_c_bypass_26_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_2_is_stationary_10 <= io_in_c_bypass_26_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_3_data_10 <= io_in_c_bypass_26_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_3_is_stationary_10 <= io_in_c_bypass_26_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_0_data_10 <= io_in_c_bypass_27_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_0_is_stationary_10 <= io_in_c_bypass_27_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_1_data_10 <= io_in_c_bypass_27_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_1_is_stationary_10 <= io_in_c_bypass_27_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_2_data_10 <= io_in_c_bypass_27_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_2_is_stationary_10 <= io_in_c_bypass_27_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_3_data_10 <= io_in_c_bypass_27_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_3_is_stationary_10 <= io_in_c_bypass_27_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_0_data_10 <= io_in_c_bypass_28_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_0_is_stationary_10 <= io_in_c_bypass_28_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_1_data_10 <= io_in_c_bypass_28_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_1_is_stationary_10 <= io_in_c_bypass_28_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_2_data_10 <= io_in_c_bypass_28_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_2_is_stationary_10 <= io_in_c_bypass_28_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_3_data_10 <= io_in_c_bypass_28_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_3_is_stationary_10 <= io_in_c_bypass_28_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_0_data_10 <= io_in_c_bypass_29_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_0_is_stationary_10 <= io_in_c_bypass_29_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_1_data_10 <= io_in_c_bypass_29_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_1_is_stationary_10 <= io_in_c_bypass_29_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_2_data_10 <= io_in_c_bypass_29_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_2_is_stationary_10 <= io_in_c_bypass_29_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_3_data_10 <= io_in_c_bypass_29_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_3_is_stationary_10 <= io_in_c_bypass_29_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_0_data_10 <= io_in_c_bypass_30_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_0_is_stationary_10 <= io_in_c_bypass_30_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_1_data_10 <= io_in_c_bypass_30_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_1_is_stationary_10 <= io_in_c_bypass_30_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_2_data_10 <= io_in_c_bypass_30_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_2_is_stationary_10 <= io_in_c_bypass_30_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_3_data_10 <= io_in_c_bypass_30_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_3_is_stationary_10 <= io_in_c_bypass_30_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_0_data_10 <= io_in_c_bypass_31_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_0_is_stationary_10 <= io_in_c_bypass_31_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_1_data_10 <= io_in_c_bypass_31_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_1_is_stationary_10 <= io_in_c_bypass_31_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_2_data_10 <= io_in_c_bypass_31_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_2_is_stationary_10 <= io_in_c_bypass_31_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_3_data_10 <= io_in_c_bypass_31_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_3_is_stationary_10 <= io_in_c_bypass_31_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_0_data_11 <= io_in_c_bypass_0_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_0_is_stationary_11 <= io_in_c_bypass_0_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_1_data_11 <= io_in_c_bypass_0_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_1_is_stationary_11 <= io_in_c_bypass_0_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_2_data_11 <= io_in_c_bypass_0_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_2_is_stationary_11 <= io_in_c_bypass_0_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_3_data_11 <= io_in_c_bypass_0_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_3_is_stationary_11 <= io_in_c_bypass_0_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_0_data_11 <= io_in_c_bypass_1_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_0_is_stationary_11 <= io_in_c_bypass_1_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_1_data_11 <= io_in_c_bypass_1_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_1_is_stationary_11 <= io_in_c_bypass_1_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_2_data_11 <= io_in_c_bypass_1_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_2_is_stationary_11 <= io_in_c_bypass_1_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_3_data_11 <= io_in_c_bypass_1_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_3_is_stationary_11 <= io_in_c_bypass_1_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_0_data_11 <= io_in_c_bypass_2_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_0_is_stationary_11 <= io_in_c_bypass_2_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_1_data_11 <= io_in_c_bypass_2_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_1_is_stationary_11 <= io_in_c_bypass_2_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_2_data_11 <= io_in_c_bypass_2_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_2_is_stationary_11 <= io_in_c_bypass_2_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_3_data_11 <= io_in_c_bypass_2_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_3_is_stationary_11 <= io_in_c_bypass_2_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_0_data_11 <= io_in_c_bypass_3_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_0_is_stationary_11 <= io_in_c_bypass_3_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_1_data_11 <= io_in_c_bypass_3_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_1_is_stationary_11 <= io_in_c_bypass_3_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_2_data_11 <= io_in_c_bypass_3_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_2_is_stationary_11 <= io_in_c_bypass_3_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_3_data_11 <= io_in_c_bypass_3_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_3_is_stationary_11 <= io_in_c_bypass_3_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_0_data_11 <= io_in_c_bypass_4_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_0_is_stationary_11 <= io_in_c_bypass_4_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_1_data_11 <= io_in_c_bypass_4_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_1_is_stationary_11 <= io_in_c_bypass_4_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_2_data_11 <= io_in_c_bypass_4_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_2_is_stationary_11 <= io_in_c_bypass_4_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_3_data_11 <= io_in_c_bypass_4_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_3_is_stationary_11 <= io_in_c_bypass_4_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_0_data_11 <= io_in_c_bypass_5_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_0_is_stationary_11 <= io_in_c_bypass_5_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_1_data_11 <= io_in_c_bypass_5_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_1_is_stationary_11 <= io_in_c_bypass_5_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_2_data_11 <= io_in_c_bypass_5_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_2_is_stationary_11 <= io_in_c_bypass_5_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_3_data_11 <= io_in_c_bypass_5_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_3_is_stationary_11 <= io_in_c_bypass_5_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_0_data_11 <= io_in_c_bypass_6_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_0_is_stationary_11 <= io_in_c_bypass_6_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_1_data_11 <= io_in_c_bypass_6_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_1_is_stationary_11 <= io_in_c_bypass_6_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_2_data_11 <= io_in_c_bypass_6_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_2_is_stationary_11 <= io_in_c_bypass_6_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_3_data_11 <= io_in_c_bypass_6_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_3_is_stationary_11 <= io_in_c_bypass_6_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_0_data_11 <= io_in_c_bypass_7_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_0_is_stationary_11 <= io_in_c_bypass_7_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_1_data_11 <= io_in_c_bypass_7_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_1_is_stationary_11 <= io_in_c_bypass_7_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_2_data_11 <= io_in_c_bypass_7_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_2_is_stationary_11 <= io_in_c_bypass_7_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_3_data_11 <= io_in_c_bypass_7_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_3_is_stationary_11 <= io_in_c_bypass_7_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_0_data_11 <= io_in_c_bypass_8_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_0_is_stationary_11 <= io_in_c_bypass_8_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_1_data_11 <= io_in_c_bypass_8_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_1_is_stationary_11 <= io_in_c_bypass_8_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_2_data_11 <= io_in_c_bypass_8_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_2_is_stationary_11 <= io_in_c_bypass_8_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_3_data_11 <= io_in_c_bypass_8_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_3_is_stationary_11 <= io_in_c_bypass_8_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_0_data_11 <= io_in_c_bypass_9_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_0_is_stationary_11 <= io_in_c_bypass_9_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_1_data_11 <= io_in_c_bypass_9_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_1_is_stationary_11 <= io_in_c_bypass_9_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_2_data_11 <= io_in_c_bypass_9_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_2_is_stationary_11 <= io_in_c_bypass_9_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_3_data_11 <= io_in_c_bypass_9_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_3_is_stationary_11 <= io_in_c_bypass_9_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_0_data_11 <= io_in_c_bypass_10_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_0_is_stationary_11 <= io_in_c_bypass_10_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_1_data_11 <= io_in_c_bypass_10_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_1_is_stationary_11 <= io_in_c_bypass_10_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_2_data_11 <= io_in_c_bypass_10_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_2_is_stationary_11 <= io_in_c_bypass_10_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_3_data_11 <= io_in_c_bypass_10_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_3_is_stationary_11 <= io_in_c_bypass_10_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_0_data_11 <= io_in_c_bypass_11_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_0_is_stationary_11 <= io_in_c_bypass_11_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_1_data_11 <= io_in_c_bypass_11_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_1_is_stationary_11 <= io_in_c_bypass_11_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_2_data_11 <= io_in_c_bypass_11_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_2_is_stationary_11 <= io_in_c_bypass_11_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_3_data_11 <= io_in_c_bypass_11_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_3_is_stationary_11 <= io_in_c_bypass_11_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_0_data_11 <= io_in_c_bypass_12_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_0_is_stationary_11 <= io_in_c_bypass_12_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_1_data_11 <= io_in_c_bypass_12_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_1_is_stationary_11 <= io_in_c_bypass_12_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_2_data_11 <= io_in_c_bypass_12_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_2_is_stationary_11 <= io_in_c_bypass_12_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_3_data_11 <= io_in_c_bypass_12_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_3_is_stationary_11 <= io_in_c_bypass_12_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_0_data_11 <= io_in_c_bypass_13_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_0_is_stationary_11 <= io_in_c_bypass_13_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_1_data_11 <= io_in_c_bypass_13_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_1_is_stationary_11 <= io_in_c_bypass_13_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_2_data_11 <= io_in_c_bypass_13_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_2_is_stationary_11 <= io_in_c_bypass_13_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_3_data_11 <= io_in_c_bypass_13_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_3_is_stationary_11 <= io_in_c_bypass_13_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_0_data_11 <= io_in_c_bypass_14_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_0_is_stationary_11 <= io_in_c_bypass_14_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_1_data_11 <= io_in_c_bypass_14_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_1_is_stationary_11 <= io_in_c_bypass_14_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_2_data_11 <= io_in_c_bypass_14_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_2_is_stationary_11 <= io_in_c_bypass_14_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_3_data_11 <= io_in_c_bypass_14_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_3_is_stationary_11 <= io_in_c_bypass_14_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_0_data_11 <= io_in_c_bypass_15_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_0_is_stationary_11 <= io_in_c_bypass_15_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_1_data_11 <= io_in_c_bypass_15_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_1_is_stationary_11 <= io_in_c_bypass_15_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_2_data_11 <= io_in_c_bypass_15_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_2_is_stationary_11 <= io_in_c_bypass_15_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_3_data_11 <= io_in_c_bypass_15_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_3_is_stationary_11 <= io_in_c_bypass_15_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_0_data_11 <= io_in_c_bypass_16_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_0_is_stationary_11 <= io_in_c_bypass_16_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_1_data_11 <= io_in_c_bypass_16_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_1_is_stationary_11 <= io_in_c_bypass_16_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_2_data_11 <= io_in_c_bypass_16_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_2_is_stationary_11 <= io_in_c_bypass_16_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_3_data_11 <= io_in_c_bypass_16_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_3_is_stationary_11 <= io_in_c_bypass_16_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_0_data_11 <= io_in_c_bypass_17_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_0_is_stationary_11 <= io_in_c_bypass_17_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_1_data_11 <= io_in_c_bypass_17_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_1_is_stationary_11 <= io_in_c_bypass_17_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_2_data_11 <= io_in_c_bypass_17_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_2_is_stationary_11 <= io_in_c_bypass_17_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_3_data_11 <= io_in_c_bypass_17_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_3_is_stationary_11 <= io_in_c_bypass_17_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_0_data_11 <= io_in_c_bypass_18_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_0_is_stationary_11 <= io_in_c_bypass_18_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_1_data_11 <= io_in_c_bypass_18_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_1_is_stationary_11 <= io_in_c_bypass_18_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_2_data_11 <= io_in_c_bypass_18_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_2_is_stationary_11 <= io_in_c_bypass_18_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_3_data_11 <= io_in_c_bypass_18_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_3_is_stationary_11 <= io_in_c_bypass_18_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_0_data_11 <= io_in_c_bypass_19_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_0_is_stationary_11 <= io_in_c_bypass_19_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_1_data_11 <= io_in_c_bypass_19_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_1_is_stationary_11 <= io_in_c_bypass_19_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_2_data_11 <= io_in_c_bypass_19_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_2_is_stationary_11 <= io_in_c_bypass_19_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_3_data_11 <= io_in_c_bypass_19_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_3_is_stationary_11 <= io_in_c_bypass_19_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_0_data_11 <= io_in_c_bypass_20_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_0_is_stationary_11 <= io_in_c_bypass_20_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_1_data_11 <= io_in_c_bypass_20_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_1_is_stationary_11 <= io_in_c_bypass_20_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_2_data_11 <= io_in_c_bypass_20_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_2_is_stationary_11 <= io_in_c_bypass_20_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_3_data_11 <= io_in_c_bypass_20_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_3_is_stationary_11 <= io_in_c_bypass_20_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_0_data_11 <= io_in_c_bypass_21_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_0_is_stationary_11 <= io_in_c_bypass_21_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_1_data_11 <= io_in_c_bypass_21_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_1_is_stationary_11 <= io_in_c_bypass_21_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_2_data_11 <= io_in_c_bypass_21_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_2_is_stationary_11 <= io_in_c_bypass_21_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_3_data_11 <= io_in_c_bypass_21_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_3_is_stationary_11 <= io_in_c_bypass_21_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_0_data_11 <= io_in_c_bypass_22_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_0_is_stationary_11 <= io_in_c_bypass_22_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_1_data_11 <= io_in_c_bypass_22_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_1_is_stationary_11 <= io_in_c_bypass_22_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_2_data_11 <= io_in_c_bypass_22_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_2_is_stationary_11 <= io_in_c_bypass_22_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_3_data_11 <= io_in_c_bypass_22_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_3_is_stationary_11 <= io_in_c_bypass_22_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_0_data_11 <= io_in_c_bypass_23_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_0_is_stationary_11 <= io_in_c_bypass_23_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_1_data_11 <= io_in_c_bypass_23_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_1_is_stationary_11 <= io_in_c_bypass_23_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_2_data_11 <= io_in_c_bypass_23_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_2_is_stationary_11 <= io_in_c_bypass_23_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_3_data_11 <= io_in_c_bypass_23_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_3_is_stationary_11 <= io_in_c_bypass_23_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_0_data_11 <= io_in_c_bypass_24_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_0_is_stationary_11 <= io_in_c_bypass_24_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_1_data_11 <= io_in_c_bypass_24_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_1_is_stationary_11 <= io_in_c_bypass_24_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_2_data_11 <= io_in_c_bypass_24_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_2_is_stationary_11 <= io_in_c_bypass_24_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_3_data_11 <= io_in_c_bypass_24_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_3_is_stationary_11 <= io_in_c_bypass_24_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_0_data_11 <= io_in_c_bypass_25_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_0_is_stationary_11 <= io_in_c_bypass_25_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_1_data_11 <= io_in_c_bypass_25_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_1_is_stationary_11 <= io_in_c_bypass_25_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_2_data_11 <= io_in_c_bypass_25_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_2_is_stationary_11 <= io_in_c_bypass_25_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_3_data_11 <= io_in_c_bypass_25_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_3_is_stationary_11 <= io_in_c_bypass_25_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_0_data_11 <= io_in_c_bypass_26_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_0_is_stationary_11 <= io_in_c_bypass_26_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_1_data_11 <= io_in_c_bypass_26_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_1_is_stationary_11 <= io_in_c_bypass_26_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_2_data_11 <= io_in_c_bypass_26_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_2_is_stationary_11 <= io_in_c_bypass_26_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_3_data_11 <= io_in_c_bypass_26_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_3_is_stationary_11 <= io_in_c_bypass_26_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_0_data_11 <= io_in_c_bypass_27_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_0_is_stationary_11 <= io_in_c_bypass_27_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_1_data_11 <= io_in_c_bypass_27_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_1_is_stationary_11 <= io_in_c_bypass_27_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_2_data_11 <= io_in_c_bypass_27_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_2_is_stationary_11 <= io_in_c_bypass_27_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_3_data_11 <= io_in_c_bypass_27_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_3_is_stationary_11 <= io_in_c_bypass_27_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_0_data_11 <= io_in_c_bypass_28_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_0_is_stationary_11 <= io_in_c_bypass_28_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_1_data_11 <= io_in_c_bypass_28_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_1_is_stationary_11 <= io_in_c_bypass_28_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_2_data_11 <= io_in_c_bypass_28_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_2_is_stationary_11 <= io_in_c_bypass_28_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_3_data_11 <= io_in_c_bypass_28_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_3_is_stationary_11 <= io_in_c_bypass_28_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_0_data_11 <= io_in_c_bypass_29_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_0_is_stationary_11 <= io_in_c_bypass_29_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_1_data_11 <= io_in_c_bypass_29_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_1_is_stationary_11 <= io_in_c_bypass_29_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_2_data_11 <= io_in_c_bypass_29_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_2_is_stationary_11 <= io_in_c_bypass_29_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_3_data_11 <= io_in_c_bypass_29_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_3_is_stationary_11 <= io_in_c_bypass_29_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_0_data_11 <= io_in_c_bypass_30_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_0_is_stationary_11 <= io_in_c_bypass_30_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_1_data_11 <= io_in_c_bypass_30_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_1_is_stationary_11 <= io_in_c_bypass_30_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_2_data_11 <= io_in_c_bypass_30_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_2_is_stationary_11 <= io_in_c_bypass_30_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_3_data_11 <= io_in_c_bypass_30_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_3_is_stationary_11 <= io_in_c_bypass_30_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_0_data_11 <= io_in_c_bypass_31_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_0_is_stationary_11 <= io_in_c_bypass_31_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_1_data_11 <= io_in_c_bypass_31_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_1_is_stationary_11 <= io_in_c_bypass_31_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_2_data_11 <= io_in_c_bypass_31_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_2_is_stationary_11 <= io_in_c_bypass_31_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_3_data_11 <= io_in_c_bypass_31_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_3_is_stationary_11 <= io_in_c_bypass_31_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_0_data_12 <= io_in_c_bypass_0_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_0_is_stationary_12 <= io_in_c_bypass_0_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_1_data_12 <= io_in_c_bypass_0_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_1_is_stationary_12 <= io_in_c_bypass_0_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_2_data_12 <= io_in_c_bypass_0_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_2_is_stationary_12 <= io_in_c_bypass_0_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_3_data_12 <= io_in_c_bypass_0_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_3_is_stationary_12 <= io_in_c_bypass_0_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_0_data_12 <= io_in_c_bypass_1_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_0_is_stationary_12 <= io_in_c_bypass_1_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_1_data_12 <= io_in_c_bypass_1_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_1_is_stationary_12 <= io_in_c_bypass_1_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_2_data_12 <= io_in_c_bypass_1_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_2_is_stationary_12 <= io_in_c_bypass_1_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_3_data_12 <= io_in_c_bypass_1_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_3_is_stationary_12 <= io_in_c_bypass_1_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_0_data_12 <= io_in_c_bypass_2_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_0_is_stationary_12 <= io_in_c_bypass_2_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_1_data_12 <= io_in_c_bypass_2_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_1_is_stationary_12 <= io_in_c_bypass_2_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_2_data_12 <= io_in_c_bypass_2_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_2_is_stationary_12 <= io_in_c_bypass_2_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_3_data_12 <= io_in_c_bypass_2_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_3_is_stationary_12 <= io_in_c_bypass_2_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_0_data_12 <= io_in_c_bypass_3_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_0_is_stationary_12 <= io_in_c_bypass_3_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_1_data_12 <= io_in_c_bypass_3_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_1_is_stationary_12 <= io_in_c_bypass_3_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_2_data_12 <= io_in_c_bypass_3_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_2_is_stationary_12 <= io_in_c_bypass_3_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_3_data_12 <= io_in_c_bypass_3_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_3_is_stationary_12 <= io_in_c_bypass_3_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_0_data_12 <= io_in_c_bypass_4_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_0_is_stationary_12 <= io_in_c_bypass_4_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_1_data_12 <= io_in_c_bypass_4_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_1_is_stationary_12 <= io_in_c_bypass_4_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_2_data_12 <= io_in_c_bypass_4_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_2_is_stationary_12 <= io_in_c_bypass_4_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_3_data_12 <= io_in_c_bypass_4_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_3_is_stationary_12 <= io_in_c_bypass_4_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_0_data_12 <= io_in_c_bypass_5_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_0_is_stationary_12 <= io_in_c_bypass_5_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_1_data_12 <= io_in_c_bypass_5_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_1_is_stationary_12 <= io_in_c_bypass_5_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_2_data_12 <= io_in_c_bypass_5_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_2_is_stationary_12 <= io_in_c_bypass_5_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_3_data_12 <= io_in_c_bypass_5_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_3_is_stationary_12 <= io_in_c_bypass_5_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_0_data_12 <= io_in_c_bypass_6_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_0_is_stationary_12 <= io_in_c_bypass_6_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_1_data_12 <= io_in_c_bypass_6_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_1_is_stationary_12 <= io_in_c_bypass_6_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_2_data_12 <= io_in_c_bypass_6_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_2_is_stationary_12 <= io_in_c_bypass_6_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_3_data_12 <= io_in_c_bypass_6_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_3_is_stationary_12 <= io_in_c_bypass_6_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_0_data_12 <= io_in_c_bypass_7_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_0_is_stationary_12 <= io_in_c_bypass_7_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_1_data_12 <= io_in_c_bypass_7_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_1_is_stationary_12 <= io_in_c_bypass_7_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_2_data_12 <= io_in_c_bypass_7_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_2_is_stationary_12 <= io_in_c_bypass_7_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_3_data_12 <= io_in_c_bypass_7_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_3_is_stationary_12 <= io_in_c_bypass_7_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_0_data_12 <= io_in_c_bypass_8_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_0_is_stationary_12 <= io_in_c_bypass_8_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_1_data_12 <= io_in_c_bypass_8_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_1_is_stationary_12 <= io_in_c_bypass_8_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_2_data_12 <= io_in_c_bypass_8_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_2_is_stationary_12 <= io_in_c_bypass_8_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_3_data_12 <= io_in_c_bypass_8_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_3_is_stationary_12 <= io_in_c_bypass_8_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_0_data_12 <= io_in_c_bypass_9_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_0_is_stationary_12 <= io_in_c_bypass_9_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_1_data_12 <= io_in_c_bypass_9_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_1_is_stationary_12 <= io_in_c_bypass_9_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_2_data_12 <= io_in_c_bypass_9_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_2_is_stationary_12 <= io_in_c_bypass_9_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_3_data_12 <= io_in_c_bypass_9_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_3_is_stationary_12 <= io_in_c_bypass_9_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_0_data_12 <= io_in_c_bypass_10_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_0_is_stationary_12 <= io_in_c_bypass_10_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_1_data_12 <= io_in_c_bypass_10_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_1_is_stationary_12 <= io_in_c_bypass_10_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_2_data_12 <= io_in_c_bypass_10_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_2_is_stationary_12 <= io_in_c_bypass_10_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_3_data_12 <= io_in_c_bypass_10_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_3_is_stationary_12 <= io_in_c_bypass_10_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_0_data_12 <= io_in_c_bypass_11_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_0_is_stationary_12 <= io_in_c_bypass_11_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_1_data_12 <= io_in_c_bypass_11_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_1_is_stationary_12 <= io_in_c_bypass_11_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_2_data_12 <= io_in_c_bypass_11_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_2_is_stationary_12 <= io_in_c_bypass_11_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_3_data_12 <= io_in_c_bypass_11_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_3_is_stationary_12 <= io_in_c_bypass_11_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_0_data_12 <= io_in_c_bypass_12_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_0_is_stationary_12 <= io_in_c_bypass_12_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_1_data_12 <= io_in_c_bypass_12_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_1_is_stationary_12 <= io_in_c_bypass_12_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_2_data_12 <= io_in_c_bypass_12_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_2_is_stationary_12 <= io_in_c_bypass_12_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_3_data_12 <= io_in_c_bypass_12_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_3_is_stationary_12 <= io_in_c_bypass_12_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_0_data_12 <= io_in_c_bypass_13_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_0_is_stationary_12 <= io_in_c_bypass_13_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_1_data_12 <= io_in_c_bypass_13_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_1_is_stationary_12 <= io_in_c_bypass_13_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_2_data_12 <= io_in_c_bypass_13_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_2_is_stationary_12 <= io_in_c_bypass_13_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_3_data_12 <= io_in_c_bypass_13_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_3_is_stationary_12 <= io_in_c_bypass_13_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_0_data_12 <= io_in_c_bypass_14_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_0_is_stationary_12 <= io_in_c_bypass_14_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_1_data_12 <= io_in_c_bypass_14_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_1_is_stationary_12 <= io_in_c_bypass_14_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_2_data_12 <= io_in_c_bypass_14_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_2_is_stationary_12 <= io_in_c_bypass_14_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_3_data_12 <= io_in_c_bypass_14_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_3_is_stationary_12 <= io_in_c_bypass_14_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_0_data_12 <= io_in_c_bypass_15_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_0_is_stationary_12 <= io_in_c_bypass_15_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_1_data_12 <= io_in_c_bypass_15_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_1_is_stationary_12 <= io_in_c_bypass_15_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_2_data_12 <= io_in_c_bypass_15_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_2_is_stationary_12 <= io_in_c_bypass_15_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_3_data_12 <= io_in_c_bypass_15_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_3_is_stationary_12 <= io_in_c_bypass_15_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_0_data_12 <= io_in_c_bypass_16_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_0_is_stationary_12 <= io_in_c_bypass_16_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_1_data_12 <= io_in_c_bypass_16_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_1_is_stationary_12 <= io_in_c_bypass_16_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_2_data_12 <= io_in_c_bypass_16_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_2_is_stationary_12 <= io_in_c_bypass_16_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_3_data_12 <= io_in_c_bypass_16_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_3_is_stationary_12 <= io_in_c_bypass_16_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_0_data_12 <= io_in_c_bypass_17_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_0_is_stationary_12 <= io_in_c_bypass_17_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_1_data_12 <= io_in_c_bypass_17_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_1_is_stationary_12 <= io_in_c_bypass_17_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_2_data_12 <= io_in_c_bypass_17_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_2_is_stationary_12 <= io_in_c_bypass_17_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_3_data_12 <= io_in_c_bypass_17_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_3_is_stationary_12 <= io_in_c_bypass_17_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_0_data_12 <= io_in_c_bypass_18_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_0_is_stationary_12 <= io_in_c_bypass_18_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_1_data_12 <= io_in_c_bypass_18_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_1_is_stationary_12 <= io_in_c_bypass_18_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_2_data_12 <= io_in_c_bypass_18_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_2_is_stationary_12 <= io_in_c_bypass_18_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_3_data_12 <= io_in_c_bypass_18_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_3_is_stationary_12 <= io_in_c_bypass_18_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_0_data_12 <= io_in_c_bypass_19_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_0_is_stationary_12 <= io_in_c_bypass_19_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_1_data_12 <= io_in_c_bypass_19_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_1_is_stationary_12 <= io_in_c_bypass_19_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_2_data_12 <= io_in_c_bypass_19_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_2_is_stationary_12 <= io_in_c_bypass_19_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_3_data_12 <= io_in_c_bypass_19_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_3_is_stationary_12 <= io_in_c_bypass_19_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_0_data_12 <= io_in_c_bypass_20_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_0_is_stationary_12 <= io_in_c_bypass_20_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_1_data_12 <= io_in_c_bypass_20_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_1_is_stationary_12 <= io_in_c_bypass_20_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_2_data_12 <= io_in_c_bypass_20_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_2_is_stationary_12 <= io_in_c_bypass_20_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_3_data_12 <= io_in_c_bypass_20_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_3_is_stationary_12 <= io_in_c_bypass_20_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_0_data_12 <= io_in_c_bypass_21_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_0_is_stationary_12 <= io_in_c_bypass_21_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_1_data_12 <= io_in_c_bypass_21_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_1_is_stationary_12 <= io_in_c_bypass_21_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_2_data_12 <= io_in_c_bypass_21_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_2_is_stationary_12 <= io_in_c_bypass_21_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_3_data_12 <= io_in_c_bypass_21_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_3_is_stationary_12 <= io_in_c_bypass_21_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_0_data_12 <= io_in_c_bypass_22_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_0_is_stationary_12 <= io_in_c_bypass_22_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_1_data_12 <= io_in_c_bypass_22_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_1_is_stationary_12 <= io_in_c_bypass_22_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_2_data_12 <= io_in_c_bypass_22_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_2_is_stationary_12 <= io_in_c_bypass_22_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_3_data_12 <= io_in_c_bypass_22_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_3_is_stationary_12 <= io_in_c_bypass_22_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_0_data_12 <= io_in_c_bypass_23_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_0_is_stationary_12 <= io_in_c_bypass_23_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_1_data_12 <= io_in_c_bypass_23_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_1_is_stationary_12 <= io_in_c_bypass_23_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_2_data_12 <= io_in_c_bypass_23_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_2_is_stationary_12 <= io_in_c_bypass_23_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_3_data_12 <= io_in_c_bypass_23_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_3_is_stationary_12 <= io_in_c_bypass_23_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_0_data_12 <= io_in_c_bypass_24_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_0_is_stationary_12 <= io_in_c_bypass_24_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_1_data_12 <= io_in_c_bypass_24_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_1_is_stationary_12 <= io_in_c_bypass_24_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_2_data_12 <= io_in_c_bypass_24_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_2_is_stationary_12 <= io_in_c_bypass_24_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_3_data_12 <= io_in_c_bypass_24_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_3_is_stationary_12 <= io_in_c_bypass_24_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_0_data_12 <= io_in_c_bypass_25_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_0_is_stationary_12 <= io_in_c_bypass_25_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_1_data_12 <= io_in_c_bypass_25_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_1_is_stationary_12 <= io_in_c_bypass_25_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_2_data_12 <= io_in_c_bypass_25_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_2_is_stationary_12 <= io_in_c_bypass_25_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_3_data_12 <= io_in_c_bypass_25_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_3_is_stationary_12 <= io_in_c_bypass_25_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_0_data_12 <= io_in_c_bypass_26_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_0_is_stationary_12 <= io_in_c_bypass_26_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_1_data_12 <= io_in_c_bypass_26_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_1_is_stationary_12 <= io_in_c_bypass_26_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_2_data_12 <= io_in_c_bypass_26_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_2_is_stationary_12 <= io_in_c_bypass_26_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_3_data_12 <= io_in_c_bypass_26_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_3_is_stationary_12 <= io_in_c_bypass_26_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_0_data_12 <= io_in_c_bypass_27_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_0_is_stationary_12 <= io_in_c_bypass_27_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_1_data_12 <= io_in_c_bypass_27_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_1_is_stationary_12 <= io_in_c_bypass_27_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_2_data_12 <= io_in_c_bypass_27_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_2_is_stationary_12 <= io_in_c_bypass_27_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_3_data_12 <= io_in_c_bypass_27_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_3_is_stationary_12 <= io_in_c_bypass_27_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_0_data_12 <= io_in_c_bypass_28_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_0_is_stationary_12 <= io_in_c_bypass_28_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_1_data_12 <= io_in_c_bypass_28_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_1_is_stationary_12 <= io_in_c_bypass_28_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_2_data_12 <= io_in_c_bypass_28_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_2_is_stationary_12 <= io_in_c_bypass_28_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_3_data_12 <= io_in_c_bypass_28_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_3_is_stationary_12 <= io_in_c_bypass_28_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_0_data_12 <= io_in_c_bypass_29_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_0_is_stationary_12 <= io_in_c_bypass_29_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_1_data_12 <= io_in_c_bypass_29_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_1_is_stationary_12 <= io_in_c_bypass_29_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_2_data_12 <= io_in_c_bypass_29_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_2_is_stationary_12 <= io_in_c_bypass_29_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_3_data_12 <= io_in_c_bypass_29_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_3_is_stationary_12 <= io_in_c_bypass_29_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_0_data_12 <= io_in_c_bypass_30_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_0_is_stationary_12 <= io_in_c_bypass_30_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_1_data_12 <= io_in_c_bypass_30_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_1_is_stationary_12 <= io_in_c_bypass_30_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_2_data_12 <= io_in_c_bypass_30_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_2_is_stationary_12 <= io_in_c_bypass_30_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_3_data_12 <= io_in_c_bypass_30_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_3_is_stationary_12 <= io_in_c_bypass_30_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_0_data_12 <= io_in_c_bypass_31_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_0_is_stationary_12 <= io_in_c_bypass_31_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_1_data_12 <= io_in_c_bypass_31_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_1_is_stationary_12 <= io_in_c_bypass_31_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_2_data_12 <= io_in_c_bypass_31_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_2_is_stationary_12 <= io_in_c_bypass_31_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_3_data_12 <= io_in_c_bypass_31_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_3_is_stationary_12 <= io_in_c_bypass_31_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_0_data_13 <= io_in_c_bypass_0_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_0_is_stationary_13 <= io_in_c_bypass_0_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_1_data_13 <= io_in_c_bypass_0_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_1_is_stationary_13 <= io_in_c_bypass_0_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_2_data_13 <= io_in_c_bypass_0_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_2_is_stationary_13 <= io_in_c_bypass_0_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_3_data_13 <= io_in_c_bypass_0_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_3_is_stationary_13 <= io_in_c_bypass_0_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_0_data_13 <= io_in_c_bypass_1_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_0_is_stationary_13 <= io_in_c_bypass_1_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_1_data_13 <= io_in_c_bypass_1_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_1_is_stationary_13 <= io_in_c_bypass_1_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_2_data_13 <= io_in_c_bypass_1_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_2_is_stationary_13 <= io_in_c_bypass_1_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_3_data_13 <= io_in_c_bypass_1_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_3_is_stationary_13 <= io_in_c_bypass_1_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_0_data_13 <= io_in_c_bypass_2_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_0_is_stationary_13 <= io_in_c_bypass_2_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_1_data_13 <= io_in_c_bypass_2_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_1_is_stationary_13 <= io_in_c_bypass_2_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_2_data_13 <= io_in_c_bypass_2_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_2_is_stationary_13 <= io_in_c_bypass_2_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_3_data_13 <= io_in_c_bypass_2_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_3_is_stationary_13 <= io_in_c_bypass_2_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_0_data_13 <= io_in_c_bypass_3_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_0_is_stationary_13 <= io_in_c_bypass_3_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_1_data_13 <= io_in_c_bypass_3_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_1_is_stationary_13 <= io_in_c_bypass_3_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_2_data_13 <= io_in_c_bypass_3_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_2_is_stationary_13 <= io_in_c_bypass_3_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_3_data_13 <= io_in_c_bypass_3_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_3_is_stationary_13 <= io_in_c_bypass_3_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_0_data_13 <= io_in_c_bypass_4_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_0_is_stationary_13 <= io_in_c_bypass_4_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_1_data_13 <= io_in_c_bypass_4_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_1_is_stationary_13 <= io_in_c_bypass_4_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_2_data_13 <= io_in_c_bypass_4_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_2_is_stationary_13 <= io_in_c_bypass_4_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_3_data_13 <= io_in_c_bypass_4_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_3_is_stationary_13 <= io_in_c_bypass_4_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_0_data_13 <= io_in_c_bypass_5_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_0_is_stationary_13 <= io_in_c_bypass_5_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_1_data_13 <= io_in_c_bypass_5_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_1_is_stationary_13 <= io_in_c_bypass_5_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_2_data_13 <= io_in_c_bypass_5_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_2_is_stationary_13 <= io_in_c_bypass_5_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_3_data_13 <= io_in_c_bypass_5_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_3_is_stationary_13 <= io_in_c_bypass_5_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_0_data_13 <= io_in_c_bypass_6_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_0_is_stationary_13 <= io_in_c_bypass_6_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_1_data_13 <= io_in_c_bypass_6_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_1_is_stationary_13 <= io_in_c_bypass_6_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_2_data_13 <= io_in_c_bypass_6_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_2_is_stationary_13 <= io_in_c_bypass_6_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_3_data_13 <= io_in_c_bypass_6_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_3_is_stationary_13 <= io_in_c_bypass_6_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_0_data_13 <= io_in_c_bypass_7_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_0_is_stationary_13 <= io_in_c_bypass_7_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_1_data_13 <= io_in_c_bypass_7_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_1_is_stationary_13 <= io_in_c_bypass_7_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_2_data_13 <= io_in_c_bypass_7_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_2_is_stationary_13 <= io_in_c_bypass_7_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_3_data_13 <= io_in_c_bypass_7_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_3_is_stationary_13 <= io_in_c_bypass_7_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_0_data_13 <= io_in_c_bypass_8_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_0_is_stationary_13 <= io_in_c_bypass_8_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_1_data_13 <= io_in_c_bypass_8_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_1_is_stationary_13 <= io_in_c_bypass_8_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_2_data_13 <= io_in_c_bypass_8_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_2_is_stationary_13 <= io_in_c_bypass_8_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_3_data_13 <= io_in_c_bypass_8_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_3_is_stationary_13 <= io_in_c_bypass_8_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_0_data_13 <= io_in_c_bypass_9_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_0_is_stationary_13 <= io_in_c_bypass_9_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_1_data_13 <= io_in_c_bypass_9_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_1_is_stationary_13 <= io_in_c_bypass_9_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_2_data_13 <= io_in_c_bypass_9_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_2_is_stationary_13 <= io_in_c_bypass_9_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_3_data_13 <= io_in_c_bypass_9_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_3_is_stationary_13 <= io_in_c_bypass_9_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_0_data_13 <= io_in_c_bypass_10_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_0_is_stationary_13 <= io_in_c_bypass_10_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_1_data_13 <= io_in_c_bypass_10_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_1_is_stationary_13 <= io_in_c_bypass_10_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_2_data_13 <= io_in_c_bypass_10_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_2_is_stationary_13 <= io_in_c_bypass_10_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_3_data_13 <= io_in_c_bypass_10_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_3_is_stationary_13 <= io_in_c_bypass_10_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_0_data_13 <= io_in_c_bypass_11_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_0_is_stationary_13 <= io_in_c_bypass_11_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_1_data_13 <= io_in_c_bypass_11_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_1_is_stationary_13 <= io_in_c_bypass_11_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_2_data_13 <= io_in_c_bypass_11_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_2_is_stationary_13 <= io_in_c_bypass_11_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_3_data_13 <= io_in_c_bypass_11_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_3_is_stationary_13 <= io_in_c_bypass_11_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_0_data_13 <= io_in_c_bypass_12_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_0_is_stationary_13 <= io_in_c_bypass_12_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_1_data_13 <= io_in_c_bypass_12_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_1_is_stationary_13 <= io_in_c_bypass_12_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_2_data_13 <= io_in_c_bypass_12_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_2_is_stationary_13 <= io_in_c_bypass_12_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_3_data_13 <= io_in_c_bypass_12_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_3_is_stationary_13 <= io_in_c_bypass_12_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_0_data_13 <= io_in_c_bypass_13_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_0_is_stationary_13 <= io_in_c_bypass_13_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_1_data_13 <= io_in_c_bypass_13_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_1_is_stationary_13 <= io_in_c_bypass_13_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_2_data_13 <= io_in_c_bypass_13_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_2_is_stationary_13 <= io_in_c_bypass_13_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_3_data_13 <= io_in_c_bypass_13_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_3_is_stationary_13 <= io_in_c_bypass_13_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_0_data_13 <= io_in_c_bypass_14_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_0_is_stationary_13 <= io_in_c_bypass_14_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_1_data_13 <= io_in_c_bypass_14_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_1_is_stationary_13 <= io_in_c_bypass_14_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_2_data_13 <= io_in_c_bypass_14_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_2_is_stationary_13 <= io_in_c_bypass_14_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_3_data_13 <= io_in_c_bypass_14_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_3_is_stationary_13 <= io_in_c_bypass_14_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_0_data_13 <= io_in_c_bypass_15_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_0_is_stationary_13 <= io_in_c_bypass_15_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_1_data_13 <= io_in_c_bypass_15_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_1_is_stationary_13 <= io_in_c_bypass_15_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_2_data_13 <= io_in_c_bypass_15_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_2_is_stationary_13 <= io_in_c_bypass_15_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_3_data_13 <= io_in_c_bypass_15_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_3_is_stationary_13 <= io_in_c_bypass_15_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_0_data_13 <= io_in_c_bypass_16_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_0_is_stationary_13 <= io_in_c_bypass_16_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_1_data_13 <= io_in_c_bypass_16_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_1_is_stationary_13 <= io_in_c_bypass_16_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_2_data_13 <= io_in_c_bypass_16_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_2_is_stationary_13 <= io_in_c_bypass_16_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_3_data_13 <= io_in_c_bypass_16_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_3_is_stationary_13 <= io_in_c_bypass_16_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_0_data_13 <= io_in_c_bypass_17_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_0_is_stationary_13 <= io_in_c_bypass_17_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_1_data_13 <= io_in_c_bypass_17_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_1_is_stationary_13 <= io_in_c_bypass_17_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_2_data_13 <= io_in_c_bypass_17_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_2_is_stationary_13 <= io_in_c_bypass_17_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_3_data_13 <= io_in_c_bypass_17_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_3_is_stationary_13 <= io_in_c_bypass_17_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_0_data_13 <= io_in_c_bypass_18_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_0_is_stationary_13 <= io_in_c_bypass_18_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_1_data_13 <= io_in_c_bypass_18_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_1_is_stationary_13 <= io_in_c_bypass_18_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_2_data_13 <= io_in_c_bypass_18_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_2_is_stationary_13 <= io_in_c_bypass_18_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_3_data_13 <= io_in_c_bypass_18_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_3_is_stationary_13 <= io_in_c_bypass_18_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_0_data_13 <= io_in_c_bypass_19_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_0_is_stationary_13 <= io_in_c_bypass_19_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_1_data_13 <= io_in_c_bypass_19_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_1_is_stationary_13 <= io_in_c_bypass_19_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_2_data_13 <= io_in_c_bypass_19_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_2_is_stationary_13 <= io_in_c_bypass_19_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_3_data_13 <= io_in_c_bypass_19_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_3_is_stationary_13 <= io_in_c_bypass_19_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_0_data_13 <= io_in_c_bypass_20_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_0_is_stationary_13 <= io_in_c_bypass_20_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_1_data_13 <= io_in_c_bypass_20_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_1_is_stationary_13 <= io_in_c_bypass_20_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_2_data_13 <= io_in_c_bypass_20_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_2_is_stationary_13 <= io_in_c_bypass_20_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_3_data_13 <= io_in_c_bypass_20_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_3_is_stationary_13 <= io_in_c_bypass_20_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_0_data_13 <= io_in_c_bypass_21_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_0_is_stationary_13 <= io_in_c_bypass_21_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_1_data_13 <= io_in_c_bypass_21_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_1_is_stationary_13 <= io_in_c_bypass_21_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_2_data_13 <= io_in_c_bypass_21_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_2_is_stationary_13 <= io_in_c_bypass_21_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_3_data_13 <= io_in_c_bypass_21_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_3_is_stationary_13 <= io_in_c_bypass_21_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_0_data_13 <= io_in_c_bypass_22_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_0_is_stationary_13 <= io_in_c_bypass_22_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_1_data_13 <= io_in_c_bypass_22_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_1_is_stationary_13 <= io_in_c_bypass_22_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_2_data_13 <= io_in_c_bypass_22_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_2_is_stationary_13 <= io_in_c_bypass_22_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_3_data_13 <= io_in_c_bypass_22_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_3_is_stationary_13 <= io_in_c_bypass_22_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_0_data_13 <= io_in_c_bypass_23_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_0_is_stationary_13 <= io_in_c_bypass_23_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_1_data_13 <= io_in_c_bypass_23_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_1_is_stationary_13 <= io_in_c_bypass_23_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_2_data_13 <= io_in_c_bypass_23_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_2_is_stationary_13 <= io_in_c_bypass_23_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_3_data_13 <= io_in_c_bypass_23_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_3_is_stationary_13 <= io_in_c_bypass_23_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_0_data_13 <= io_in_c_bypass_24_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_0_is_stationary_13 <= io_in_c_bypass_24_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_1_data_13 <= io_in_c_bypass_24_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_1_is_stationary_13 <= io_in_c_bypass_24_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_2_data_13 <= io_in_c_bypass_24_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_2_is_stationary_13 <= io_in_c_bypass_24_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_3_data_13 <= io_in_c_bypass_24_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_3_is_stationary_13 <= io_in_c_bypass_24_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_0_data_13 <= io_in_c_bypass_25_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_0_is_stationary_13 <= io_in_c_bypass_25_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_1_data_13 <= io_in_c_bypass_25_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_1_is_stationary_13 <= io_in_c_bypass_25_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_2_data_13 <= io_in_c_bypass_25_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_2_is_stationary_13 <= io_in_c_bypass_25_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_3_data_13 <= io_in_c_bypass_25_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_3_is_stationary_13 <= io_in_c_bypass_25_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_0_data_13 <= io_in_c_bypass_26_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_0_is_stationary_13 <= io_in_c_bypass_26_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_1_data_13 <= io_in_c_bypass_26_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_1_is_stationary_13 <= io_in_c_bypass_26_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_2_data_13 <= io_in_c_bypass_26_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_2_is_stationary_13 <= io_in_c_bypass_26_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_3_data_13 <= io_in_c_bypass_26_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_3_is_stationary_13 <= io_in_c_bypass_26_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_0_data_13 <= io_in_c_bypass_27_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_0_is_stationary_13 <= io_in_c_bypass_27_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_1_data_13 <= io_in_c_bypass_27_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_1_is_stationary_13 <= io_in_c_bypass_27_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_2_data_13 <= io_in_c_bypass_27_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_2_is_stationary_13 <= io_in_c_bypass_27_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_3_data_13 <= io_in_c_bypass_27_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_3_is_stationary_13 <= io_in_c_bypass_27_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_0_data_13 <= io_in_c_bypass_28_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_0_is_stationary_13 <= io_in_c_bypass_28_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_1_data_13 <= io_in_c_bypass_28_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_1_is_stationary_13 <= io_in_c_bypass_28_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_2_data_13 <= io_in_c_bypass_28_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_2_is_stationary_13 <= io_in_c_bypass_28_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_3_data_13 <= io_in_c_bypass_28_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_3_is_stationary_13 <= io_in_c_bypass_28_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_0_data_13 <= io_in_c_bypass_29_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_0_is_stationary_13 <= io_in_c_bypass_29_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_1_data_13 <= io_in_c_bypass_29_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_1_is_stationary_13 <= io_in_c_bypass_29_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_2_data_13 <= io_in_c_bypass_29_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_2_is_stationary_13 <= io_in_c_bypass_29_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_3_data_13 <= io_in_c_bypass_29_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_3_is_stationary_13 <= io_in_c_bypass_29_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_0_data_13 <= io_in_c_bypass_30_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_0_is_stationary_13 <= io_in_c_bypass_30_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_1_data_13 <= io_in_c_bypass_30_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_1_is_stationary_13 <= io_in_c_bypass_30_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_2_data_13 <= io_in_c_bypass_30_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_2_is_stationary_13 <= io_in_c_bypass_30_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_3_data_13 <= io_in_c_bypass_30_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_3_is_stationary_13 <= io_in_c_bypass_30_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_0_data_13 <= io_in_c_bypass_31_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_0_is_stationary_13 <= io_in_c_bypass_31_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_1_data_13 <= io_in_c_bypass_31_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_1_is_stationary_13 <= io_in_c_bypass_31_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_2_data_13 <= io_in_c_bypass_31_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_2_is_stationary_13 <= io_in_c_bypass_31_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_3_data_13 <= io_in_c_bypass_31_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_3_is_stationary_13 <= io_in_c_bypass_31_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_0_data_14 <= io_in_c_bypass_0_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_0_is_stationary_14 <= io_in_c_bypass_0_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_1_data_14 <= io_in_c_bypass_0_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_1_is_stationary_14 <= io_in_c_bypass_0_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_2_data_14 <= io_in_c_bypass_0_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_2_is_stationary_14 <= io_in_c_bypass_0_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_3_data_14 <= io_in_c_bypass_0_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_3_is_stationary_14 <= io_in_c_bypass_0_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_0_data_14 <= io_in_c_bypass_1_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_0_is_stationary_14 <= io_in_c_bypass_1_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_1_data_14 <= io_in_c_bypass_1_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_1_is_stationary_14 <= io_in_c_bypass_1_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_2_data_14 <= io_in_c_bypass_1_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_2_is_stationary_14 <= io_in_c_bypass_1_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_3_data_14 <= io_in_c_bypass_1_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_3_is_stationary_14 <= io_in_c_bypass_1_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_0_data_14 <= io_in_c_bypass_2_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_0_is_stationary_14 <= io_in_c_bypass_2_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_1_data_14 <= io_in_c_bypass_2_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_1_is_stationary_14 <= io_in_c_bypass_2_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_2_data_14 <= io_in_c_bypass_2_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_2_is_stationary_14 <= io_in_c_bypass_2_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_3_data_14 <= io_in_c_bypass_2_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_3_is_stationary_14 <= io_in_c_bypass_2_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_0_data_14 <= io_in_c_bypass_3_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_0_is_stationary_14 <= io_in_c_bypass_3_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_1_data_14 <= io_in_c_bypass_3_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_1_is_stationary_14 <= io_in_c_bypass_3_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_2_data_14 <= io_in_c_bypass_3_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_2_is_stationary_14 <= io_in_c_bypass_3_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_3_data_14 <= io_in_c_bypass_3_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_3_is_stationary_14 <= io_in_c_bypass_3_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_0_data_14 <= io_in_c_bypass_4_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_0_is_stationary_14 <= io_in_c_bypass_4_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_1_data_14 <= io_in_c_bypass_4_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_1_is_stationary_14 <= io_in_c_bypass_4_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_2_data_14 <= io_in_c_bypass_4_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_2_is_stationary_14 <= io_in_c_bypass_4_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_3_data_14 <= io_in_c_bypass_4_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_3_is_stationary_14 <= io_in_c_bypass_4_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_0_data_14 <= io_in_c_bypass_5_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_0_is_stationary_14 <= io_in_c_bypass_5_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_1_data_14 <= io_in_c_bypass_5_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_1_is_stationary_14 <= io_in_c_bypass_5_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_2_data_14 <= io_in_c_bypass_5_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_2_is_stationary_14 <= io_in_c_bypass_5_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_3_data_14 <= io_in_c_bypass_5_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_3_is_stationary_14 <= io_in_c_bypass_5_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_0_data_14 <= io_in_c_bypass_6_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_0_is_stationary_14 <= io_in_c_bypass_6_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_1_data_14 <= io_in_c_bypass_6_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_1_is_stationary_14 <= io_in_c_bypass_6_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_2_data_14 <= io_in_c_bypass_6_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_2_is_stationary_14 <= io_in_c_bypass_6_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_3_data_14 <= io_in_c_bypass_6_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_3_is_stationary_14 <= io_in_c_bypass_6_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_0_data_14 <= io_in_c_bypass_7_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_0_is_stationary_14 <= io_in_c_bypass_7_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_1_data_14 <= io_in_c_bypass_7_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_1_is_stationary_14 <= io_in_c_bypass_7_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_2_data_14 <= io_in_c_bypass_7_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_2_is_stationary_14 <= io_in_c_bypass_7_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_3_data_14 <= io_in_c_bypass_7_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_3_is_stationary_14 <= io_in_c_bypass_7_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_0_data_14 <= io_in_c_bypass_8_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_0_is_stationary_14 <= io_in_c_bypass_8_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_1_data_14 <= io_in_c_bypass_8_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_1_is_stationary_14 <= io_in_c_bypass_8_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_2_data_14 <= io_in_c_bypass_8_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_2_is_stationary_14 <= io_in_c_bypass_8_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_3_data_14 <= io_in_c_bypass_8_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_3_is_stationary_14 <= io_in_c_bypass_8_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_0_data_14 <= io_in_c_bypass_9_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_0_is_stationary_14 <= io_in_c_bypass_9_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_1_data_14 <= io_in_c_bypass_9_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_1_is_stationary_14 <= io_in_c_bypass_9_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_2_data_14 <= io_in_c_bypass_9_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_2_is_stationary_14 <= io_in_c_bypass_9_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_3_data_14 <= io_in_c_bypass_9_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_3_is_stationary_14 <= io_in_c_bypass_9_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_0_data_14 <= io_in_c_bypass_10_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_0_is_stationary_14 <= io_in_c_bypass_10_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_1_data_14 <= io_in_c_bypass_10_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_1_is_stationary_14 <= io_in_c_bypass_10_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_2_data_14 <= io_in_c_bypass_10_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_2_is_stationary_14 <= io_in_c_bypass_10_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_3_data_14 <= io_in_c_bypass_10_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_3_is_stationary_14 <= io_in_c_bypass_10_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_0_data_14 <= io_in_c_bypass_11_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_0_is_stationary_14 <= io_in_c_bypass_11_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_1_data_14 <= io_in_c_bypass_11_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_1_is_stationary_14 <= io_in_c_bypass_11_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_2_data_14 <= io_in_c_bypass_11_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_2_is_stationary_14 <= io_in_c_bypass_11_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_3_data_14 <= io_in_c_bypass_11_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_3_is_stationary_14 <= io_in_c_bypass_11_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_0_data_14 <= io_in_c_bypass_12_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_0_is_stationary_14 <= io_in_c_bypass_12_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_1_data_14 <= io_in_c_bypass_12_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_1_is_stationary_14 <= io_in_c_bypass_12_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_2_data_14 <= io_in_c_bypass_12_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_2_is_stationary_14 <= io_in_c_bypass_12_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_3_data_14 <= io_in_c_bypass_12_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_3_is_stationary_14 <= io_in_c_bypass_12_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_0_data_14 <= io_in_c_bypass_13_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_0_is_stationary_14 <= io_in_c_bypass_13_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_1_data_14 <= io_in_c_bypass_13_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_1_is_stationary_14 <= io_in_c_bypass_13_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_2_data_14 <= io_in_c_bypass_13_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_2_is_stationary_14 <= io_in_c_bypass_13_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_3_data_14 <= io_in_c_bypass_13_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_3_is_stationary_14 <= io_in_c_bypass_13_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_0_data_14 <= io_in_c_bypass_14_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_0_is_stationary_14 <= io_in_c_bypass_14_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_1_data_14 <= io_in_c_bypass_14_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_1_is_stationary_14 <= io_in_c_bypass_14_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_2_data_14 <= io_in_c_bypass_14_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_2_is_stationary_14 <= io_in_c_bypass_14_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_3_data_14 <= io_in_c_bypass_14_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_3_is_stationary_14 <= io_in_c_bypass_14_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_0_data_14 <= io_in_c_bypass_15_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_0_is_stationary_14 <= io_in_c_bypass_15_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_1_data_14 <= io_in_c_bypass_15_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_1_is_stationary_14 <= io_in_c_bypass_15_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_2_data_14 <= io_in_c_bypass_15_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_2_is_stationary_14 <= io_in_c_bypass_15_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_3_data_14 <= io_in_c_bypass_15_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_3_is_stationary_14 <= io_in_c_bypass_15_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_0_data_14 <= io_in_c_bypass_16_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_0_is_stationary_14 <= io_in_c_bypass_16_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_1_data_14 <= io_in_c_bypass_16_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_1_is_stationary_14 <= io_in_c_bypass_16_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_2_data_14 <= io_in_c_bypass_16_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_2_is_stationary_14 <= io_in_c_bypass_16_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_3_data_14 <= io_in_c_bypass_16_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_3_is_stationary_14 <= io_in_c_bypass_16_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_0_data_14 <= io_in_c_bypass_17_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_0_is_stationary_14 <= io_in_c_bypass_17_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_1_data_14 <= io_in_c_bypass_17_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_1_is_stationary_14 <= io_in_c_bypass_17_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_2_data_14 <= io_in_c_bypass_17_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_2_is_stationary_14 <= io_in_c_bypass_17_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_3_data_14 <= io_in_c_bypass_17_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_3_is_stationary_14 <= io_in_c_bypass_17_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_0_data_14 <= io_in_c_bypass_18_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_0_is_stationary_14 <= io_in_c_bypass_18_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_1_data_14 <= io_in_c_bypass_18_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_1_is_stationary_14 <= io_in_c_bypass_18_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_2_data_14 <= io_in_c_bypass_18_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_2_is_stationary_14 <= io_in_c_bypass_18_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_3_data_14 <= io_in_c_bypass_18_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_3_is_stationary_14 <= io_in_c_bypass_18_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_0_data_14 <= io_in_c_bypass_19_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_0_is_stationary_14 <= io_in_c_bypass_19_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_1_data_14 <= io_in_c_bypass_19_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_1_is_stationary_14 <= io_in_c_bypass_19_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_2_data_14 <= io_in_c_bypass_19_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_2_is_stationary_14 <= io_in_c_bypass_19_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_3_data_14 <= io_in_c_bypass_19_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_3_is_stationary_14 <= io_in_c_bypass_19_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_0_data_14 <= io_in_c_bypass_20_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_0_is_stationary_14 <= io_in_c_bypass_20_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_1_data_14 <= io_in_c_bypass_20_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_1_is_stationary_14 <= io_in_c_bypass_20_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_2_data_14 <= io_in_c_bypass_20_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_2_is_stationary_14 <= io_in_c_bypass_20_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_3_data_14 <= io_in_c_bypass_20_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_3_is_stationary_14 <= io_in_c_bypass_20_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_0_data_14 <= io_in_c_bypass_21_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_0_is_stationary_14 <= io_in_c_bypass_21_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_1_data_14 <= io_in_c_bypass_21_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_1_is_stationary_14 <= io_in_c_bypass_21_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_2_data_14 <= io_in_c_bypass_21_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_2_is_stationary_14 <= io_in_c_bypass_21_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_3_data_14 <= io_in_c_bypass_21_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_3_is_stationary_14 <= io_in_c_bypass_21_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_0_data_14 <= io_in_c_bypass_22_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_0_is_stationary_14 <= io_in_c_bypass_22_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_1_data_14 <= io_in_c_bypass_22_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_1_is_stationary_14 <= io_in_c_bypass_22_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_2_data_14 <= io_in_c_bypass_22_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_2_is_stationary_14 <= io_in_c_bypass_22_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_3_data_14 <= io_in_c_bypass_22_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_3_is_stationary_14 <= io_in_c_bypass_22_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_0_data_14 <= io_in_c_bypass_23_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_0_is_stationary_14 <= io_in_c_bypass_23_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_1_data_14 <= io_in_c_bypass_23_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_1_is_stationary_14 <= io_in_c_bypass_23_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_2_data_14 <= io_in_c_bypass_23_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_2_is_stationary_14 <= io_in_c_bypass_23_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_3_data_14 <= io_in_c_bypass_23_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_3_is_stationary_14 <= io_in_c_bypass_23_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_0_data_14 <= io_in_c_bypass_24_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_0_is_stationary_14 <= io_in_c_bypass_24_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_1_data_14 <= io_in_c_bypass_24_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_1_is_stationary_14 <= io_in_c_bypass_24_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_2_data_14 <= io_in_c_bypass_24_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_2_is_stationary_14 <= io_in_c_bypass_24_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_3_data_14 <= io_in_c_bypass_24_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_3_is_stationary_14 <= io_in_c_bypass_24_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_0_data_14 <= io_in_c_bypass_25_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_0_is_stationary_14 <= io_in_c_bypass_25_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_1_data_14 <= io_in_c_bypass_25_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_1_is_stationary_14 <= io_in_c_bypass_25_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_2_data_14 <= io_in_c_bypass_25_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_2_is_stationary_14 <= io_in_c_bypass_25_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_3_data_14 <= io_in_c_bypass_25_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_3_is_stationary_14 <= io_in_c_bypass_25_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_0_data_14 <= io_in_c_bypass_26_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_0_is_stationary_14 <= io_in_c_bypass_26_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_1_data_14 <= io_in_c_bypass_26_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_1_is_stationary_14 <= io_in_c_bypass_26_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_2_data_14 <= io_in_c_bypass_26_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_2_is_stationary_14 <= io_in_c_bypass_26_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_3_data_14 <= io_in_c_bypass_26_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_3_is_stationary_14 <= io_in_c_bypass_26_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_0_data_14 <= io_in_c_bypass_27_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_0_is_stationary_14 <= io_in_c_bypass_27_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_1_data_14 <= io_in_c_bypass_27_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_1_is_stationary_14 <= io_in_c_bypass_27_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_2_data_14 <= io_in_c_bypass_27_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_2_is_stationary_14 <= io_in_c_bypass_27_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_3_data_14 <= io_in_c_bypass_27_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_3_is_stationary_14 <= io_in_c_bypass_27_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_0_data_14 <= io_in_c_bypass_28_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_0_is_stationary_14 <= io_in_c_bypass_28_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_1_data_14 <= io_in_c_bypass_28_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_1_is_stationary_14 <= io_in_c_bypass_28_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_2_data_14 <= io_in_c_bypass_28_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_2_is_stationary_14 <= io_in_c_bypass_28_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_3_data_14 <= io_in_c_bypass_28_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_3_is_stationary_14 <= io_in_c_bypass_28_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_0_data_14 <= io_in_c_bypass_29_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_0_is_stationary_14 <= io_in_c_bypass_29_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_1_data_14 <= io_in_c_bypass_29_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_1_is_stationary_14 <= io_in_c_bypass_29_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_2_data_14 <= io_in_c_bypass_29_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_2_is_stationary_14 <= io_in_c_bypass_29_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_3_data_14 <= io_in_c_bypass_29_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_3_is_stationary_14 <= io_in_c_bypass_29_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_0_data_14 <= io_in_c_bypass_30_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_0_is_stationary_14 <= io_in_c_bypass_30_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_1_data_14 <= io_in_c_bypass_30_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_1_is_stationary_14 <= io_in_c_bypass_30_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_2_data_14 <= io_in_c_bypass_30_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_2_is_stationary_14 <= io_in_c_bypass_30_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_3_data_14 <= io_in_c_bypass_30_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_3_is_stationary_14 <= io_in_c_bypass_30_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_0_data_14 <= io_in_c_bypass_31_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_0_is_stationary_14 <= io_in_c_bypass_31_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_1_data_14 <= io_in_c_bypass_31_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_1_is_stationary_14 <= io_in_c_bypass_31_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_2_data_14 <= io_in_c_bypass_31_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_2_is_stationary_14 <= io_in_c_bypass_31_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_3_data_14 <= io_in_c_bypass_31_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_3_is_stationary_14 <= io_in_c_bypass_31_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_0_data_15 <= io_in_c_bypass_0_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_0_is_stationary_15 <= io_in_c_bypass_0_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_1_data_15 <= io_in_c_bypass_0_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_1_is_stationary_15 <= io_in_c_bypass_0_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_2_data_15 <= io_in_c_bypass_0_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_2_is_stationary_15 <= io_in_c_bypass_0_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_3_data_15 <= io_in_c_bypass_0_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_3_is_stationary_15 <= io_in_c_bypass_0_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_0_data_15 <= io_in_c_bypass_1_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_0_is_stationary_15 <= io_in_c_bypass_1_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_1_data_15 <= io_in_c_bypass_1_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_1_is_stationary_15 <= io_in_c_bypass_1_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_2_data_15 <= io_in_c_bypass_1_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_2_is_stationary_15 <= io_in_c_bypass_1_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_3_data_15 <= io_in_c_bypass_1_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_3_is_stationary_15 <= io_in_c_bypass_1_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_0_data_15 <= io_in_c_bypass_2_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_0_is_stationary_15 <= io_in_c_bypass_2_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_1_data_15 <= io_in_c_bypass_2_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_1_is_stationary_15 <= io_in_c_bypass_2_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_2_data_15 <= io_in_c_bypass_2_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_2_is_stationary_15 <= io_in_c_bypass_2_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_3_data_15 <= io_in_c_bypass_2_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_3_is_stationary_15 <= io_in_c_bypass_2_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_0_data_15 <= io_in_c_bypass_3_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_0_is_stationary_15 <= io_in_c_bypass_3_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_1_data_15 <= io_in_c_bypass_3_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_1_is_stationary_15 <= io_in_c_bypass_3_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_2_data_15 <= io_in_c_bypass_3_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_2_is_stationary_15 <= io_in_c_bypass_3_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_3_data_15 <= io_in_c_bypass_3_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_3_is_stationary_15 <= io_in_c_bypass_3_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_0_data_15 <= io_in_c_bypass_4_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_0_is_stationary_15 <= io_in_c_bypass_4_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_1_data_15 <= io_in_c_bypass_4_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_1_is_stationary_15 <= io_in_c_bypass_4_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_2_data_15 <= io_in_c_bypass_4_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_2_is_stationary_15 <= io_in_c_bypass_4_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_3_data_15 <= io_in_c_bypass_4_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_3_is_stationary_15 <= io_in_c_bypass_4_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_0_data_15 <= io_in_c_bypass_5_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_0_is_stationary_15 <= io_in_c_bypass_5_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_1_data_15 <= io_in_c_bypass_5_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_1_is_stationary_15 <= io_in_c_bypass_5_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_2_data_15 <= io_in_c_bypass_5_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_2_is_stationary_15 <= io_in_c_bypass_5_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_3_data_15 <= io_in_c_bypass_5_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_3_is_stationary_15 <= io_in_c_bypass_5_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_0_data_15 <= io_in_c_bypass_6_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_0_is_stationary_15 <= io_in_c_bypass_6_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_1_data_15 <= io_in_c_bypass_6_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_1_is_stationary_15 <= io_in_c_bypass_6_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_2_data_15 <= io_in_c_bypass_6_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_2_is_stationary_15 <= io_in_c_bypass_6_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_3_data_15 <= io_in_c_bypass_6_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_3_is_stationary_15 <= io_in_c_bypass_6_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_0_data_15 <= io_in_c_bypass_7_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_0_is_stationary_15 <= io_in_c_bypass_7_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_1_data_15 <= io_in_c_bypass_7_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_1_is_stationary_15 <= io_in_c_bypass_7_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_2_data_15 <= io_in_c_bypass_7_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_2_is_stationary_15 <= io_in_c_bypass_7_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_3_data_15 <= io_in_c_bypass_7_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_3_is_stationary_15 <= io_in_c_bypass_7_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_0_data_15 <= io_in_c_bypass_8_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_0_is_stationary_15 <= io_in_c_bypass_8_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_1_data_15 <= io_in_c_bypass_8_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_1_is_stationary_15 <= io_in_c_bypass_8_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_2_data_15 <= io_in_c_bypass_8_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_2_is_stationary_15 <= io_in_c_bypass_8_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_3_data_15 <= io_in_c_bypass_8_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_3_is_stationary_15 <= io_in_c_bypass_8_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_0_data_15 <= io_in_c_bypass_9_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_0_is_stationary_15 <= io_in_c_bypass_9_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_1_data_15 <= io_in_c_bypass_9_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_1_is_stationary_15 <= io_in_c_bypass_9_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_2_data_15 <= io_in_c_bypass_9_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_2_is_stationary_15 <= io_in_c_bypass_9_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_3_data_15 <= io_in_c_bypass_9_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_3_is_stationary_15 <= io_in_c_bypass_9_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_0_data_15 <= io_in_c_bypass_10_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_0_is_stationary_15 <= io_in_c_bypass_10_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_1_data_15 <= io_in_c_bypass_10_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_1_is_stationary_15 <= io_in_c_bypass_10_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_2_data_15 <= io_in_c_bypass_10_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_2_is_stationary_15 <= io_in_c_bypass_10_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_3_data_15 <= io_in_c_bypass_10_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_3_is_stationary_15 <= io_in_c_bypass_10_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_0_data_15 <= io_in_c_bypass_11_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_0_is_stationary_15 <= io_in_c_bypass_11_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_1_data_15 <= io_in_c_bypass_11_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_1_is_stationary_15 <= io_in_c_bypass_11_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_2_data_15 <= io_in_c_bypass_11_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_2_is_stationary_15 <= io_in_c_bypass_11_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_3_data_15 <= io_in_c_bypass_11_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_3_is_stationary_15 <= io_in_c_bypass_11_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_0_data_15 <= io_in_c_bypass_12_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_0_is_stationary_15 <= io_in_c_bypass_12_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_1_data_15 <= io_in_c_bypass_12_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_1_is_stationary_15 <= io_in_c_bypass_12_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_2_data_15 <= io_in_c_bypass_12_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_2_is_stationary_15 <= io_in_c_bypass_12_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_3_data_15 <= io_in_c_bypass_12_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_3_is_stationary_15 <= io_in_c_bypass_12_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_0_data_15 <= io_in_c_bypass_13_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_0_is_stationary_15 <= io_in_c_bypass_13_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_1_data_15 <= io_in_c_bypass_13_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_1_is_stationary_15 <= io_in_c_bypass_13_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_2_data_15 <= io_in_c_bypass_13_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_2_is_stationary_15 <= io_in_c_bypass_13_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_3_data_15 <= io_in_c_bypass_13_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_3_is_stationary_15 <= io_in_c_bypass_13_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_0_data_15 <= io_in_c_bypass_14_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_0_is_stationary_15 <= io_in_c_bypass_14_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_1_data_15 <= io_in_c_bypass_14_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_1_is_stationary_15 <= io_in_c_bypass_14_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_2_data_15 <= io_in_c_bypass_14_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_2_is_stationary_15 <= io_in_c_bypass_14_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_3_data_15 <= io_in_c_bypass_14_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_3_is_stationary_15 <= io_in_c_bypass_14_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_0_data_15 <= io_in_c_bypass_15_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_0_is_stationary_15 <= io_in_c_bypass_15_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_1_data_15 <= io_in_c_bypass_15_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_1_is_stationary_15 <= io_in_c_bypass_15_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_2_data_15 <= io_in_c_bypass_15_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_2_is_stationary_15 <= io_in_c_bypass_15_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_3_data_15 <= io_in_c_bypass_15_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_3_is_stationary_15 <= io_in_c_bypass_15_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_0_data_15 <= io_in_c_bypass_16_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_0_is_stationary_15 <= io_in_c_bypass_16_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_1_data_15 <= io_in_c_bypass_16_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_1_is_stationary_15 <= io_in_c_bypass_16_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_2_data_15 <= io_in_c_bypass_16_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_2_is_stationary_15 <= io_in_c_bypass_16_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_3_data_15 <= io_in_c_bypass_16_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_3_is_stationary_15 <= io_in_c_bypass_16_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_0_data_15 <= io_in_c_bypass_17_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_0_is_stationary_15 <= io_in_c_bypass_17_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_1_data_15 <= io_in_c_bypass_17_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_1_is_stationary_15 <= io_in_c_bypass_17_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_2_data_15 <= io_in_c_bypass_17_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_2_is_stationary_15 <= io_in_c_bypass_17_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_3_data_15 <= io_in_c_bypass_17_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_3_is_stationary_15 <= io_in_c_bypass_17_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_0_data_15 <= io_in_c_bypass_18_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_0_is_stationary_15 <= io_in_c_bypass_18_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_1_data_15 <= io_in_c_bypass_18_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_1_is_stationary_15 <= io_in_c_bypass_18_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_2_data_15 <= io_in_c_bypass_18_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_2_is_stationary_15 <= io_in_c_bypass_18_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_3_data_15 <= io_in_c_bypass_18_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_3_is_stationary_15 <= io_in_c_bypass_18_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_0_data_15 <= io_in_c_bypass_19_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_0_is_stationary_15 <= io_in_c_bypass_19_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_1_data_15 <= io_in_c_bypass_19_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_1_is_stationary_15 <= io_in_c_bypass_19_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_2_data_15 <= io_in_c_bypass_19_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_2_is_stationary_15 <= io_in_c_bypass_19_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_3_data_15 <= io_in_c_bypass_19_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_3_is_stationary_15 <= io_in_c_bypass_19_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_0_data_15 <= io_in_c_bypass_20_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_0_is_stationary_15 <= io_in_c_bypass_20_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_1_data_15 <= io_in_c_bypass_20_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_1_is_stationary_15 <= io_in_c_bypass_20_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_2_data_15 <= io_in_c_bypass_20_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_2_is_stationary_15 <= io_in_c_bypass_20_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_3_data_15 <= io_in_c_bypass_20_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_3_is_stationary_15 <= io_in_c_bypass_20_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_0_data_15 <= io_in_c_bypass_21_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_0_is_stationary_15 <= io_in_c_bypass_21_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_1_data_15 <= io_in_c_bypass_21_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_1_is_stationary_15 <= io_in_c_bypass_21_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_2_data_15 <= io_in_c_bypass_21_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_2_is_stationary_15 <= io_in_c_bypass_21_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_3_data_15 <= io_in_c_bypass_21_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_3_is_stationary_15 <= io_in_c_bypass_21_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_0_data_15 <= io_in_c_bypass_22_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_0_is_stationary_15 <= io_in_c_bypass_22_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_1_data_15 <= io_in_c_bypass_22_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_1_is_stationary_15 <= io_in_c_bypass_22_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_2_data_15 <= io_in_c_bypass_22_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_2_is_stationary_15 <= io_in_c_bypass_22_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_3_data_15 <= io_in_c_bypass_22_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_3_is_stationary_15 <= io_in_c_bypass_22_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_0_data_15 <= io_in_c_bypass_23_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_0_is_stationary_15 <= io_in_c_bypass_23_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_1_data_15 <= io_in_c_bypass_23_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_1_is_stationary_15 <= io_in_c_bypass_23_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_2_data_15 <= io_in_c_bypass_23_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_2_is_stationary_15 <= io_in_c_bypass_23_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_3_data_15 <= io_in_c_bypass_23_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_3_is_stationary_15 <= io_in_c_bypass_23_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_0_data_15 <= io_in_c_bypass_24_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_0_is_stationary_15 <= io_in_c_bypass_24_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_1_data_15 <= io_in_c_bypass_24_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_1_is_stationary_15 <= io_in_c_bypass_24_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_2_data_15 <= io_in_c_bypass_24_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_2_is_stationary_15 <= io_in_c_bypass_24_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_3_data_15 <= io_in_c_bypass_24_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_3_is_stationary_15 <= io_in_c_bypass_24_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_0_data_15 <= io_in_c_bypass_25_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_0_is_stationary_15 <= io_in_c_bypass_25_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_1_data_15 <= io_in_c_bypass_25_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_1_is_stationary_15 <= io_in_c_bypass_25_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_2_data_15 <= io_in_c_bypass_25_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_2_is_stationary_15 <= io_in_c_bypass_25_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_3_data_15 <= io_in_c_bypass_25_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_3_is_stationary_15 <= io_in_c_bypass_25_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_0_data_15 <= io_in_c_bypass_26_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_0_is_stationary_15 <= io_in_c_bypass_26_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_1_data_15 <= io_in_c_bypass_26_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_1_is_stationary_15 <= io_in_c_bypass_26_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_2_data_15 <= io_in_c_bypass_26_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_2_is_stationary_15 <= io_in_c_bypass_26_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_3_data_15 <= io_in_c_bypass_26_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_3_is_stationary_15 <= io_in_c_bypass_26_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_0_data_15 <= io_in_c_bypass_27_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_0_is_stationary_15 <= io_in_c_bypass_27_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_1_data_15 <= io_in_c_bypass_27_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_1_is_stationary_15 <= io_in_c_bypass_27_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_2_data_15 <= io_in_c_bypass_27_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_2_is_stationary_15 <= io_in_c_bypass_27_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_3_data_15 <= io_in_c_bypass_27_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_3_is_stationary_15 <= io_in_c_bypass_27_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_0_data_15 <= io_in_c_bypass_28_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_0_is_stationary_15 <= io_in_c_bypass_28_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_1_data_15 <= io_in_c_bypass_28_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_1_is_stationary_15 <= io_in_c_bypass_28_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_2_data_15 <= io_in_c_bypass_28_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_2_is_stationary_15 <= io_in_c_bypass_28_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_3_data_15 <= io_in_c_bypass_28_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_3_is_stationary_15 <= io_in_c_bypass_28_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_0_data_15 <= io_in_c_bypass_29_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_0_is_stationary_15 <= io_in_c_bypass_29_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_1_data_15 <= io_in_c_bypass_29_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_1_is_stationary_15 <= io_in_c_bypass_29_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_2_data_15 <= io_in_c_bypass_29_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_2_is_stationary_15 <= io_in_c_bypass_29_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_3_data_15 <= io_in_c_bypass_29_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_3_is_stationary_15 <= io_in_c_bypass_29_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_0_data_15 <= io_in_c_bypass_30_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_0_is_stationary_15 <= io_in_c_bypass_30_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_1_data_15 <= io_in_c_bypass_30_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_1_is_stationary_15 <= io_in_c_bypass_30_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_2_data_15 <= io_in_c_bypass_30_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_2_is_stationary_15 <= io_in_c_bypass_30_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_3_data_15 <= io_in_c_bypass_30_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_3_is_stationary_15 <= io_in_c_bypass_30_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_0_data_15 <= io_in_c_bypass_31_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_0_is_stationary_15 <= io_in_c_bypass_31_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_1_data_15 <= io_in_c_bypass_31_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_1_is_stationary_15 <= io_in_c_bypass_31_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_2_data_15 <= io_in_c_bypass_31_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_2_is_stationary_15 <= io_in_c_bypass_31_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_3_data_15 <= io_in_c_bypass_31_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_3_is_stationary_15 <= io_in_c_bypass_31_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_0_data_16 <= io_in_c_bypass_0_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_0_is_stationary_16 <= io_in_c_bypass_0_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_1_data_16 <= io_in_c_bypass_0_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_1_is_stationary_16 <= io_in_c_bypass_0_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_2_data_16 <= io_in_c_bypass_0_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_2_is_stationary_16 <= io_in_c_bypass_0_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_3_data_16 <= io_in_c_bypass_0_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_3_is_stationary_16 <= io_in_c_bypass_0_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_0_data_16 <= io_in_c_bypass_1_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_0_is_stationary_16 <= io_in_c_bypass_1_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_1_data_16 <= io_in_c_bypass_1_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_1_is_stationary_16 <= io_in_c_bypass_1_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_2_data_16 <= io_in_c_bypass_1_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_2_is_stationary_16 <= io_in_c_bypass_1_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_3_data_16 <= io_in_c_bypass_1_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_3_is_stationary_16 <= io_in_c_bypass_1_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_0_data_16 <= io_in_c_bypass_2_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_0_is_stationary_16 <= io_in_c_bypass_2_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_1_data_16 <= io_in_c_bypass_2_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_1_is_stationary_16 <= io_in_c_bypass_2_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_2_data_16 <= io_in_c_bypass_2_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_2_is_stationary_16 <= io_in_c_bypass_2_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_3_data_16 <= io_in_c_bypass_2_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_3_is_stationary_16 <= io_in_c_bypass_2_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_0_data_16 <= io_in_c_bypass_3_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_0_is_stationary_16 <= io_in_c_bypass_3_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_1_data_16 <= io_in_c_bypass_3_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_1_is_stationary_16 <= io_in_c_bypass_3_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_2_data_16 <= io_in_c_bypass_3_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_2_is_stationary_16 <= io_in_c_bypass_3_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_3_data_16 <= io_in_c_bypass_3_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_3_is_stationary_16 <= io_in_c_bypass_3_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_0_data_16 <= io_in_c_bypass_4_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_0_is_stationary_16 <= io_in_c_bypass_4_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_1_data_16 <= io_in_c_bypass_4_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_1_is_stationary_16 <= io_in_c_bypass_4_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_2_data_16 <= io_in_c_bypass_4_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_2_is_stationary_16 <= io_in_c_bypass_4_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_3_data_16 <= io_in_c_bypass_4_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_3_is_stationary_16 <= io_in_c_bypass_4_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_0_data_16 <= io_in_c_bypass_5_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_0_is_stationary_16 <= io_in_c_bypass_5_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_1_data_16 <= io_in_c_bypass_5_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_1_is_stationary_16 <= io_in_c_bypass_5_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_2_data_16 <= io_in_c_bypass_5_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_2_is_stationary_16 <= io_in_c_bypass_5_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_3_data_16 <= io_in_c_bypass_5_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_3_is_stationary_16 <= io_in_c_bypass_5_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_0_data_16 <= io_in_c_bypass_6_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_0_is_stationary_16 <= io_in_c_bypass_6_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_1_data_16 <= io_in_c_bypass_6_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_1_is_stationary_16 <= io_in_c_bypass_6_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_2_data_16 <= io_in_c_bypass_6_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_2_is_stationary_16 <= io_in_c_bypass_6_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_3_data_16 <= io_in_c_bypass_6_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_3_is_stationary_16 <= io_in_c_bypass_6_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_0_data_16 <= io_in_c_bypass_7_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_0_is_stationary_16 <= io_in_c_bypass_7_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_1_data_16 <= io_in_c_bypass_7_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_1_is_stationary_16 <= io_in_c_bypass_7_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_2_data_16 <= io_in_c_bypass_7_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_2_is_stationary_16 <= io_in_c_bypass_7_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_3_data_16 <= io_in_c_bypass_7_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_3_is_stationary_16 <= io_in_c_bypass_7_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_0_data_16 <= io_in_c_bypass_8_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_0_is_stationary_16 <= io_in_c_bypass_8_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_1_data_16 <= io_in_c_bypass_8_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_1_is_stationary_16 <= io_in_c_bypass_8_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_2_data_16 <= io_in_c_bypass_8_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_2_is_stationary_16 <= io_in_c_bypass_8_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_3_data_16 <= io_in_c_bypass_8_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_3_is_stationary_16 <= io_in_c_bypass_8_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_0_data_16 <= io_in_c_bypass_9_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_0_is_stationary_16 <= io_in_c_bypass_9_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_1_data_16 <= io_in_c_bypass_9_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_1_is_stationary_16 <= io_in_c_bypass_9_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_2_data_16 <= io_in_c_bypass_9_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_2_is_stationary_16 <= io_in_c_bypass_9_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_3_data_16 <= io_in_c_bypass_9_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_3_is_stationary_16 <= io_in_c_bypass_9_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_0_data_16 <= io_in_c_bypass_10_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_0_is_stationary_16 <= io_in_c_bypass_10_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_1_data_16 <= io_in_c_bypass_10_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_1_is_stationary_16 <= io_in_c_bypass_10_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_2_data_16 <= io_in_c_bypass_10_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_2_is_stationary_16 <= io_in_c_bypass_10_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_3_data_16 <= io_in_c_bypass_10_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_3_is_stationary_16 <= io_in_c_bypass_10_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_0_data_16 <= io_in_c_bypass_11_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_0_is_stationary_16 <= io_in_c_bypass_11_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_1_data_16 <= io_in_c_bypass_11_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_1_is_stationary_16 <= io_in_c_bypass_11_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_2_data_16 <= io_in_c_bypass_11_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_2_is_stationary_16 <= io_in_c_bypass_11_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_3_data_16 <= io_in_c_bypass_11_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_3_is_stationary_16 <= io_in_c_bypass_11_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_0_data_16 <= io_in_c_bypass_12_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_0_is_stationary_16 <= io_in_c_bypass_12_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_1_data_16 <= io_in_c_bypass_12_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_1_is_stationary_16 <= io_in_c_bypass_12_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_2_data_16 <= io_in_c_bypass_12_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_2_is_stationary_16 <= io_in_c_bypass_12_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_3_data_16 <= io_in_c_bypass_12_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_3_is_stationary_16 <= io_in_c_bypass_12_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_0_data_16 <= io_in_c_bypass_13_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_0_is_stationary_16 <= io_in_c_bypass_13_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_1_data_16 <= io_in_c_bypass_13_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_1_is_stationary_16 <= io_in_c_bypass_13_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_2_data_16 <= io_in_c_bypass_13_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_2_is_stationary_16 <= io_in_c_bypass_13_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_3_data_16 <= io_in_c_bypass_13_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_3_is_stationary_16 <= io_in_c_bypass_13_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_0_data_16 <= io_in_c_bypass_14_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_0_is_stationary_16 <= io_in_c_bypass_14_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_1_data_16 <= io_in_c_bypass_14_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_1_is_stationary_16 <= io_in_c_bypass_14_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_2_data_16 <= io_in_c_bypass_14_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_2_is_stationary_16 <= io_in_c_bypass_14_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_3_data_16 <= io_in_c_bypass_14_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_3_is_stationary_16 <= io_in_c_bypass_14_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_0_data_16 <= io_in_c_bypass_15_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_0_is_stationary_16 <= io_in_c_bypass_15_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_1_data_16 <= io_in_c_bypass_15_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_1_is_stationary_16 <= io_in_c_bypass_15_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_2_data_16 <= io_in_c_bypass_15_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_2_is_stationary_16 <= io_in_c_bypass_15_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_3_data_16 <= io_in_c_bypass_15_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_3_is_stationary_16 <= io_in_c_bypass_15_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_0_data_16 <= io_in_c_bypass_16_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_0_is_stationary_16 <= io_in_c_bypass_16_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_1_data_16 <= io_in_c_bypass_16_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_1_is_stationary_16 <= io_in_c_bypass_16_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_2_data_16 <= io_in_c_bypass_16_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_2_is_stationary_16 <= io_in_c_bypass_16_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_3_data_16 <= io_in_c_bypass_16_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_3_is_stationary_16 <= io_in_c_bypass_16_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_0_data_16 <= io_in_c_bypass_17_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_0_is_stationary_16 <= io_in_c_bypass_17_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_1_data_16 <= io_in_c_bypass_17_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_1_is_stationary_16 <= io_in_c_bypass_17_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_2_data_16 <= io_in_c_bypass_17_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_2_is_stationary_16 <= io_in_c_bypass_17_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_3_data_16 <= io_in_c_bypass_17_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_3_is_stationary_16 <= io_in_c_bypass_17_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_0_data_16 <= io_in_c_bypass_18_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_0_is_stationary_16 <= io_in_c_bypass_18_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_1_data_16 <= io_in_c_bypass_18_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_1_is_stationary_16 <= io_in_c_bypass_18_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_2_data_16 <= io_in_c_bypass_18_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_2_is_stationary_16 <= io_in_c_bypass_18_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_3_data_16 <= io_in_c_bypass_18_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_3_is_stationary_16 <= io_in_c_bypass_18_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_0_data_16 <= io_in_c_bypass_19_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_0_is_stationary_16 <= io_in_c_bypass_19_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_1_data_16 <= io_in_c_bypass_19_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_1_is_stationary_16 <= io_in_c_bypass_19_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_2_data_16 <= io_in_c_bypass_19_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_2_is_stationary_16 <= io_in_c_bypass_19_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_3_data_16 <= io_in_c_bypass_19_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_3_is_stationary_16 <= io_in_c_bypass_19_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_0_data_16 <= io_in_c_bypass_20_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_0_is_stationary_16 <= io_in_c_bypass_20_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_1_data_16 <= io_in_c_bypass_20_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_1_is_stationary_16 <= io_in_c_bypass_20_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_2_data_16 <= io_in_c_bypass_20_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_2_is_stationary_16 <= io_in_c_bypass_20_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_3_data_16 <= io_in_c_bypass_20_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_3_is_stationary_16 <= io_in_c_bypass_20_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_0_data_16 <= io_in_c_bypass_21_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_0_is_stationary_16 <= io_in_c_bypass_21_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_1_data_16 <= io_in_c_bypass_21_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_1_is_stationary_16 <= io_in_c_bypass_21_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_2_data_16 <= io_in_c_bypass_21_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_2_is_stationary_16 <= io_in_c_bypass_21_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_3_data_16 <= io_in_c_bypass_21_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_3_is_stationary_16 <= io_in_c_bypass_21_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_0_data_16 <= io_in_c_bypass_22_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_0_is_stationary_16 <= io_in_c_bypass_22_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_1_data_16 <= io_in_c_bypass_22_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_1_is_stationary_16 <= io_in_c_bypass_22_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_2_data_16 <= io_in_c_bypass_22_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_2_is_stationary_16 <= io_in_c_bypass_22_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_3_data_16 <= io_in_c_bypass_22_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_3_is_stationary_16 <= io_in_c_bypass_22_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_0_data_16 <= io_in_c_bypass_23_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_0_is_stationary_16 <= io_in_c_bypass_23_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_1_data_16 <= io_in_c_bypass_23_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_1_is_stationary_16 <= io_in_c_bypass_23_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_2_data_16 <= io_in_c_bypass_23_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_2_is_stationary_16 <= io_in_c_bypass_23_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_3_data_16 <= io_in_c_bypass_23_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_3_is_stationary_16 <= io_in_c_bypass_23_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_0_data_16 <= io_in_c_bypass_24_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_0_is_stationary_16 <= io_in_c_bypass_24_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_1_data_16 <= io_in_c_bypass_24_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_1_is_stationary_16 <= io_in_c_bypass_24_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_2_data_16 <= io_in_c_bypass_24_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_2_is_stationary_16 <= io_in_c_bypass_24_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_3_data_16 <= io_in_c_bypass_24_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_3_is_stationary_16 <= io_in_c_bypass_24_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_0_data_16 <= io_in_c_bypass_25_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_0_is_stationary_16 <= io_in_c_bypass_25_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_1_data_16 <= io_in_c_bypass_25_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_1_is_stationary_16 <= io_in_c_bypass_25_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_2_data_16 <= io_in_c_bypass_25_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_2_is_stationary_16 <= io_in_c_bypass_25_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_3_data_16 <= io_in_c_bypass_25_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_3_is_stationary_16 <= io_in_c_bypass_25_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_0_data_16 <= io_in_c_bypass_26_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_0_is_stationary_16 <= io_in_c_bypass_26_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_1_data_16 <= io_in_c_bypass_26_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_1_is_stationary_16 <= io_in_c_bypass_26_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_2_data_16 <= io_in_c_bypass_26_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_2_is_stationary_16 <= io_in_c_bypass_26_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_3_data_16 <= io_in_c_bypass_26_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_3_is_stationary_16 <= io_in_c_bypass_26_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_0_data_16 <= io_in_c_bypass_27_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_0_is_stationary_16 <= io_in_c_bypass_27_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_1_data_16 <= io_in_c_bypass_27_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_1_is_stationary_16 <= io_in_c_bypass_27_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_2_data_16 <= io_in_c_bypass_27_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_2_is_stationary_16 <= io_in_c_bypass_27_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_3_data_16 <= io_in_c_bypass_27_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_3_is_stationary_16 <= io_in_c_bypass_27_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_0_data_16 <= io_in_c_bypass_28_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_0_is_stationary_16 <= io_in_c_bypass_28_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_1_data_16 <= io_in_c_bypass_28_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_1_is_stationary_16 <= io_in_c_bypass_28_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_2_data_16 <= io_in_c_bypass_28_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_2_is_stationary_16 <= io_in_c_bypass_28_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_3_data_16 <= io_in_c_bypass_28_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_3_is_stationary_16 <= io_in_c_bypass_28_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_0_data_16 <= io_in_c_bypass_29_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_0_is_stationary_16 <= io_in_c_bypass_29_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_1_data_16 <= io_in_c_bypass_29_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_1_is_stationary_16 <= io_in_c_bypass_29_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_2_data_16 <= io_in_c_bypass_29_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_2_is_stationary_16 <= io_in_c_bypass_29_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_3_data_16 <= io_in_c_bypass_29_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_3_is_stationary_16 <= io_in_c_bypass_29_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_0_data_16 <= io_in_c_bypass_30_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_0_is_stationary_16 <= io_in_c_bypass_30_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_1_data_16 <= io_in_c_bypass_30_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_1_is_stationary_16 <= io_in_c_bypass_30_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_2_data_16 <= io_in_c_bypass_30_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_2_is_stationary_16 <= io_in_c_bypass_30_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_3_data_16 <= io_in_c_bypass_30_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_3_is_stationary_16 <= io_in_c_bypass_30_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_0_data_16 <= io_in_c_bypass_31_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_0_is_stationary_16 <= io_in_c_bypass_31_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_1_data_16 <= io_in_c_bypass_31_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_1_is_stationary_16 <= io_in_c_bypass_31_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_2_data_16 <= io_in_c_bypass_31_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_2_is_stationary_16 <= io_in_c_bypass_31_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_3_data_16 <= io_in_c_bypass_31_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_3_is_stationary_16 <= io_in_c_bypass_31_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_0_data_17 <= io_in_c_bypass_0_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_0_is_stationary_17 <= io_in_c_bypass_0_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_1_data_17 <= io_in_c_bypass_0_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_1_is_stationary_17 <= io_in_c_bypass_0_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_2_data_17 <= io_in_c_bypass_0_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_2_is_stationary_17 <= io_in_c_bypass_0_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_3_data_17 <= io_in_c_bypass_0_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_3_is_stationary_17 <= io_in_c_bypass_0_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_0_data_17 <= io_in_c_bypass_1_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_0_is_stationary_17 <= io_in_c_bypass_1_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_1_data_17 <= io_in_c_bypass_1_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_1_is_stationary_17 <= io_in_c_bypass_1_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_2_data_17 <= io_in_c_bypass_1_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_2_is_stationary_17 <= io_in_c_bypass_1_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_3_data_17 <= io_in_c_bypass_1_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_3_is_stationary_17 <= io_in_c_bypass_1_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_0_data_17 <= io_in_c_bypass_2_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_0_is_stationary_17 <= io_in_c_bypass_2_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_1_data_17 <= io_in_c_bypass_2_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_1_is_stationary_17 <= io_in_c_bypass_2_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_2_data_17 <= io_in_c_bypass_2_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_2_is_stationary_17 <= io_in_c_bypass_2_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_3_data_17 <= io_in_c_bypass_2_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_3_is_stationary_17 <= io_in_c_bypass_2_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_0_data_17 <= io_in_c_bypass_3_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_0_is_stationary_17 <= io_in_c_bypass_3_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_1_data_17 <= io_in_c_bypass_3_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_1_is_stationary_17 <= io_in_c_bypass_3_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_2_data_17 <= io_in_c_bypass_3_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_2_is_stationary_17 <= io_in_c_bypass_3_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_3_data_17 <= io_in_c_bypass_3_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_3_is_stationary_17 <= io_in_c_bypass_3_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_0_data_17 <= io_in_c_bypass_4_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_0_is_stationary_17 <= io_in_c_bypass_4_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_1_data_17 <= io_in_c_bypass_4_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_1_is_stationary_17 <= io_in_c_bypass_4_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_2_data_17 <= io_in_c_bypass_4_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_2_is_stationary_17 <= io_in_c_bypass_4_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_3_data_17 <= io_in_c_bypass_4_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_3_is_stationary_17 <= io_in_c_bypass_4_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_0_data_17 <= io_in_c_bypass_5_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_0_is_stationary_17 <= io_in_c_bypass_5_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_1_data_17 <= io_in_c_bypass_5_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_1_is_stationary_17 <= io_in_c_bypass_5_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_2_data_17 <= io_in_c_bypass_5_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_2_is_stationary_17 <= io_in_c_bypass_5_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_3_data_17 <= io_in_c_bypass_5_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_3_is_stationary_17 <= io_in_c_bypass_5_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_0_data_17 <= io_in_c_bypass_6_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_0_is_stationary_17 <= io_in_c_bypass_6_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_1_data_17 <= io_in_c_bypass_6_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_1_is_stationary_17 <= io_in_c_bypass_6_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_2_data_17 <= io_in_c_bypass_6_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_2_is_stationary_17 <= io_in_c_bypass_6_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_3_data_17 <= io_in_c_bypass_6_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_3_is_stationary_17 <= io_in_c_bypass_6_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_0_data_17 <= io_in_c_bypass_7_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_0_is_stationary_17 <= io_in_c_bypass_7_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_1_data_17 <= io_in_c_bypass_7_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_1_is_stationary_17 <= io_in_c_bypass_7_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_2_data_17 <= io_in_c_bypass_7_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_2_is_stationary_17 <= io_in_c_bypass_7_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_3_data_17 <= io_in_c_bypass_7_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_3_is_stationary_17 <= io_in_c_bypass_7_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_0_data_17 <= io_in_c_bypass_8_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_0_is_stationary_17 <= io_in_c_bypass_8_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_1_data_17 <= io_in_c_bypass_8_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_1_is_stationary_17 <= io_in_c_bypass_8_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_2_data_17 <= io_in_c_bypass_8_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_2_is_stationary_17 <= io_in_c_bypass_8_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_3_data_17 <= io_in_c_bypass_8_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_3_is_stationary_17 <= io_in_c_bypass_8_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_0_data_17 <= io_in_c_bypass_9_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_0_is_stationary_17 <= io_in_c_bypass_9_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_1_data_17 <= io_in_c_bypass_9_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_1_is_stationary_17 <= io_in_c_bypass_9_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_2_data_17 <= io_in_c_bypass_9_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_2_is_stationary_17 <= io_in_c_bypass_9_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_3_data_17 <= io_in_c_bypass_9_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_3_is_stationary_17 <= io_in_c_bypass_9_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_0_data_17 <= io_in_c_bypass_10_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_0_is_stationary_17 <= io_in_c_bypass_10_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_1_data_17 <= io_in_c_bypass_10_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_1_is_stationary_17 <= io_in_c_bypass_10_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_2_data_17 <= io_in_c_bypass_10_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_2_is_stationary_17 <= io_in_c_bypass_10_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_3_data_17 <= io_in_c_bypass_10_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_3_is_stationary_17 <= io_in_c_bypass_10_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_0_data_17 <= io_in_c_bypass_11_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_0_is_stationary_17 <= io_in_c_bypass_11_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_1_data_17 <= io_in_c_bypass_11_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_1_is_stationary_17 <= io_in_c_bypass_11_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_2_data_17 <= io_in_c_bypass_11_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_2_is_stationary_17 <= io_in_c_bypass_11_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_3_data_17 <= io_in_c_bypass_11_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_3_is_stationary_17 <= io_in_c_bypass_11_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_0_data_17 <= io_in_c_bypass_12_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_0_is_stationary_17 <= io_in_c_bypass_12_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_1_data_17 <= io_in_c_bypass_12_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_1_is_stationary_17 <= io_in_c_bypass_12_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_2_data_17 <= io_in_c_bypass_12_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_2_is_stationary_17 <= io_in_c_bypass_12_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_3_data_17 <= io_in_c_bypass_12_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_3_is_stationary_17 <= io_in_c_bypass_12_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_0_data_17 <= io_in_c_bypass_13_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_0_is_stationary_17 <= io_in_c_bypass_13_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_1_data_17 <= io_in_c_bypass_13_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_1_is_stationary_17 <= io_in_c_bypass_13_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_2_data_17 <= io_in_c_bypass_13_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_2_is_stationary_17 <= io_in_c_bypass_13_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_3_data_17 <= io_in_c_bypass_13_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_3_is_stationary_17 <= io_in_c_bypass_13_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_0_data_17 <= io_in_c_bypass_14_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_0_is_stationary_17 <= io_in_c_bypass_14_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_1_data_17 <= io_in_c_bypass_14_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_1_is_stationary_17 <= io_in_c_bypass_14_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_2_data_17 <= io_in_c_bypass_14_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_2_is_stationary_17 <= io_in_c_bypass_14_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_3_data_17 <= io_in_c_bypass_14_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_3_is_stationary_17 <= io_in_c_bypass_14_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_0_data_17 <= io_in_c_bypass_15_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_0_is_stationary_17 <= io_in_c_bypass_15_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_1_data_17 <= io_in_c_bypass_15_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_1_is_stationary_17 <= io_in_c_bypass_15_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_2_data_17 <= io_in_c_bypass_15_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_2_is_stationary_17 <= io_in_c_bypass_15_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_3_data_17 <= io_in_c_bypass_15_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_3_is_stationary_17 <= io_in_c_bypass_15_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_0_data_17 <= io_in_c_bypass_16_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_0_is_stationary_17 <= io_in_c_bypass_16_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_1_data_17 <= io_in_c_bypass_16_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_1_is_stationary_17 <= io_in_c_bypass_16_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_2_data_17 <= io_in_c_bypass_16_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_2_is_stationary_17 <= io_in_c_bypass_16_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_3_data_17 <= io_in_c_bypass_16_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_3_is_stationary_17 <= io_in_c_bypass_16_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_0_data_17 <= io_in_c_bypass_17_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_0_is_stationary_17 <= io_in_c_bypass_17_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_1_data_17 <= io_in_c_bypass_17_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_1_is_stationary_17 <= io_in_c_bypass_17_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_2_data_17 <= io_in_c_bypass_17_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_2_is_stationary_17 <= io_in_c_bypass_17_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_3_data_17 <= io_in_c_bypass_17_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_3_is_stationary_17 <= io_in_c_bypass_17_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_0_data_17 <= io_in_c_bypass_18_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_0_is_stationary_17 <= io_in_c_bypass_18_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_1_data_17 <= io_in_c_bypass_18_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_1_is_stationary_17 <= io_in_c_bypass_18_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_2_data_17 <= io_in_c_bypass_18_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_2_is_stationary_17 <= io_in_c_bypass_18_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_3_data_17 <= io_in_c_bypass_18_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_3_is_stationary_17 <= io_in_c_bypass_18_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_0_data_17 <= io_in_c_bypass_19_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_0_is_stationary_17 <= io_in_c_bypass_19_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_1_data_17 <= io_in_c_bypass_19_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_1_is_stationary_17 <= io_in_c_bypass_19_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_2_data_17 <= io_in_c_bypass_19_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_2_is_stationary_17 <= io_in_c_bypass_19_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_3_data_17 <= io_in_c_bypass_19_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_3_is_stationary_17 <= io_in_c_bypass_19_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_0_data_17 <= io_in_c_bypass_20_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_0_is_stationary_17 <= io_in_c_bypass_20_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_1_data_17 <= io_in_c_bypass_20_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_1_is_stationary_17 <= io_in_c_bypass_20_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_2_data_17 <= io_in_c_bypass_20_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_2_is_stationary_17 <= io_in_c_bypass_20_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_3_data_17 <= io_in_c_bypass_20_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_3_is_stationary_17 <= io_in_c_bypass_20_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_0_data_17 <= io_in_c_bypass_21_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_0_is_stationary_17 <= io_in_c_bypass_21_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_1_data_17 <= io_in_c_bypass_21_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_1_is_stationary_17 <= io_in_c_bypass_21_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_2_data_17 <= io_in_c_bypass_21_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_2_is_stationary_17 <= io_in_c_bypass_21_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_3_data_17 <= io_in_c_bypass_21_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_3_is_stationary_17 <= io_in_c_bypass_21_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_0_data_17 <= io_in_c_bypass_22_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_0_is_stationary_17 <= io_in_c_bypass_22_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_1_data_17 <= io_in_c_bypass_22_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_1_is_stationary_17 <= io_in_c_bypass_22_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_2_data_17 <= io_in_c_bypass_22_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_2_is_stationary_17 <= io_in_c_bypass_22_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_3_data_17 <= io_in_c_bypass_22_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_3_is_stationary_17 <= io_in_c_bypass_22_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_0_data_17 <= io_in_c_bypass_23_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_0_is_stationary_17 <= io_in_c_bypass_23_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_1_data_17 <= io_in_c_bypass_23_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_1_is_stationary_17 <= io_in_c_bypass_23_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_2_data_17 <= io_in_c_bypass_23_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_2_is_stationary_17 <= io_in_c_bypass_23_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_3_data_17 <= io_in_c_bypass_23_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_3_is_stationary_17 <= io_in_c_bypass_23_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_0_data_17 <= io_in_c_bypass_24_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_0_is_stationary_17 <= io_in_c_bypass_24_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_1_data_17 <= io_in_c_bypass_24_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_1_is_stationary_17 <= io_in_c_bypass_24_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_2_data_17 <= io_in_c_bypass_24_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_2_is_stationary_17 <= io_in_c_bypass_24_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_3_data_17 <= io_in_c_bypass_24_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_3_is_stationary_17 <= io_in_c_bypass_24_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_0_data_17 <= io_in_c_bypass_25_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_0_is_stationary_17 <= io_in_c_bypass_25_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_1_data_17 <= io_in_c_bypass_25_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_1_is_stationary_17 <= io_in_c_bypass_25_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_2_data_17 <= io_in_c_bypass_25_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_2_is_stationary_17 <= io_in_c_bypass_25_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_3_data_17 <= io_in_c_bypass_25_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_3_is_stationary_17 <= io_in_c_bypass_25_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_0_data_17 <= io_in_c_bypass_26_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_0_is_stationary_17 <= io_in_c_bypass_26_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_1_data_17 <= io_in_c_bypass_26_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_1_is_stationary_17 <= io_in_c_bypass_26_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_2_data_17 <= io_in_c_bypass_26_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_2_is_stationary_17 <= io_in_c_bypass_26_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_3_data_17 <= io_in_c_bypass_26_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_3_is_stationary_17 <= io_in_c_bypass_26_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_0_data_17 <= io_in_c_bypass_27_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_0_is_stationary_17 <= io_in_c_bypass_27_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_1_data_17 <= io_in_c_bypass_27_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_1_is_stationary_17 <= io_in_c_bypass_27_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_2_data_17 <= io_in_c_bypass_27_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_2_is_stationary_17 <= io_in_c_bypass_27_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_3_data_17 <= io_in_c_bypass_27_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_3_is_stationary_17 <= io_in_c_bypass_27_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_0_data_17 <= io_in_c_bypass_28_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_0_is_stationary_17 <= io_in_c_bypass_28_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_1_data_17 <= io_in_c_bypass_28_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_1_is_stationary_17 <= io_in_c_bypass_28_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_2_data_17 <= io_in_c_bypass_28_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_2_is_stationary_17 <= io_in_c_bypass_28_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_3_data_17 <= io_in_c_bypass_28_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_3_is_stationary_17 <= io_in_c_bypass_28_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_0_data_17 <= io_in_c_bypass_29_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_0_is_stationary_17 <= io_in_c_bypass_29_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_1_data_17 <= io_in_c_bypass_29_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_1_is_stationary_17 <= io_in_c_bypass_29_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_2_data_17 <= io_in_c_bypass_29_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_2_is_stationary_17 <= io_in_c_bypass_29_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_3_data_17 <= io_in_c_bypass_29_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_3_is_stationary_17 <= io_in_c_bypass_29_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_0_data_17 <= io_in_c_bypass_30_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_0_is_stationary_17 <= io_in_c_bypass_30_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_1_data_17 <= io_in_c_bypass_30_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_1_is_stationary_17 <= io_in_c_bypass_30_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_2_data_17 <= io_in_c_bypass_30_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_2_is_stationary_17 <= io_in_c_bypass_30_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_3_data_17 <= io_in_c_bypass_30_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_3_is_stationary_17 <= io_in_c_bypass_30_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_0_data_17 <= io_in_c_bypass_31_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_0_is_stationary_17 <= io_in_c_bypass_31_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_1_data_17 <= io_in_c_bypass_31_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_1_is_stationary_17 <= io_in_c_bypass_31_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_2_data_17 <= io_in_c_bypass_31_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_2_is_stationary_17 <= io_in_c_bypass_31_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_3_data_17 <= io_in_c_bypass_31_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_3_is_stationary_17 <= io_in_c_bypass_31_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_0_data_18 <= io_in_c_bypass_0_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_0_is_stationary_18 <= io_in_c_bypass_0_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_1_data_18 <= io_in_c_bypass_0_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_1_is_stationary_18 <= io_in_c_bypass_0_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_2_data_18 <= io_in_c_bypass_0_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_2_is_stationary_18 <= io_in_c_bypass_0_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_3_data_18 <= io_in_c_bypass_0_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_3_is_stationary_18 <= io_in_c_bypass_0_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_0_data_18 <= io_in_c_bypass_1_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_0_is_stationary_18 <= io_in_c_bypass_1_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_1_data_18 <= io_in_c_bypass_1_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_1_is_stationary_18 <= io_in_c_bypass_1_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_2_data_18 <= io_in_c_bypass_1_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_2_is_stationary_18 <= io_in_c_bypass_1_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_3_data_18 <= io_in_c_bypass_1_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_3_is_stationary_18 <= io_in_c_bypass_1_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_0_data_18 <= io_in_c_bypass_2_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_0_is_stationary_18 <= io_in_c_bypass_2_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_1_data_18 <= io_in_c_bypass_2_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_1_is_stationary_18 <= io_in_c_bypass_2_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_2_data_18 <= io_in_c_bypass_2_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_2_is_stationary_18 <= io_in_c_bypass_2_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_3_data_18 <= io_in_c_bypass_2_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_3_is_stationary_18 <= io_in_c_bypass_2_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_0_data_18 <= io_in_c_bypass_3_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_0_is_stationary_18 <= io_in_c_bypass_3_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_1_data_18 <= io_in_c_bypass_3_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_1_is_stationary_18 <= io_in_c_bypass_3_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_2_data_18 <= io_in_c_bypass_3_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_2_is_stationary_18 <= io_in_c_bypass_3_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_3_data_18 <= io_in_c_bypass_3_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_3_is_stationary_18 <= io_in_c_bypass_3_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_0_data_18 <= io_in_c_bypass_4_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_0_is_stationary_18 <= io_in_c_bypass_4_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_1_data_18 <= io_in_c_bypass_4_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_1_is_stationary_18 <= io_in_c_bypass_4_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_2_data_18 <= io_in_c_bypass_4_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_2_is_stationary_18 <= io_in_c_bypass_4_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_3_data_18 <= io_in_c_bypass_4_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_3_is_stationary_18 <= io_in_c_bypass_4_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_0_data_18 <= io_in_c_bypass_5_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_0_is_stationary_18 <= io_in_c_bypass_5_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_1_data_18 <= io_in_c_bypass_5_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_1_is_stationary_18 <= io_in_c_bypass_5_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_2_data_18 <= io_in_c_bypass_5_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_2_is_stationary_18 <= io_in_c_bypass_5_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_3_data_18 <= io_in_c_bypass_5_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_3_is_stationary_18 <= io_in_c_bypass_5_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_0_data_18 <= io_in_c_bypass_6_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_0_is_stationary_18 <= io_in_c_bypass_6_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_1_data_18 <= io_in_c_bypass_6_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_1_is_stationary_18 <= io_in_c_bypass_6_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_2_data_18 <= io_in_c_bypass_6_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_2_is_stationary_18 <= io_in_c_bypass_6_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_3_data_18 <= io_in_c_bypass_6_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_3_is_stationary_18 <= io_in_c_bypass_6_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_0_data_18 <= io_in_c_bypass_7_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_0_is_stationary_18 <= io_in_c_bypass_7_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_1_data_18 <= io_in_c_bypass_7_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_1_is_stationary_18 <= io_in_c_bypass_7_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_2_data_18 <= io_in_c_bypass_7_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_2_is_stationary_18 <= io_in_c_bypass_7_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_3_data_18 <= io_in_c_bypass_7_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_3_is_stationary_18 <= io_in_c_bypass_7_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_0_data_18 <= io_in_c_bypass_8_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_0_is_stationary_18 <= io_in_c_bypass_8_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_1_data_18 <= io_in_c_bypass_8_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_1_is_stationary_18 <= io_in_c_bypass_8_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_2_data_18 <= io_in_c_bypass_8_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_2_is_stationary_18 <= io_in_c_bypass_8_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_3_data_18 <= io_in_c_bypass_8_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_3_is_stationary_18 <= io_in_c_bypass_8_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_0_data_18 <= io_in_c_bypass_9_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_0_is_stationary_18 <= io_in_c_bypass_9_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_1_data_18 <= io_in_c_bypass_9_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_1_is_stationary_18 <= io_in_c_bypass_9_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_2_data_18 <= io_in_c_bypass_9_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_2_is_stationary_18 <= io_in_c_bypass_9_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_3_data_18 <= io_in_c_bypass_9_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_3_is_stationary_18 <= io_in_c_bypass_9_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_0_data_18 <= io_in_c_bypass_10_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_0_is_stationary_18 <= io_in_c_bypass_10_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_1_data_18 <= io_in_c_bypass_10_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_1_is_stationary_18 <= io_in_c_bypass_10_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_2_data_18 <= io_in_c_bypass_10_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_2_is_stationary_18 <= io_in_c_bypass_10_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_3_data_18 <= io_in_c_bypass_10_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_3_is_stationary_18 <= io_in_c_bypass_10_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_0_data_18 <= io_in_c_bypass_11_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_0_is_stationary_18 <= io_in_c_bypass_11_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_1_data_18 <= io_in_c_bypass_11_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_1_is_stationary_18 <= io_in_c_bypass_11_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_2_data_18 <= io_in_c_bypass_11_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_2_is_stationary_18 <= io_in_c_bypass_11_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_3_data_18 <= io_in_c_bypass_11_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_3_is_stationary_18 <= io_in_c_bypass_11_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_0_data_18 <= io_in_c_bypass_12_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_0_is_stationary_18 <= io_in_c_bypass_12_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_1_data_18 <= io_in_c_bypass_12_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_1_is_stationary_18 <= io_in_c_bypass_12_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_2_data_18 <= io_in_c_bypass_12_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_2_is_stationary_18 <= io_in_c_bypass_12_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_3_data_18 <= io_in_c_bypass_12_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_3_is_stationary_18 <= io_in_c_bypass_12_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_0_data_18 <= io_in_c_bypass_13_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_0_is_stationary_18 <= io_in_c_bypass_13_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_1_data_18 <= io_in_c_bypass_13_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_1_is_stationary_18 <= io_in_c_bypass_13_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_2_data_18 <= io_in_c_bypass_13_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_2_is_stationary_18 <= io_in_c_bypass_13_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_3_data_18 <= io_in_c_bypass_13_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_3_is_stationary_18 <= io_in_c_bypass_13_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_0_data_18 <= io_in_c_bypass_14_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_0_is_stationary_18 <= io_in_c_bypass_14_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_1_data_18 <= io_in_c_bypass_14_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_1_is_stationary_18 <= io_in_c_bypass_14_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_2_data_18 <= io_in_c_bypass_14_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_2_is_stationary_18 <= io_in_c_bypass_14_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_3_data_18 <= io_in_c_bypass_14_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_3_is_stationary_18 <= io_in_c_bypass_14_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_0_data_18 <= io_in_c_bypass_15_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_0_is_stationary_18 <= io_in_c_bypass_15_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_1_data_18 <= io_in_c_bypass_15_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_1_is_stationary_18 <= io_in_c_bypass_15_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_2_data_18 <= io_in_c_bypass_15_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_2_is_stationary_18 <= io_in_c_bypass_15_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_3_data_18 <= io_in_c_bypass_15_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_3_is_stationary_18 <= io_in_c_bypass_15_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_0_data_18 <= io_in_c_bypass_16_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_0_is_stationary_18 <= io_in_c_bypass_16_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_1_data_18 <= io_in_c_bypass_16_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_1_is_stationary_18 <= io_in_c_bypass_16_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_2_data_18 <= io_in_c_bypass_16_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_2_is_stationary_18 <= io_in_c_bypass_16_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_3_data_18 <= io_in_c_bypass_16_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_3_is_stationary_18 <= io_in_c_bypass_16_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_0_data_18 <= io_in_c_bypass_17_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_0_is_stationary_18 <= io_in_c_bypass_17_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_1_data_18 <= io_in_c_bypass_17_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_1_is_stationary_18 <= io_in_c_bypass_17_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_2_data_18 <= io_in_c_bypass_17_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_2_is_stationary_18 <= io_in_c_bypass_17_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_3_data_18 <= io_in_c_bypass_17_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_3_is_stationary_18 <= io_in_c_bypass_17_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_0_data_18 <= io_in_c_bypass_18_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_0_is_stationary_18 <= io_in_c_bypass_18_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_1_data_18 <= io_in_c_bypass_18_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_1_is_stationary_18 <= io_in_c_bypass_18_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_2_data_18 <= io_in_c_bypass_18_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_2_is_stationary_18 <= io_in_c_bypass_18_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_3_data_18 <= io_in_c_bypass_18_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_3_is_stationary_18 <= io_in_c_bypass_18_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_0_data_18 <= io_in_c_bypass_19_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_0_is_stationary_18 <= io_in_c_bypass_19_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_1_data_18 <= io_in_c_bypass_19_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_1_is_stationary_18 <= io_in_c_bypass_19_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_2_data_18 <= io_in_c_bypass_19_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_2_is_stationary_18 <= io_in_c_bypass_19_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_3_data_18 <= io_in_c_bypass_19_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_3_is_stationary_18 <= io_in_c_bypass_19_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_0_data_18 <= io_in_c_bypass_20_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_0_is_stationary_18 <= io_in_c_bypass_20_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_1_data_18 <= io_in_c_bypass_20_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_1_is_stationary_18 <= io_in_c_bypass_20_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_2_data_18 <= io_in_c_bypass_20_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_2_is_stationary_18 <= io_in_c_bypass_20_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_3_data_18 <= io_in_c_bypass_20_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_3_is_stationary_18 <= io_in_c_bypass_20_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_0_data_18 <= io_in_c_bypass_21_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_0_is_stationary_18 <= io_in_c_bypass_21_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_1_data_18 <= io_in_c_bypass_21_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_1_is_stationary_18 <= io_in_c_bypass_21_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_2_data_18 <= io_in_c_bypass_21_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_2_is_stationary_18 <= io_in_c_bypass_21_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_3_data_18 <= io_in_c_bypass_21_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_3_is_stationary_18 <= io_in_c_bypass_21_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_0_data_18 <= io_in_c_bypass_22_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_0_is_stationary_18 <= io_in_c_bypass_22_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_1_data_18 <= io_in_c_bypass_22_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_1_is_stationary_18 <= io_in_c_bypass_22_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_2_data_18 <= io_in_c_bypass_22_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_2_is_stationary_18 <= io_in_c_bypass_22_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_3_data_18 <= io_in_c_bypass_22_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_3_is_stationary_18 <= io_in_c_bypass_22_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_0_data_18 <= io_in_c_bypass_23_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_0_is_stationary_18 <= io_in_c_bypass_23_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_1_data_18 <= io_in_c_bypass_23_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_1_is_stationary_18 <= io_in_c_bypass_23_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_2_data_18 <= io_in_c_bypass_23_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_2_is_stationary_18 <= io_in_c_bypass_23_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_3_data_18 <= io_in_c_bypass_23_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_3_is_stationary_18 <= io_in_c_bypass_23_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_0_data_18 <= io_in_c_bypass_24_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_0_is_stationary_18 <= io_in_c_bypass_24_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_1_data_18 <= io_in_c_bypass_24_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_1_is_stationary_18 <= io_in_c_bypass_24_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_2_data_18 <= io_in_c_bypass_24_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_2_is_stationary_18 <= io_in_c_bypass_24_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_3_data_18 <= io_in_c_bypass_24_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_3_is_stationary_18 <= io_in_c_bypass_24_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_0_data_18 <= io_in_c_bypass_25_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_0_is_stationary_18 <= io_in_c_bypass_25_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_1_data_18 <= io_in_c_bypass_25_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_1_is_stationary_18 <= io_in_c_bypass_25_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_2_data_18 <= io_in_c_bypass_25_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_2_is_stationary_18 <= io_in_c_bypass_25_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_3_data_18 <= io_in_c_bypass_25_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_3_is_stationary_18 <= io_in_c_bypass_25_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_0_data_18 <= io_in_c_bypass_26_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_0_is_stationary_18 <= io_in_c_bypass_26_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_1_data_18 <= io_in_c_bypass_26_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_1_is_stationary_18 <= io_in_c_bypass_26_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_2_data_18 <= io_in_c_bypass_26_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_2_is_stationary_18 <= io_in_c_bypass_26_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_3_data_18 <= io_in_c_bypass_26_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_3_is_stationary_18 <= io_in_c_bypass_26_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_0_data_18 <= io_in_c_bypass_27_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_0_is_stationary_18 <= io_in_c_bypass_27_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_1_data_18 <= io_in_c_bypass_27_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_1_is_stationary_18 <= io_in_c_bypass_27_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_2_data_18 <= io_in_c_bypass_27_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_2_is_stationary_18 <= io_in_c_bypass_27_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_3_data_18 <= io_in_c_bypass_27_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_3_is_stationary_18 <= io_in_c_bypass_27_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_0_data_18 <= io_in_c_bypass_28_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_0_is_stationary_18 <= io_in_c_bypass_28_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_1_data_18 <= io_in_c_bypass_28_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_1_is_stationary_18 <= io_in_c_bypass_28_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_2_data_18 <= io_in_c_bypass_28_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_2_is_stationary_18 <= io_in_c_bypass_28_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_3_data_18 <= io_in_c_bypass_28_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_3_is_stationary_18 <= io_in_c_bypass_28_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_0_data_18 <= io_in_c_bypass_29_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_0_is_stationary_18 <= io_in_c_bypass_29_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_1_data_18 <= io_in_c_bypass_29_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_1_is_stationary_18 <= io_in_c_bypass_29_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_2_data_18 <= io_in_c_bypass_29_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_2_is_stationary_18 <= io_in_c_bypass_29_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_3_data_18 <= io_in_c_bypass_29_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_3_is_stationary_18 <= io_in_c_bypass_29_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_0_data_18 <= io_in_c_bypass_30_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_0_is_stationary_18 <= io_in_c_bypass_30_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_1_data_18 <= io_in_c_bypass_30_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_1_is_stationary_18 <= io_in_c_bypass_30_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_2_data_18 <= io_in_c_bypass_30_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_2_is_stationary_18 <= io_in_c_bypass_30_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_3_data_18 <= io_in_c_bypass_30_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_3_is_stationary_18 <= io_in_c_bypass_30_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_0_data_18 <= io_in_c_bypass_31_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_0_is_stationary_18 <= io_in_c_bypass_31_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_1_data_18 <= io_in_c_bypass_31_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_1_is_stationary_18 <= io_in_c_bypass_31_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_2_data_18 <= io_in_c_bypass_31_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_2_is_stationary_18 <= io_in_c_bypass_31_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_3_data_18 <= io_in_c_bypass_31_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_3_is_stationary_18 <= io_in_c_bypass_31_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_0_data_19 <= io_in_c_bypass_0_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_0_is_stationary_19 <= io_in_c_bypass_0_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_1_data_19 <= io_in_c_bypass_0_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_1_is_stationary_19 <= io_in_c_bypass_0_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_2_data_19 <= io_in_c_bypass_0_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_2_is_stationary_19 <= io_in_c_bypass_0_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_3_data_19 <= io_in_c_bypass_0_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_3_is_stationary_19 <= io_in_c_bypass_0_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_0_data_19 <= io_in_c_bypass_1_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_0_is_stationary_19 <= io_in_c_bypass_1_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_1_data_19 <= io_in_c_bypass_1_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_1_is_stationary_19 <= io_in_c_bypass_1_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_2_data_19 <= io_in_c_bypass_1_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_2_is_stationary_19 <= io_in_c_bypass_1_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_3_data_19 <= io_in_c_bypass_1_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_3_is_stationary_19 <= io_in_c_bypass_1_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_0_data_19 <= io_in_c_bypass_2_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_0_is_stationary_19 <= io_in_c_bypass_2_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_1_data_19 <= io_in_c_bypass_2_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_1_is_stationary_19 <= io_in_c_bypass_2_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_2_data_19 <= io_in_c_bypass_2_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_2_is_stationary_19 <= io_in_c_bypass_2_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_3_data_19 <= io_in_c_bypass_2_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_3_is_stationary_19 <= io_in_c_bypass_2_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_0_data_19 <= io_in_c_bypass_3_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_0_is_stationary_19 <= io_in_c_bypass_3_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_1_data_19 <= io_in_c_bypass_3_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_1_is_stationary_19 <= io_in_c_bypass_3_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_2_data_19 <= io_in_c_bypass_3_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_2_is_stationary_19 <= io_in_c_bypass_3_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_3_data_19 <= io_in_c_bypass_3_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_3_is_stationary_19 <= io_in_c_bypass_3_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_0_data_19 <= io_in_c_bypass_4_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_0_is_stationary_19 <= io_in_c_bypass_4_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_1_data_19 <= io_in_c_bypass_4_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_1_is_stationary_19 <= io_in_c_bypass_4_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_2_data_19 <= io_in_c_bypass_4_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_2_is_stationary_19 <= io_in_c_bypass_4_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_3_data_19 <= io_in_c_bypass_4_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_3_is_stationary_19 <= io_in_c_bypass_4_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_0_data_19 <= io_in_c_bypass_5_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_0_is_stationary_19 <= io_in_c_bypass_5_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_1_data_19 <= io_in_c_bypass_5_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_1_is_stationary_19 <= io_in_c_bypass_5_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_2_data_19 <= io_in_c_bypass_5_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_2_is_stationary_19 <= io_in_c_bypass_5_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_3_data_19 <= io_in_c_bypass_5_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_3_is_stationary_19 <= io_in_c_bypass_5_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_0_data_19 <= io_in_c_bypass_6_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_0_is_stationary_19 <= io_in_c_bypass_6_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_1_data_19 <= io_in_c_bypass_6_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_1_is_stationary_19 <= io_in_c_bypass_6_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_2_data_19 <= io_in_c_bypass_6_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_2_is_stationary_19 <= io_in_c_bypass_6_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_3_data_19 <= io_in_c_bypass_6_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_3_is_stationary_19 <= io_in_c_bypass_6_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_0_data_19 <= io_in_c_bypass_7_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_0_is_stationary_19 <= io_in_c_bypass_7_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_1_data_19 <= io_in_c_bypass_7_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_1_is_stationary_19 <= io_in_c_bypass_7_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_2_data_19 <= io_in_c_bypass_7_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_2_is_stationary_19 <= io_in_c_bypass_7_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_3_data_19 <= io_in_c_bypass_7_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_3_is_stationary_19 <= io_in_c_bypass_7_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_0_data_19 <= io_in_c_bypass_8_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_0_is_stationary_19 <= io_in_c_bypass_8_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_1_data_19 <= io_in_c_bypass_8_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_1_is_stationary_19 <= io_in_c_bypass_8_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_2_data_19 <= io_in_c_bypass_8_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_2_is_stationary_19 <= io_in_c_bypass_8_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_3_data_19 <= io_in_c_bypass_8_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_3_is_stationary_19 <= io_in_c_bypass_8_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_0_data_19 <= io_in_c_bypass_9_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_0_is_stationary_19 <= io_in_c_bypass_9_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_1_data_19 <= io_in_c_bypass_9_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_1_is_stationary_19 <= io_in_c_bypass_9_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_2_data_19 <= io_in_c_bypass_9_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_2_is_stationary_19 <= io_in_c_bypass_9_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_3_data_19 <= io_in_c_bypass_9_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_3_is_stationary_19 <= io_in_c_bypass_9_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_0_data_19 <= io_in_c_bypass_10_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_0_is_stationary_19 <= io_in_c_bypass_10_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_1_data_19 <= io_in_c_bypass_10_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_1_is_stationary_19 <= io_in_c_bypass_10_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_2_data_19 <= io_in_c_bypass_10_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_2_is_stationary_19 <= io_in_c_bypass_10_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_3_data_19 <= io_in_c_bypass_10_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_3_is_stationary_19 <= io_in_c_bypass_10_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_0_data_19 <= io_in_c_bypass_11_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_0_is_stationary_19 <= io_in_c_bypass_11_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_1_data_19 <= io_in_c_bypass_11_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_1_is_stationary_19 <= io_in_c_bypass_11_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_2_data_19 <= io_in_c_bypass_11_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_2_is_stationary_19 <= io_in_c_bypass_11_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_3_data_19 <= io_in_c_bypass_11_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_3_is_stationary_19 <= io_in_c_bypass_11_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_0_data_19 <= io_in_c_bypass_12_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_0_is_stationary_19 <= io_in_c_bypass_12_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_1_data_19 <= io_in_c_bypass_12_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_1_is_stationary_19 <= io_in_c_bypass_12_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_2_data_19 <= io_in_c_bypass_12_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_2_is_stationary_19 <= io_in_c_bypass_12_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_3_data_19 <= io_in_c_bypass_12_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_3_is_stationary_19 <= io_in_c_bypass_12_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_0_data_19 <= io_in_c_bypass_13_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_0_is_stationary_19 <= io_in_c_bypass_13_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_1_data_19 <= io_in_c_bypass_13_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_1_is_stationary_19 <= io_in_c_bypass_13_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_2_data_19 <= io_in_c_bypass_13_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_2_is_stationary_19 <= io_in_c_bypass_13_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_3_data_19 <= io_in_c_bypass_13_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_3_is_stationary_19 <= io_in_c_bypass_13_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_0_data_19 <= io_in_c_bypass_14_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_0_is_stationary_19 <= io_in_c_bypass_14_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_1_data_19 <= io_in_c_bypass_14_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_1_is_stationary_19 <= io_in_c_bypass_14_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_2_data_19 <= io_in_c_bypass_14_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_2_is_stationary_19 <= io_in_c_bypass_14_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_3_data_19 <= io_in_c_bypass_14_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_3_is_stationary_19 <= io_in_c_bypass_14_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_0_data_19 <= io_in_c_bypass_15_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_0_is_stationary_19 <= io_in_c_bypass_15_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_1_data_19 <= io_in_c_bypass_15_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_1_is_stationary_19 <= io_in_c_bypass_15_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_2_data_19 <= io_in_c_bypass_15_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_2_is_stationary_19 <= io_in_c_bypass_15_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_3_data_19 <= io_in_c_bypass_15_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_3_is_stationary_19 <= io_in_c_bypass_15_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_0_data_19 <= io_in_c_bypass_16_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_0_is_stationary_19 <= io_in_c_bypass_16_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_1_data_19 <= io_in_c_bypass_16_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_1_is_stationary_19 <= io_in_c_bypass_16_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_2_data_19 <= io_in_c_bypass_16_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_2_is_stationary_19 <= io_in_c_bypass_16_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_3_data_19 <= io_in_c_bypass_16_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_3_is_stationary_19 <= io_in_c_bypass_16_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_0_data_19 <= io_in_c_bypass_17_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_0_is_stationary_19 <= io_in_c_bypass_17_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_1_data_19 <= io_in_c_bypass_17_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_1_is_stationary_19 <= io_in_c_bypass_17_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_2_data_19 <= io_in_c_bypass_17_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_2_is_stationary_19 <= io_in_c_bypass_17_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_3_data_19 <= io_in_c_bypass_17_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_3_is_stationary_19 <= io_in_c_bypass_17_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_0_data_19 <= io_in_c_bypass_18_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_0_is_stationary_19 <= io_in_c_bypass_18_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_1_data_19 <= io_in_c_bypass_18_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_1_is_stationary_19 <= io_in_c_bypass_18_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_2_data_19 <= io_in_c_bypass_18_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_2_is_stationary_19 <= io_in_c_bypass_18_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_3_data_19 <= io_in_c_bypass_18_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_3_is_stationary_19 <= io_in_c_bypass_18_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_0_data_19 <= io_in_c_bypass_19_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_0_is_stationary_19 <= io_in_c_bypass_19_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_1_data_19 <= io_in_c_bypass_19_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_1_is_stationary_19 <= io_in_c_bypass_19_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_2_data_19 <= io_in_c_bypass_19_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_2_is_stationary_19 <= io_in_c_bypass_19_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_3_data_19 <= io_in_c_bypass_19_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_3_is_stationary_19 <= io_in_c_bypass_19_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_0_data_19 <= io_in_c_bypass_20_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_0_is_stationary_19 <= io_in_c_bypass_20_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_1_data_19 <= io_in_c_bypass_20_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_1_is_stationary_19 <= io_in_c_bypass_20_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_2_data_19 <= io_in_c_bypass_20_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_2_is_stationary_19 <= io_in_c_bypass_20_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_3_data_19 <= io_in_c_bypass_20_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_3_is_stationary_19 <= io_in_c_bypass_20_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_0_data_19 <= io_in_c_bypass_21_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_0_is_stationary_19 <= io_in_c_bypass_21_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_1_data_19 <= io_in_c_bypass_21_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_1_is_stationary_19 <= io_in_c_bypass_21_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_2_data_19 <= io_in_c_bypass_21_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_2_is_stationary_19 <= io_in_c_bypass_21_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_3_data_19 <= io_in_c_bypass_21_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_3_is_stationary_19 <= io_in_c_bypass_21_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_0_data_19 <= io_in_c_bypass_22_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_0_is_stationary_19 <= io_in_c_bypass_22_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_1_data_19 <= io_in_c_bypass_22_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_1_is_stationary_19 <= io_in_c_bypass_22_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_2_data_19 <= io_in_c_bypass_22_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_2_is_stationary_19 <= io_in_c_bypass_22_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_3_data_19 <= io_in_c_bypass_22_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_3_is_stationary_19 <= io_in_c_bypass_22_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_0_data_19 <= io_in_c_bypass_23_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_0_is_stationary_19 <= io_in_c_bypass_23_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_1_data_19 <= io_in_c_bypass_23_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_1_is_stationary_19 <= io_in_c_bypass_23_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_2_data_19 <= io_in_c_bypass_23_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_2_is_stationary_19 <= io_in_c_bypass_23_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_3_data_19 <= io_in_c_bypass_23_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_3_is_stationary_19 <= io_in_c_bypass_23_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_0_data_19 <= io_in_c_bypass_24_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_0_is_stationary_19 <= io_in_c_bypass_24_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_1_data_19 <= io_in_c_bypass_24_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_1_is_stationary_19 <= io_in_c_bypass_24_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_2_data_19 <= io_in_c_bypass_24_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_2_is_stationary_19 <= io_in_c_bypass_24_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_3_data_19 <= io_in_c_bypass_24_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_3_is_stationary_19 <= io_in_c_bypass_24_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_0_data_19 <= io_in_c_bypass_25_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_0_is_stationary_19 <= io_in_c_bypass_25_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_1_data_19 <= io_in_c_bypass_25_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_1_is_stationary_19 <= io_in_c_bypass_25_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_2_data_19 <= io_in_c_bypass_25_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_2_is_stationary_19 <= io_in_c_bypass_25_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_3_data_19 <= io_in_c_bypass_25_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_3_is_stationary_19 <= io_in_c_bypass_25_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_0_data_19 <= io_in_c_bypass_26_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_0_is_stationary_19 <= io_in_c_bypass_26_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_1_data_19 <= io_in_c_bypass_26_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_1_is_stationary_19 <= io_in_c_bypass_26_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_2_data_19 <= io_in_c_bypass_26_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_2_is_stationary_19 <= io_in_c_bypass_26_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_3_data_19 <= io_in_c_bypass_26_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_3_is_stationary_19 <= io_in_c_bypass_26_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_0_data_19 <= io_in_c_bypass_27_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_0_is_stationary_19 <= io_in_c_bypass_27_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_1_data_19 <= io_in_c_bypass_27_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_1_is_stationary_19 <= io_in_c_bypass_27_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_2_data_19 <= io_in_c_bypass_27_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_2_is_stationary_19 <= io_in_c_bypass_27_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_3_data_19 <= io_in_c_bypass_27_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_3_is_stationary_19 <= io_in_c_bypass_27_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_0_data_19 <= io_in_c_bypass_28_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_0_is_stationary_19 <= io_in_c_bypass_28_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_1_data_19 <= io_in_c_bypass_28_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_1_is_stationary_19 <= io_in_c_bypass_28_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_2_data_19 <= io_in_c_bypass_28_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_2_is_stationary_19 <= io_in_c_bypass_28_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_3_data_19 <= io_in_c_bypass_28_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_3_is_stationary_19 <= io_in_c_bypass_28_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_0_data_19 <= io_in_c_bypass_29_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_0_is_stationary_19 <= io_in_c_bypass_29_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_1_data_19 <= io_in_c_bypass_29_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_1_is_stationary_19 <= io_in_c_bypass_29_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_2_data_19 <= io_in_c_bypass_29_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_2_is_stationary_19 <= io_in_c_bypass_29_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_3_data_19 <= io_in_c_bypass_29_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_3_is_stationary_19 <= io_in_c_bypass_29_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_0_data_19 <= io_in_c_bypass_30_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_0_is_stationary_19 <= io_in_c_bypass_30_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_1_data_19 <= io_in_c_bypass_30_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_1_is_stationary_19 <= io_in_c_bypass_30_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_2_data_19 <= io_in_c_bypass_30_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_2_is_stationary_19 <= io_in_c_bypass_30_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_3_data_19 <= io_in_c_bypass_30_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_3_is_stationary_19 <= io_in_c_bypass_30_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_0_data_19 <= io_in_c_bypass_31_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_0_is_stationary_19 <= io_in_c_bypass_31_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_1_data_19 <= io_in_c_bypass_31_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_1_is_stationary_19 <= io_in_c_bypass_31_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_2_data_19 <= io_in_c_bypass_31_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_2_is_stationary_19 <= io_in_c_bypass_31_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_3_data_19 <= io_in_c_bypass_31_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_3_is_stationary_19 <= io_in_c_bypass_31_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_0_data_20 <= io_in_c_bypass_0_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_0_is_stationary_20 <= io_in_c_bypass_0_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_1_data_20 <= io_in_c_bypass_0_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_1_is_stationary_20 <= io_in_c_bypass_0_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_2_data_20 <= io_in_c_bypass_0_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_2_is_stationary_20 <= io_in_c_bypass_0_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_3_data_20 <= io_in_c_bypass_0_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_3_is_stationary_20 <= io_in_c_bypass_0_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_0_data_20 <= io_in_c_bypass_1_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_0_is_stationary_20 <= io_in_c_bypass_1_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_1_data_20 <= io_in_c_bypass_1_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_1_is_stationary_20 <= io_in_c_bypass_1_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_2_data_20 <= io_in_c_bypass_1_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_2_is_stationary_20 <= io_in_c_bypass_1_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_3_data_20 <= io_in_c_bypass_1_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_3_is_stationary_20 <= io_in_c_bypass_1_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_0_data_20 <= io_in_c_bypass_2_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_0_is_stationary_20 <= io_in_c_bypass_2_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_1_data_20 <= io_in_c_bypass_2_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_1_is_stationary_20 <= io_in_c_bypass_2_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_2_data_20 <= io_in_c_bypass_2_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_2_is_stationary_20 <= io_in_c_bypass_2_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_3_data_20 <= io_in_c_bypass_2_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_3_is_stationary_20 <= io_in_c_bypass_2_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_0_data_20 <= io_in_c_bypass_3_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_0_is_stationary_20 <= io_in_c_bypass_3_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_1_data_20 <= io_in_c_bypass_3_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_1_is_stationary_20 <= io_in_c_bypass_3_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_2_data_20 <= io_in_c_bypass_3_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_2_is_stationary_20 <= io_in_c_bypass_3_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_3_data_20 <= io_in_c_bypass_3_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_3_is_stationary_20 <= io_in_c_bypass_3_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_0_data_20 <= io_in_c_bypass_4_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_0_is_stationary_20 <= io_in_c_bypass_4_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_1_data_20 <= io_in_c_bypass_4_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_1_is_stationary_20 <= io_in_c_bypass_4_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_2_data_20 <= io_in_c_bypass_4_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_2_is_stationary_20 <= io_in_c_bypass_4_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_3_data_20 <= io_in_c_bypass_4_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_3_is_stationary_20 <= io_in_c_bypass_4_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_0_data_20 <= io_in_c_bypass_5_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_0_is_stationary_20 <= io_in_c_bypass_5_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_1_data_20 <= io_in_c_bypass_5_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_1_is_stationary_20 <= io_in_c_bypass_5_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_2_data_20 <= io_in_c_bypass_5_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_2_is_stationary_20 <= io_in_c_bypass_5_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_3_data_20 <= io_in_c_bypass_5_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_3_is_stationary_20 <= io_in_c_bypass_5_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_0_data_20 <= io_in_c_bypass_6_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_0_is_stationary_20 <= io_in_c_bypass_6_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_1_data_20 <= io_in_c_bypass_6_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_1_is_stationary_20 <= io_in_c_bypass_6_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_2_data_20 <= io_in_c_bypass_6_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_2_is_stationary_20 <= io_in_c_bypass_6_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_3_data_20 <= io_in_c_bypass_6_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_3_is_stationary_20 <= io_in_c_bypass_6_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_0_data_20 <= io_in_c_bypass_7_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_0_is_stationary_20 <= io_in_c_bypass_7_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_1_data_20 <= io_in_c_bypass_7_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_1_is_stationary_20 <= io_in_c_bypass_7_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_2_data_20 <= io_in_c_bypass_7_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_2_is_stationary_20 <= io_in_c_bypass_7_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_3_data_20 <= io_in_c_bypass_7_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_3_is_stationary_20 <= io_in_c_bypass_7_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_0_data_20 <= io_in_c_bypass_8_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_0_is_stationary_20 <= io_in_c_bypass_8_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_1_data_20 <= io_in_c_bypass_8_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_1_is_stationary_20 <= io_in_c_bypass_8_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_2_data_20 <= io_in_c_bypass_8_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_2_is_stationary_20 <= io_in_c_bypass_8_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_3_data_20 <= io_in_c_bypass_8_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_3_is_stationary_20 <= io_in_c_bypass_8_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_0_data_20 <= io_in_c_bypass_9_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_0_is_stationary_20 <= io_in_c_bypass_9_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_1_data_20 <= io_in_c_bypass_9_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_1_is_stationary_20 <= io_in_c_bypass_9_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_2_data_20 <= io_in_c_bypass_9_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_2_is_stationary_20 <= io_in_c_bypass_9_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_3_data_20 <= io_in_c_bypass_9_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_3_is_stationary_20 <= io_in_c_bypass_9_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_0_data_20 <= io_in_c_bypass_10_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_0_is_stationary_20 <= io_in_c_bypass_10_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_1_data_20 <= io_in_c_bypass_10_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_1_is_stationary_20 <= io_in_c_bypass_10_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_2_data_20 <= io_in_c_bypass_10_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_2_is_stationary_20 <= io_in_c_bypass_10_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_3_data_20 <= io_in_c_bypass_10_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_3_is_stationary_20 <= io_in_c_bypass_10_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_0_data_20 <= io_in_c_bypass_11_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_0_is_stationary_20 <= io_in_c_bypass_11_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_1_data_20 <= io_in_c_bypass_11_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_1_is_stationary_20 <= io_in_c_bypass_11_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_2_data_20 <= io_in_c_bypass_11_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_2_is_stationary_20 <= io_in_c_bypass_11_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_3_data_20 <= io_in_c_bypass_11_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_3_is_stationary_20 <= io_in_c_bypass_11_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_0_data_20 <= io_in_c_bypass_12_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_0_is_stationary_20 <= io_in_c_bypass_12_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_1_data_20 <= io_in_c_bypass_12_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_1_is_stationary_20 <= io_in_c_bypass_12_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_2_data_20 <= io_in_c_bypass_12_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_2_is_stationary_20 <= io_in_c_bypass_12_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_3_data_20 <= io_in_c_bypass_12_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_3_is_stationary_20 <= io_in_c_bypass_12_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_0_data_20 <= io_in_c_bypass_13_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_0_is_stationary_20 <= io_in_c_bypass_13_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_1_data_20 <= io_in_c_bypass_13_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_1_is_stationary_20 <= io_in_c_bypass_13_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_2_data_20 <= io_in_c_bypass_13_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_2_is_stationary_20 <= io_in_c_bypass_13_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_3_data_20 <= io_in_c_bypass_13_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_3_is_stationary_20 <= io_in_c_bypass_13_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_0_data_20 <= io_in_c_bypass_14_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_0_is_stationary_20 <= io_in_c_bypass_14_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_1_data_20 <= io_in_c_bypass_14_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_1_is_stationary_20 <= io_in_c_bypass_14_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_2_data_20 <= io_in_c_bypass_14_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_2_is_stationary_20 <= io_in_c_bypass_14_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_3_data_20 <= io_in_c_bypass_14_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_3_is_stationary_20 <= io_in_c_bypass_14_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_0_data_20 <= io_in_c_bypass_15_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_0_is_stationary_20 <= io_in_c_bypass_15_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_1_data_20 <= io_in_c_bypass_15_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_1_is_stationary_20 <= io_in_c_bypass_15_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_2_data_20 <= io_in_c_bypass_15_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_2_is_stationary_20 <= io_in_c_bypass_15_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_3_data_20 <= io_in_c_bypass_15_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_3_is_stationary_20 <= io_in_c_bypass_15_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_0_data_20 <= io_in_c_bypass_16_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_0_is_stationary_20 <= io_in_c_bypass_16_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_1_data_20 <= io_in_c_bypass_16_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_1_is_stationary_20 <= io_in_c_bypass_16_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_2_data_20 <= io_in_c_bypass_16_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_2_is_stationary_20 <= io_in_c_bypass_16_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_3_data_20 <= io_in_c_bypass_16_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_3_is_stationary_20 <= io_in_c_bypass_16_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_0_data_20 <= io_in_c_bypass_17_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_0_is_stationary_20 <= io_in_c_bypass_17_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_1_data_20 <= io_in_c_bypass_17_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_1_is_stationary_20 <= io_in_c_bypass_17_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_2_data_20 <= io_in_c_bypass_17_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_2_is_stationary_20 <= io_in_c_bypass_17_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_3_data_20 <= io_in_c_bypass_17_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_3_is_stationary_20 <= io_in_c_bypass_17_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_0_data_20 <= io_in_c_bypass_18_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_0_is_stationary_20 <= io_in_c_bypass_18_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_1_data_20 <= io_in_c_bypass_18_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_1_is_stationary_20 <= io_in_c_bypass_18_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_2_data_20 <= io_in_c_bypass_18_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_2_is_stationary_20 <= io_in_c_bypass_18_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_3_data_20 <= io_in_c_bypass_18_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_3_is_stationary_20 <= io_in_c_bypass_18_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_0_data_20 <= io_in_c_bypass_19_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_0_is_stationary_20 <= io_in_c_bypass_19_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_1_data_20 <= io_in_c_bypass_19_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_1_is_stationary_20 <= io_in_c_bypass_19_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_2_data_20 <= io_in_c_bypass_19_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_2_is_stationary_20 <= io_in_c_bypass_19_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_3_data_20 <= io_in_c_bypass_19_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_3_is_stationary_20 <= io_in_c_bypass_19_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_0_data_20 <= io_in_c_bypass_20_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_0_is_stationary_20 <= io_in_c_bypass_20_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_1_data_20 <= io_in_c_bypass_20_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_1_is_stationary_20 <= io_in_c_bypass_20_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_2_data_20 <= io_in_c_bypass_20_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_2_is_stationary_20 <= io_in_c_bypass_20_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_3_data_20 <= io_in_c_bypass_20_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_3_is_stationary_20 <= io_in_c_bypass_20_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_0_data_20 <= io_in_c_bypass_21_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_0_is_stationary_20 <= io_in_c_bypass_21_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_1_data_20 <= io_in_c_bypass_21_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_1_is_stationary_20 <= io_in_c_bypass_21_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_2_data_20 <= io_in_c_bypass_21_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_2_is_stationary_20 <= io_in_c_bypass_21_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_3_data_20 <= io_in_c_bypass_21_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_3_is_stationary_20 <= io_in_c_bypass_21_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_0_data_20 <= io_in_c_bypass_22_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_0_is_stationary_20 <= io_in_c_bypass_22_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_1_data_20 <= io_in_c_bypass_22_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_1_is_stationary_20 <= io_in_c_bypass_22_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_2_data_20 <= io_in_c_bypass_22_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_2_is_stationary_20 <= io_in_c_bypass_22_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_3_data_20 <= io_in_c_bypass_22_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_3_is_stationary_20 <= io_in_c_bypass_22_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_0_data_20 <= io_in_c_bypass_23_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_0_is_stationary_20 <= io_in_c_bypass_23_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_1_data_20 <= io_in_c_bypass_23_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_1_is_stationary_20 <= io_in_c_bypass_23_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_2_data_20 <= io_in_c_bypass_23_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_2_is_stationary_20 <= io_in_c_bypass_23_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_3_data_20 <= io_in_c_bypass_23_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_3_is_stationary_20 <= io_in_c_bypass_23_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_0_data_20 <= io_in_c_bypass_24_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_0_is_stationary_20 <= io_in_c_bypass_24_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_1_data_20 <= io_in_c_bypass_24_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_1_is_stationary_20 <= io_in_c_bypass_24_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_2_data_20 <= io_in_c_bypass_24_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_2_is_stationary_20 <= io_in_c_bypass_24_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_3_data_20 <= io_in_c_bypass_24_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_3_is_stationary_20 <= io_in_c_bypass_24_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_0_data_20 <= io_in_c_bypass_25_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_0_is_stationary_20 <= io_in_c_bypass_25_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_1_data_20 <= io_in_c_bypass_25_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_1_is_stationary_20 <= io_in_c_bypass_25_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_2_data_20 <= io_in_c_bypass_25_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_2_is_stationary_20 <= io_in_c_bypass_25_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_3_data_20 <= io_in_c_bypass_25_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_3_is_stationary_20 <= io_in_c_bypass_25_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_0_data_20 <= io_in_c_bypass_26_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_0_is_stationary_20 <= io_in_c_bypass_26_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_1_data_20 <= io_in_c_bypass_26_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_1_is_stationary_20 <= io_in_c_bypass_26_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_2_data_20 <= io_in_c_bypass_26_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_2_is_stationary_20 <= io_in_c_bypass_26_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_3_data_20 <= io_in_c_bypass_26_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_3_is_stationary_20 <= io_in_c_bypass_26_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_0_data_20 <= io_in_c_bypass_27_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_0_is_stationary_20 <= io_in_c_bypass_27_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_1_data_20 <= io_in_c_bypass_27_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_1_is_stationary_20 <= io_in_c_bypass_27_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_2_data_20 <= io_in_c_bypass_27_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_2_is_stationary_20 <= io_in_c_bypass_27_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_3_data_20 <= io_in_c_bypass_27_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_3_is_stationary_20 <= io_in_c_bypass_27_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_0_data_20 <= io_in_c_bypass_28_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_0_is_stationary_20 <= io_in_c_bypass_28_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_1_data_20 <= io_in_c_bypass_28_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_1_is_stationary_20 <= io_in_c_bypass_28_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_2_data_20 <= io_in_c_bypass_28_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_2_is_stationary_20 <= io_in_c_bypass_28_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_3_data_20 <= io_in_c_bypass_28_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_3_is_stationary_20 <= io_in_c_bypass_28_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_0_data_20 <= io_in_c_bypass_29_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_0_is_stationary_20 <= io_in_c_bypass_29_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_1_data_20 <= io_in_c_bypass_29_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_1_is_stationary_20 <= io_in_c_bypass_29_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_2_data_20 <= io_in_c_bypass_29_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_2_is_stationary_20 <= io_in_c_bypass_29_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_3_data_20 <= io_in_c_bypass_29_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_3_is_stationary_20 <= io_in_c_bypass_29_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_0_data_20 <= io_in_c_bypass_30_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_0_is_stationary_20 <= io_in_c_bypass_30_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_1_data_20 <= io_in_c_bypass_30_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_1_is_stationary_20 <= io_in_c_bypass_30_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_2_data_20 <= io_in_c_bypass_30_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_2_is_stationary_20 <= io_in_c_bypass_30_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_3_data_20 <= io_in_c_bypass_30_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_3_is_stationary_20 <= io_in_c_bypass_30_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_0_data_20 <= io_in_c_bypass_31_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_0_is_stationary_20 <= io_in_c_bypass_31_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_1_data_20 <= io_in_c_bypass_31_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_1_is_stationary_20 <= io_in_c_bypass_31_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_2_data_20 <= io_in_c_bypass_31_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_2_is_stationary_20 <= io_in_c_bypass_31_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_3_data_20 <= io_in_c_bypass_31_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_3_is_stationary_20 <= io_in_c_bypass_31_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_0_data_21 <= io_in_c_bypass_0_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_0_is_stationary_21 <= io_in_c_bypass_0_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_1_data_21 <= io_in_c_bypass_0_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_1_is_stationary_21 <= io_in_c_bypass_0_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_2_data_21 <= io_in_c_bypass_0_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_2_is_stationary_21 <= io_in_c_bypass_0_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_3_data_21 <= io_in_c_bypass_0_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_3_is_stationary_21 <= io_in_c_bypass_0_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_0_data_21 <= io_in_c_bypass_1_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_0_is_stationary_21 <= io_in_c_bypass_1_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_1_data_21 <= io_in_c_bypass_1_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_1_is_stationary_21 <= io_in_c_bypass_1_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_2_data_21 <= io_in_c_bypass_1_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_2_is_stationary_21 <= io_in_c_bypass_1_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_3_data_21 <= io_in_c_bypass_1_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_3_is_stationary_21 <= io_in_c_bypass_1_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_0_data_21 <= io_in_c_bypass_2_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_0_is_stationary_21 <= io_in_c_bypass_2_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_1_data_21 <= io_in_c_bypass_2_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_1_is_stationary_21 <= io_in_c_bypass_2_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_2_data_21 <= io_in_c_bypass_2_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_2_is_stationary_21 <= io_in_c_bypass_2_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_3_data_21 <= io_in_c_bypass_2_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_3_is_stationary_21 <= io_in_c_bypass_2_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_0_data_21 <= io_in_c_bypass_3_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_0_is_stationary_21 <= io_in_c_bypass_3_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_1_data_21 <= io_in_c_bypass_3_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_1_is_stationary_21 <= io_in_c_bypass_3_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_2_data_21 <= io_in_c_bypass_3_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_2_is_stationary_21 <= io_in_c_bypass_3_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_3_data_21 <= io_in_c_bypass_3_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_3_is_stationary_21 <= io_in_c_bypass_3_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_0_data_21 <= io_in_c_bypass_4_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_0_is_stationary_21 <= io_in_c_bypass_4_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_1_data_21 <= io_in_c_bypass_4_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_1_is_stationary_21 <= io_in_c_bypass_4_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_2_data_21 <= io_in_c_bypass_4_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_2_is_stationary_21 <= io_in_c_bypass_4_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_3_data_21 <= io_in_c_bypass_4_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_3_is_stationary_21 <= io_in_c_bypass_4_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_0_data_21 <= io_in_c_bypass_5_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_0_is_stationary_21 <= io_in_c_bypass_5_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_1_data_21 <= io_in_c_bypass_5_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_1_is_stationary_21 <= io_in_c_bypass_5_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_2_data_21 <= io_in_c_bypass_5_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_2_is_stationary_21 <= io_in_c_bypass_5_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_3_data_21 <= io_in_c_bypass_5_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_3_is_stationary_21 <= io_in_c_bypass_5_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_0_data_21 <= io_in_c_bypass_6_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_0_is_stationary_21 <= io_in_c_bypass_6_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_1_data_21 <= io_in_c_bypass_6_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_1_is_stationary_21 <= io_in_c_bypass_6_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_2_data_21 <= io_in_c_bypass_6_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_2_is_stationary_21 <= io_in_c_bypass_6_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_3_data_21 <= io_in_c_bypass_6_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_3_is_stationary_21 <= io_in_c_bypass_6_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_0_data_21 <= io_in_c_bypass_7_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_0_is_stationary_21 <= io_in_c_bypass_7_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_1_data_21 <= io_in_c_bypass_7_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_1_is_stationary_21 <= io_in_c_bypass_7_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_2_data_21 <= io_in_c_bypass_7_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_2_is_stationary_21 <= io_in_c_bypass_7_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_3_data_21 <= io_in_c_bypass_7_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_3_is_stationary_21 <= io_in_c_bypass_7_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_0_data_21 <= io_in_c_bypass_8_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_0_is_stationary_21 <= io_in_c_bypass_8_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_1_data_21 <= io_in_c_bypass_8_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_1_is_stationary_21 <= io_in_c_bypass_8_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_2_data_21 <= io_in_c_bypass_8_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_2_is_stationary_21 <= io_in_c_bypass_8_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_3_data_21 <= io_in_c_bypass_8_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_3_is_stationary_21 <= io_in_c_bypass_8_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_0_data_21 <= io_in_c_bypass_9_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_0_is_stationary_21 <= io_in_c_bypass_9_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_1_data_21 <= io_in_c_bypass_9_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_1_is_stationary_21 <= io_in_c_bypass_9_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_2_data_21 <= io_in_c_bypass_9_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_2_is_stationary_21 <= io_in_c_bypass_9_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_3_data_21 <= io_in_c_bypass_9_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_3_is_stationary_21 <= io_in_c_bypass_9_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_0_data_21 <= io_in_c_bypass_10_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_0_is_stationary_21 <= io_in_c_bypass_10_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_1_data_21 <= io_in_c_bypass_10_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_1_is_stationary_21 <= io_in_c_bypass_10_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_2_data_21 <= io_in_c_bypass_10_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_2_is_stationary_21 <= io_in_c_bypass_10_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_3_data_21 <= io_in_c_bypass_10_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_3_is_stationary_21 <= io_in_c_bypass_10_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_0_data_21 <= io_in_c_bypass_11_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_0_is_stationary_21 <= io_in_c_bypass_11_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_1_data_21 <= io_in_c_bypass_11_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_1_is_stationary_21 <= io_in_c_bypass_11_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_2_data_21 <= io_in_c_bypass_11_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_2_is_stationary_21 <= io_in_c_bypass_11_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_3_data_21 <= io_in_c_bypass_11_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_3_is_stationary_21 <= io_in_c_bypass_11_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_0_data_21 <= io_in_c_bypass_12_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_0_is_stationary_21 <= io_in_c_bypass_12_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_1_data_21 <= io_in_c_bypass_12_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_1_is_stationary_21 <= io_in_c_bypass_12_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_2_data_21 <= io_in_c_bypass_12_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_2_is_stationary_21 <= io_in_c_bypass_12_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_3_data_21 <= io_in_c_bypass_12_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_3_is_stationary_21 <= io_in_c_bypass_12_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_0_data_21 <= io_in_c_bypass_13_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_0_is_stationary_21 <= io_in_c_bypass_13_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_1_data_21 <= io_in_c_bypass_13_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_1_is_stationary_21 <= io_in_c_bypass_13_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_2_data_21 <= io_in_c_bypass_13_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_2_is_stationary_21 <= io_in_c_bypass_13_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_3_data_21 <= io_in_c_bypass_13_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_3_is_stationary_21 <= io_in_c_bypass_13_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_0_data_21 <= io_in_c_bypass_14_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_0_is_stationary_21 <= io_in_c_bypass_14_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_1_data_21 <= io_in_c_bypass_14_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_1_is_stationary_21 <= io_in_c_bypass_14_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_2_data_21 <= io_in_c_bypass_14_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_2_is_stationary_21 <= io_in_c_bypass_14_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_3_data_21 <= io_in_c_bypass_14_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_3_is_stationary_21 <= io_in_c_bypass_14_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_0_data_21 <= io_in_c_bypass_15_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_0_is_stationary_21 <= io_in_c_bypass_15_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_1_data_21 <= io_in_c_bypass_15_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_1_is_stationary_21 <= io_in_c_bypass_15_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_2_data_21 <= io_in_c_bypass_15_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_2_is_stationary_21 <= io_in_c_bypass_15_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_3_data_21 <= io_in_c_bypass_15_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_3_is_stationary_21 <= io_in_c_bypass_15_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_0_data_21 <= io_in_c_bypass_16_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_0_is_stationary_21 <= io_in_c_bypass_16_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_1_data_21 <= io_in_c_bypass_16_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_1_is_stationary_21 <= io_in_c_bypass_16_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_2_data_21 <= io_in_c_bypass_16_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_2_is_stationary_21 <= io_in_c_bypass_16_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_3_data_21 <= io_in_c_bypass_16_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_3_is_stationary_21 <= io_in_c_bypass_16_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_0_data_21 <= io_in_c_bypass_17_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_0_is_stationary_21 <= io_in_c_bypass_17_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_1_data_21 <= io_in_c_bypass_17_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_1_is_stationary_21 <= io_in_c_bypass_17_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_2_data_21 <= io_in_c_bypass_17_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_2_is_stationary_21 <= io_in_c_bypass_17_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_3_data_21 <= io_in_c_bypass_17_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_3_is_stationary_21 <= io_in_c_bypass_17_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_0_data_21 <= io_in_c_bypass_18_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_0_is_stationary_21 <= io_in_c_bypass_18_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_1_data_21 <= io_in_c_bypass_18_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_1_is_stationary_21 <= io_in_c_bypass_18_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_2_data_21 <= io_in_c_bypass_18_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_2_is_stationary_21 <= io_in_c_bypass_18_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_3_data_21 <= io_in_c_bypass_18_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_3_is_stationary_21 <= io_in_c_bypass_18_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_0_data_21 <= io_in_c_bypass_19_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_0_is_stationary_21 <= io_in_c_bypass_19_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_1_data_21 <= io_in_c_bypass_19_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_1_is_stationary_21 <= io_in_c_bypass_19_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_2_data_21 <= io_in_c_bypass_19_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_2_is_stationary_21 <= io_in_c_bypass_19_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_3_data_21 <= io_in_c_bypass_19_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_3_is_stationary_21 <= io_in_c_bypass_19_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_0_data_21 <= io_in_c_bypass_20_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_0_is_stationary_21 <= io_in_c_bypass_20_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_1_data_21 <= io_in_c_bypass_20_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_1_is_stationary_21 <= io_in_c_bypass_20_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_2_data_21 <= io_in_c_bypass_20_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_2_is_stationary_21 <= io_in_c_bypass_20_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_3_data_21 <= io_in_c_bypass_20_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_3_is_stationary_21 <= io_in_c_bypass_20_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_0_data_21 <= io_in_c_bypass_21_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_0_is_stationary_21 <= io_in_c_bypass_21_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_1_data_21 <= io_in_c_bypass_21_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_1_is_stationary_21 <= io_in_c_bypass_21_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_2_data_21 <= io_in_c_bypass_21_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_2_is_stationary_21 <= io_in_c_bypass_21_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_3_data_21 <= io_in_c_bypass_21_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_3_is_stationary_21 <= io_in_c_bypass_21_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_0_data_21 <= io_in_c_bypass_22_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_0_is_stationary_21 <= io_in_c_bypass_22_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_1_data_21 <= io_in_c_bypass_22_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_1_is_stationary_21 <= io_in_c_bypass_22_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_2_data_21 <= io_in_c_bypass_22_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_2_is_stationary_21 <= io_in_c_bypass_22_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_3_data_21 <= io_in_c_bypass_22_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_3_is_stationary_21 <= io_in_c_bypass_22_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_0_data_21 <= io_in_c_bypass_23_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_0_is_stationary_21 <= io_in_c_bypass_23_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_1_data_21 <= io_in_c_bypass_23_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_1_is_stationary_21 <= io_in_c_bypass_23_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_2_data_21 <= io_in_c_bypass_23_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_2_is_stationary_21 <= io_in_c_bypass_23_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_3_data_21 <= io_in_c_bypass_23_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_3_is_stationary_21 <= io_in_c_bypass_23_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_0_data_21 <= io_in_c_bypass_24_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_0_is_stationary_21 <= io_in_c_bypass_24_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_1_data_21 <= io_in_c_bypass_24_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_1_is_stationary_21 <= io_in_c_bypass_24_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_2_data_21 <= io_in_c_bypass_24_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_2_is_stationary_21 <= io_in_c_bypass_24_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_3_data_21 <= io_in_c_bypass_24_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_3_is_stationary_21 <= io_in_c_bypass_24_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_0_data_21 <= io_in_c_bypass_25_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_0_is_stationary_21 <= io_in_c_bypass_25_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_1_data_21 <= io_in_c_bypass_25_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_1_is_stationary_21 <= io_in_c_bypass_25_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_2_data_21 <= io_in_c_bypass_25_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_2_is_stationary_21 <= io_in_c_bypass_25_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_3_data_21 <= io_in_c_bypass_25_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_3_is_stationary_21 <= io_in_c_bypass_25_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_0_data_21 <= io_in_c_bypass_26_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_0_is_stationary_21 <= io_in_c_bypass_26_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_1_data_21 <= io_in_c_bypass_26_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_1_is_stationary_21 <= io_in_c_bypass_26_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_2_data_21 <= io_in_c_bypass_26_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_2_is_stationary_21 <= io_in_c_bypass_26_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_3_data_21 <= io_in_c_bypass_26_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_3_is_stationary_21 <= io_in_c_bypass_26_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_0_data_21 <= io_in_c_bypass_27_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_0_is_stationary_21 <= io_in_c_bypass_27_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_1_data_21 <= io_in_c_bypass_27_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_1_is_stationary_21 <= io_in_c_bypass_27_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_2_data_21 <= io_in_c_bypass_27_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_2_is_stationary_21 <= io_in_c_bypass_27_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_3_data_21 <= io_in_c_bypass_27_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_3_is_stationary_21 <= io_in_c_bypass_27_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_0_data_21 <= io_in_c_bypass_28_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_0_is_stationary_21 <= io_in_c_bypass_28_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_1_data_21 <= io_in_c_bypass_28_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_1_is_stationary_21 <= io_in_c_bypass_28_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_2_data_21 <= io_in_c_bypass_28_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_2_is_stationary_21 <= io_in_c_bypass_28_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_3_data_21 <= io_in_c_bypass_28_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_3_is_stationary_21 <= io_in_c_bypass_28_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_0_data_21 <= io_in_c_bypass_29_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_0_is_stationary_21 <= io_in_c_bypass_29_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_1_data_21 <= io_in_c_bypass_29_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_1_is_stationary_21 <= io_in_c_bypass_29_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_2_data_21 <= io_in_c_bypass_29_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_2_is_stationary_21 <= io_in_c_bypass_29_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_3_data_21 <= io_in_c_bypass_29_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_3_is_stationary_21 <= io_in_c_bypass_29_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_0_data_21 <= io_in_c_bypass_30_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_0_is_stationary_21 <= io_in_c_bypass_30_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_1_data_21 <= io_in_c_bypass_30_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_1_is_stationary_21 <= io_in_c_bypass_30_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_2_data_21 <= io_in_c_bypass_30_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_2_is_stationary_21 <= io_in_c_bypass_30_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_3_data_21 <= io_in_c_bypass_30_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_3_is_stationary_21 <= io_in_c_bypass_30_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_0_data_21 <= io_in_c_bypass_31_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_0_is_stationary_21 <= io_in_c_bypass_31_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_1_data_21 <= io_in_c_bypass_31_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_1_is_stationary_21 <= io_in_c_bypass_31_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_2_data_21 <= io_in_c_bypass_31_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_2_is_stationary_21 <= io_in_c_bypass_31_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_3_data_21 <= io_in_c_bypass_31_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_3_is_stationary_21 <= io_in_c_bypass_31_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_0_data_22 <= io_in_c_bypass_0_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_0_is_stationary_22 <= io_in_c_bypass_0_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_1_data_22 <= io_in_c_bypass_0_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_1_is_stationary_22 <= io_in_c_bypass_0_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_2_data_22 <= io_in_c_bypass_0_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_2_is_stationary_22 <= io_in_c_bypass_0_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_3_data_22 <= io_in_c_bypass_0_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_3_is_stationary_22 <= io_in_c_bypass_0_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_0_data_22 <= io_in_c_bypass_1_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_0_is_stationary_22 <= io_in_c_bypass_1_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_1_data_22 <= io_in_c_bypass_1_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_1_is_stationary_22 <= io_in_c_bypass_1_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_2_data_22 <= io_in_c_bypass_1_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_2_is_stationary_22 <= io_in_c_bypass_1_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_3_data_22 <= io_in_c_bypass_1_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_3_is_stationary_22 <= io_in_c_bypass_1_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_0_data_22 <= io_in_c_bypass_2_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_0_is_stationary_22 <= io_in_c_bypass_2_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_1_data_22 <= io_in_c_bypass_2_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_1_is_stationary_22 <= io_in_c_bypass_2_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_2_data_22 <= io_in_c_bypass_2_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_2_is_stationary_22 <= io_in_c_bypass_2_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_3_data_22 <= io_in_c_bypass_2_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_3_is_stationary_22 <= io_in_c_bypass_2_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_0_data_22 <= io_in_c_bypass_3_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_0_is_stationary_22 <= io_in_c_bypass_3_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_1_data_22 <= io_in_c_bypass_3_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_1_is_stationary_22 <= io_in_c_bypass_3_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_2_data_22 <= io_in_c_bypass_3_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_2_is_stationary_22 <= io_in_c_bypass_3_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_3_data_22 <= io_in_c_bypass_3_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_3_is_stationary_22 <= io_in_c_bypass_3_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_0_data_22 <= io_in_c_bypass_4_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_0_is_stationary_22 <= io_in_c_bypass_4_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_1_data_22 <= io_in_c_bypass_4_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_1_is_stationary_22 <= io_in_c_bypass_4_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_2_data_22 <= io_in_c_bypass_4_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_2_is_stationary_22 <= io_in_c_bypass_4_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_3_data_22 <= io_in_c_bypass_4_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_3_is_stationary_22 <= io_in_c_bypass_4_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_0_data_22 <= io_in_c_bypass_5_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_0_is_stationary_22 <= io_in_c_bypass_5_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_1_data_22 <= io_in_c_bypass_5_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_1_is_stationary_22 <= io_in_c_bypass_5_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_2_data_22 <= io_in_c_bypass_5_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_2_is_stationary_22 <= io_in_c_bypass_5_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_3_data_22 <= io_in_c_bypass_5_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_3_is_stationary_22 <= io_in_c_bypass_5_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_0_data_22 <= io_in_c_bypass_6_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_0_is_stationary_22 <= io_in_c_bypass_6_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_1_data_22 <= io_in_c_bypass_6_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_1_is_stationary_22 <= io_in_c_bypass_6_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_2_data_22 <= io_in_c_bypass_6_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_2_is_stationary_22 <= io_in_c_bypass_6_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_3_data_22 <= io_in_c_bypass_6_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_3_is_stationary_22 <= io_in_c_bypass_6_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_0_data_22 <= io_in_c_bypass_7_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_0_is_stationary_22 <= io_in_c_bypass_7_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_1_data_22 <= io_in_c_bypass_7_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_1_is_stationary_22 <= io_in_c_bypass_7_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_2_data_22 <= io_in_c_bypass_7_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_2_is_stationary_22 <= io_in_c_bypass_7_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_3_data_22 <= io_in_c_bypass_7_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_3_is_stationary_22 <= io_in_c_bypass_7_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_0_data_22 <= io_in_c_bypass_8_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_0_is_stationary_22 <= io_in_c_bypass_8_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_1_data_22 <= io_in_c_bypass_8_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_1_is_stationary_22 <= io_in_c_bypass_8_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_2_data_22 <= io_in_c_bypass_8_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_2_is_stationary_22 <= io_in_c_bypass_8_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_3_data_22 <= io_in_c_bypass_8_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_3_is_stationary_22 <= io_in_c_bypass_8_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_0_data_22 <= io_in_c_bypass_9_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_0_is_stationary_22 <= io_in_c_bypass_9_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_1_data_22 <= io_in_c_bypass_9_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_1_is_stationary_22 <= io_in_c_bypass_9_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_2_data_22 <= io_in_c_bypass_9_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_2_is_stationary_22 <= io_in_c_bypass_9_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_3_data_22 <= io_in_c_bypass_9_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_3_is_stationary_22 <= io_in_c_bypass_9_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_0_data_22 <= io_in_c_bypass_10_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_0_is_stationary_22 <= io_in_c_bypass_10_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_1_data_22 <= io_in_c_bypass_10_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_1_is_stationary_22 <= io_in_c_bypass_10_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_2_data_22 <= io_in_c_bypass_10_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_2_is_stationary_22 <= io_in_c_bypass_10_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_3_data_22 <= io_in_c_bypass_10_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_3_is_stationary_22 <= io_in_c_bypass_10_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_0_data_22 <= io_in_c_bypass_11_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_0_is_stationary_22 <= io_in_c_bypass_11_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_1_data_22 <= io_in_c_bypass_11_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_1_is_stationary_22 <= io_in_c_bypass_11_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_2_data_22 <= io_in_c_bypass_11_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_2_is_stationary_22 <= io_in_c_bypass_11_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_3_data_22 <= io_in_c_bypass_11_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_3_is_stationary_22 <= io_in_c_bypass_11_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_0_data_22 <= io_in_c_bypass_12_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_0_is_stationary_22 <= io_in_c_bypass_12_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_1_data_22 <= io_in_c_bypass_12_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_1_is_stationary_22 <= io_in_c_bypass_12_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_2_data_22 <= io_in_c_bypass_12_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_2_is_stationary_22 <= io_in_c_bypass_12_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_3_data_22 <= io_in_c_bypass_12_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_3_is_stationary_22 <= io_in_c_bypass_12_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_0_data_22 <= io_in_c_bypass_13_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_0_is_stationary_22 <= io_in_c_bypass_13_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_1_data_22 <= io_in_c_bypass_13_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_1_is_stationary_22 <= io_in_c_bypass_13_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_2_data_22 <= io_in_c_bypass_13_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_2_is_stationary_22 <= io_in_c_bypass_13_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_3_data_22 <= io_in_c_bypass_13_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_3_is_stationary_22 <= io_in_c_bypass_13_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_0_data_22 <= io_in_c_bypass_14_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_0_is_stationary_22 <= io_in_c_bypass_14_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_1_data_22 <= io_in_c_bypass_14_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_1_is_stationary_22 <= io_in_c_bypass_14_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_2_data_22 <= io_in_c_bypass_14_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_2_is_stationary_22 <= io_in_c_bypass_14_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_3_data_22 <= io_in_c_bypass_14_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_3_is_stationary_22 <= io_in_c_bypass_14_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_0_data_22 <= io_in_c_bypass_15_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_0_is_stationary_22 <= io_in_c_bypass_15_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_1_data_22 <= io_in_c_bypass_15_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_1_is_stationary_22 <= io_in_c_bypass_15_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_2_data_22 <= io_in_c_bypass_15_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_2_is_stationary_22 <= io_in_c_bypass_15_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_3_data_22 <= io_in_c_bypass_15_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_3_is_stationary_22 <= io_in_c_bypass_15_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_0_data_22 <= io_in_c_bypass_16_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_0_is_stationary_22 <= io_in_c_bypass_16_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_1_data_22 <= io_in_c_bypass_16_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_1_is_stationary_22 <= io_in_c_bypass_16_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_2_data_22 <= io_in_c_bypass_16_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_2_is_stationary_22 <= io_in_c_bypass_16_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_3_data_22 <= io_in_c_bypass_16_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_3_is_stationary_22 <= io_in_c_bypass_16_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_0_data_22 <= io_in_c_bypass_17_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_0_is_stationary_22 <= io_in_c_bypass_17_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_1_data_22 <= io_in_c_bypass_17_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_1_is_stationary_22 <= io_in_c_bypass_17_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_2_data_22 <= io_in_c_bypass_17_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_2_is_stationary_22 <= io_in_c_bypass_17_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_3_data_22 <= io_in_c_bypass_17_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_3_is_stationary_22 <= io_in_c_bypass_17_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_0_data_22 <= io_in_c_bypass_18_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_0_is_stationary_22 <= io_in_c_bypass_18_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_1_data_22 <= io_in_c_bypass_18_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_1_is_stationary_22 <= io_in_c_bypass_18_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_2_data_22 <= io_in_c_bypass_18_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_2_is_stationary_22 <= io_in_c_bypass_18_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_3_data_22 <= io_in_c_bypass_18_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_3_is_stationary_22 <= io_in_c_bypass_18_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_0_data_22 <= io_in_c_bypass_19_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_0_is_stationary_22 <= io_in_c_bypass_19_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_1_data_22 <= io_in_c_bypass_19_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_1_is_stationary_22 <= io_in_c_bypass_19_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_2_data_22 <= io_in_c_bypass_19_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_2_is_stationary_22 <= io_in_c_bypass_19_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_3_data_22 <= io_in_c_bypass_19_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_3_is_stationary_22 <= io_in_c_bypass_19_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_0_data_22 <= io_in_c_bypass_20_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_0_is_stationary_22 <= io_in_c_bypass_20_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_1_data_22 <= io_in_c_bypass_20_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_1_is_stationary_22 <= io_in_c_bypass_20_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_2_data_22 <= io_in_c_bypass_20_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_2_is_stationary_22 <= io_in_c_bypass_20_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_3_data_22 <= io_in_c_bypass_20_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_3_is_stationary_22 <= io_in_c_bypass_20_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_0_data_22 <= io_in_c_bypass_21_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_0_is_stationary_22 <= io_in_c_bypass_21_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_1_data_22 <= io_in_c_bypass_21_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_1_is_stationary_22 <= io_in_c_bypass_21_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_2_data_22 <= io_in_c_bypass_21_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_2_is_stationary_22 <= io_in_c_bypass_21_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_3_data_22 <= io_in_c_bypass_21_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_3_is_stationary_22 <= io_in_c_bypass_21_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_0_data_22 <= io_in_c_bypass_22_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_0_is_stationary_22 <= io_in_c_bypass_22_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_1_data_22 <= io_in_c_bypass_22_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_1_is_stationary_22 <= io_in_c_bypass_22_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_2_data_22 <= io_in_c_bypass_22_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_2_is_stationary_22 <= io_in_c_bypass_22_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_3_data_22 <= io_in_c_bypass_22_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_3_is_stationary_22 <= io_in_c_bypass_22_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_0_data_22 <= io_in_c_bypass_23_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_0_is_stationary_22 <= io_in_c_bypass_23_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_1_data_22 <= io_in_c_bypass_23_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_1_is_stationary_22 <= io_in_c_bypass_23_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_2_data_22 <= io_in_c_bypass_23_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_2_is_stationary_22 <= io_in_c_bypass_23_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_3_data_22 <= io_in_c_bypass_23_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_3_is_stationary_22 <= io_in_c_bypass_23_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_0_data_22 <= io_in_c_bypass_24_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_0_is_stationary_22 <= io_in_c_bypass_24_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_1_data_22 <= io_in_c_bypass_24_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_1_is_stationary_22 <= io_in_c_bypass_24_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_2_data_22 <= io_in_c_bypass_24_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_2_is_stationary_22 <= io_in_c_bypass_24_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_3_data_22 <= io_in_c_bypass_24_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_3_is_stationary_22 <= io_in_c_bypass_24_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_0_data_22 <= io_in_c_bypass_25_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_0_is_stationary_22 <= io_in_c_bypass_25_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_1_data_22 <= io_in_c_bypass_25_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_1_is_stationary_22 <= io_in_c_bypass_25_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_2_data_22 <= io_in_c_bypass_25_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_2_is_stationary_22 <= io_in_c_bypass_25_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_3_data_22 <= io_in_c_bypass_25_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_3_is_stationary_22 <= io_in_c_bypass_25_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_0_data_22 <= io_in_c_bypass_26_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_0_is_stationary_22 <= io_in_c_bypass_26_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_1_data_22 <= io_in_c_bypass_26_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_1_is_stationary_22 <= io_in_c_bypass_26_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_2_data_22 <= io_in_c_bypass_26_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_2_is_stationary_22 <= io_in_c_bypass_26_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_3_data_22 <= io_in_c_bypass_26_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_3_is_stationary_22 <= io_in_c_bypass_26_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_0_data_22 <= io_in_c_bypass_27_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_0_is_stationary_22 <= io_in_c_bypass_27_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_1_data_22 <= io_in_c_bypass_27_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_1_is_stationary_22 <= io_in_c_bypass_27_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_2_data_22 <= io_in_c_bypass_27_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_2_is_stationary_22 <= io_in_c_bypass_27_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_3_data_22 <= io_in_c_bypass_27_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_3_is_stationary_22 <= io_in_c_bypass_27_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_0_data_22 <= io_in_c_bypass_28_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_0_is_stationary_22 <= io_in_c_bypass_28_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_1_data_22 <= io_in_c_bypass_28_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_1_is_stationary_22 <= io_in_c_bypass_28_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_2_data_22 <= io_in_c_bypass_28_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_2_is_stationary_22 <= io_in_c_bypass_28_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_3_data_22 <= io_in_c_bypass_28_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_3_is_stationary_22 <= io_in_c_bypass_28_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_0_data_22 <= io_in_c_bypass_29_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_0_is_stationary_22 <= io_in_c_bypass_29_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_1_data_22 <= io_in_c_bypass_29_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_1_is_stationary_22 <= io_in_c_bypass_29_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_2_data_22 <= io_in_c_bypass_29_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_2_is_stationary_22 <= io_in_c_bypass_29_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_3_data_22 <= io_in_c_bypass_29_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_3_is_stationary_22 <= io_in_c_bypass_29_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_0_data_22 <= io_in_c_bypass_30_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_0_is_stationary_22 <= io_in_c_bypass_30_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_1_data_22 <= io_in_c_bypass_30_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_1_is_stationary_22 <= io_in_c_bypass_30_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_2_data_22 <= io_in_c_bypass_30_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_2_is_stationary_22 <= io_in_c_bypass_30_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_3_data_22 <= io_in_c_bypass_30_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_3_is_stationary_22 <= io_in_c_bypass_30_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_0_data_22 <= io_in_c_bypass_31_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_0_is_stationary_22 <= io_in_c_bypass_31_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_1_data_22 <= io_in_c_bypass_31_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_1_is_stationary_22 <= io_in_c_bypass_31_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_2_data_22 <= io_in_c_bypass_31_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_2_is_stationary_22 <= io_in_c_bypass_31_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_3_data_22 <= io_in_c_bypass_31_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_3_is_stationary_22 <= io_in_c_bypass_31_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_0_data_23 <= io_in_c_bypass_0_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_0_is_stationary_23 <= io_in_c_bypass_0_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_1_data_23 <= io_in_c_bypass_0_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_1_is_stationary_23 <= io_in_c_bypass_0_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_2_data_23 <= io_in_c_bypass_0_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_2_is_stationary_23 <= io_in_c_bypass_0_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_3_data_23 <= io_in_c_bypass_0_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_3_is_stationary_23 <= io_in_c_bypass_0_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_0_data_23 <= io_in_c_bypass_1_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_0_is_stationary_23 <= io_in_c_bypass_1_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_1_data_23 <= io_in_c_bypass_1_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_1_is_stationary_23 <= io_in_c_bypass_1_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_2_data_23 <= io_in_c_bypass_1_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_2_is_stationary_23 <= io_in_c_bypass_1_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_3_data_23 <= io_in_c_bypass_1_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_3_is_stationary_23 <= io_in_c_bypass_1_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_0_data_23 <= io_in_c_bypass_2_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_0_is_stationary_23 <= io_in_c_bypass_2_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_1_data_23 <= io_in_c_bypass_2_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_1_is_stationary_23 <= io_in_c_bypass_2_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_2_data_23 <= io_in_c_bypass_2_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_2_is_stationary_23 <= io_in_c_bypass_2_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_3_data_23 <= io_in_c_bypass_2_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_3_is_stationary_23 <= io_in_c_bypass_2_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_0_data_23 <= io_in_c_bypass_3_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_0_is_stationary_23 <= io_in_c_bypass_3_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_1_data_23 <= io_in_c_bypass_3_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_1_is_stationary_23 <= io_in_c_bypass_3_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_2_data_23 <= io_in_c_bypass_3_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_2_is_stationary_23 <= io_in_c_bypass_3_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_3_data_23 <= io_in_c_bypass_3_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_3_is_stationary_23 <= io_in_c_bypass_3_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_0_data_23 <= io_in_c_bypass_4_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_0_is_stationary_23 <= io_in_c_bypass_4_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_1_data_23 <= io_in_c_bypass_4_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_1_is_stationary_23 <= io_in_c_bypass_4_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_2_data_23 <= io_in_c_bypass_4_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_2_is_stationary_23 <= io_in_c_bypass_4_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_3_data_23 <= io_in_c_bypass_4_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_3_is_stationary_23 <= io_in_c_bypass_4_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_0_data_23 <= io_in_c_bypass_5_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_0_is_stationary_23 <= io_in_c_bypass_5_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_1_data_23 <= io_in_c_bypass_5_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_1_is_stationary_23 <= io_in_c_bypass_5_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_2_data_23 <= io_in_c_bypass_5_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_2_is_stationary_23 <= io_in_c_bypass_5_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_3_data_23 <= io_in_c_bypass_5_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_3_is_stationary_23 <= io_in_c_bypass_5_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_0_data_23 <= io_in_c_bypass_6_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_0_is_stationary_23 <= io_in_c_bypass_6_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_1_data_23 <= io_in_c_bypass_6_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_1_is_stationary_23 <= io_in_c_bypass_6_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_2_data_23 <= io_in_c_bypass_6_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_2_is_stationary_23 <= io_in_c_bypass_6_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_3_data_23 <= io_in_c_bypass_6_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_3_is_stationary_23 <= io_in_c_bypass_6_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_0_data_23 <= io_in_c_bypass_7_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_0_is_stationary_23 <= io_in_c_bypass_7_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_1_data_23 <= io_in_c_bypass_7_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_1_is_stationary_23 <= io_in_c_bypass_7_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_2_data_23 <= io_in_c_bypass_7_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_2_is_stationary_23 <= io_in_c_bypass_7_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_3_data_23 <= io_in_c_bypass_7_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_3_is_stationary_23 <= io_in_c_bypass_7_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_0_data_23 <= io_in_c_bypass_8_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_0_is_stationary_23 <= io_in_c_bypass_8_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_1_data_23 <= io_in_c_bypass_8_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_1_is_stationary_23 <= io_in_c_bypass_8_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_2_data_23 <= io_in_c_bypass_8_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_2_is_stationary_23 <= io_in_c_bypass_8_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_3_data_23 <= io_in_c_bypass_8_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_3_is_stationary_23 <= io_in_c_bypass_8_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_0_data_23 <= io_in_c_bypass_9_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_0_is_stationary_23 <= io_in_c_bypass_9_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_1_data_23 <= io_in_c_bypass_9_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_1_is_stationary_23 <= io_in_c_bypass_9_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_2_data_23 <= io_in_c_bypass_9_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_2_is_stationary_23 <= io_in_c_bypass_9_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_3_data_23 <= io_in_c_bypass_9_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_3_is_stationary_23 <= io_in_c_bypass_9_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_0_data_23 <= io_in_c_bypass_10_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_0_is_stationary_23 <= io_in_c_bypass_10_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_1_data_23 <= io_in_c_bypass_10_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_1_is_stationary_23 <= io_in_c_bypass_10_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_2_data_23 <= io_in_c_bypass_10_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_2_is_stationary_23 <= io_in_c_bypass_10_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_3_data_23 <= io_in_c_bypass_10_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_3_is_stationary_23 <= io_in_c_bypass_10_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_0_data_23 <= io_in_c_bypass_11_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_0_is_stationary_23 <= io_in_c_bypass_11_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_1_data_23 <= io_in_c_bypass_11_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_1_is_stationary_23 <= io_in_c_bypass_11_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_2_data_23 <= io_in_c_bypass_11_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_2_is_stationary_23 <= io_in_c_bypass_11_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_3_data_23 <= io_in_c_bypass_11_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_3_is_stationary_23 <= io_in_c_bypass_11_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_0_data_23 <= io_in_c_bypass_12_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_0_is_stationary_23 <= io_in_c_bypass_12_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_1_data_23 <= io_in_c_bypass_12_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_1_is_stationary_23 <= io_in_c_bypass_12_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_2_data_23 <= io_in_c_bypass_12_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_2_is_stationary_23 <= io_in_c_bypass_12_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_3_data_23 <= io_in_c_bypass_12_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_3_is_stationary_23 <= io_in_c_bypass_12_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_0_data_23 <= io_in_c_bypass_13_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_0_is_stationary_23 <= io_in_c_bypass_13_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_1_data_23 <= io_in_c_bypass_13_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_1_is_stationary_23 <= io_in_c_bypass_13_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_2_data_23 <= io_in_c_bypass_13_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_2_is_stationary_23 <= io_in_c_bypass_13_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_3_data_23 <= io_in_c_bypass_13_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_3_is_stationary_23 <= io_in_c_bypass_13_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_0_data_23 <= io_in_c_bypass_14_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_0_is_stationary_23 <= io_in_c_bypass_14_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_1_data_23 <= io_in_c_bypass_14_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_1_is_stationary_23 <= io_in_c_bypass_14_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_2_data_23 <= io_in_c_bypass_14_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_2_is_stationary_23 <= io_in_c_bypass_14_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_3_data_23 <= io_in_c_bypass_14_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_3_is_stationary_23 <= io_in_c_bypass_14_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_0_data_23 <= io_in_c_bypass_15_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_0_is_stationary_23 <= io_in_c_bypass_15_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_1_data_23 <= io_in_c_bypass_15_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_1_is_stationary_23 <= io_in_c_bypass_15_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_2_data_23 <= io_in_c_bypass_15_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_2_is_stationary_23 <= io_in_c_bypass_15_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_3_data_23 <= io_in_c_bypass_15_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_3_is_stationary_23 <= io_in_c_bypass_15_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_0_data_23 <= io_in_c_bypass_16_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_0_is_stationary_23 <= io_in_c_bypass_16_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_1_data_23 <= io_in_c_bypass_16_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_1_is_stationary_23 <= io_in_c_bypass_16_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_2_data_23 <= io_in_c_bypass_16_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_2_is_stationary_23 <= io_in_c_bypass_16_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_3_data_23 <= io_in_c_bypass_16_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_3_is_stationary_23 <= io_in_c_bypass_16_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_0_data_23 <= io_in_c_bypass_17_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_0_is_stationary_23 <= io_in_c_bypass_17_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_1_data_23 <= io_in_c_bypass_17_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_1_is_stationary_23 <= io_in_c_bypass_17_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_2_data_23 <= io_in_c_bypass_17_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_2_is_stationary_23 <= io_in_c_bypass_17_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_3_data_23 <= io_in_c_bypass_17_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_3_is_stationary_23 <= io_in_c_bypass_17_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_0_data_23 <= io_in_c_bypass_18_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_0_is_stationary_23 <= io_in_c_bypass_18_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_1_data_23 <= io_in_c_bypass_18_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_1_is_stationary_23 <= io_in_c_bypass_18_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_2_data_23 <= io_in_c_bypass_18_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_2_is_stationary_23 <= io_in_c_bypass_18_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_3_data_23 <= io_in_c_bypass_18_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_3_is_stationary_23 <= io_in_c_bypass_18_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_0_data_23 <= io_in_c_bypass_19_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_0_is_stationary_23 <= io_in_c_bypass_19_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_1_data_23 <= io_in_c_bypass_19_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_1_is_stationary_23 <= io_in_c_bypass_19_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_2_data_23 <= io_in_c_bypass_19_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_2_is_stationary_23 <= io_in_c_bypass_19_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_3_data_23 <= io_in_c_bypass_19_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_3_is_stationary_23 <= io_in_c_bypass_19_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_0_data_23 <= io_in_c_bypass_20_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_0_is_stationary_23 <= io_in_c_bypass_20_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_1_data_23 <= io_in_c_bypass_20_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_1_is_stationary_23 <= io_in_c_bypass_20_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_2_data_23 <= io_in_c_bypass_20_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_2_is_stationary_23 <= io_in_c_bypass_20_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_3_data_23 <= io_in_c_bypass_20_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_3_is_stationary_23 <= io_in_c_bypass_20_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_0_data_23 <= io_in_c_bypass_21_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_0_is_stationary_23 <= io_in_c_bypass_21_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_1_data_23 <= io_in_c_bypass_21_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_1_is_stationary_23 <= io_in_c_bypass_21_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_2_data_23 <= io_in_c_bypass_21_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_2_is_stationary_23 <= io_in_c_bypass_21_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_3_data_23 <= io_in_c_bypass_21_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_3_is_stationary_23 <= io_in_c_bypass_21_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_0_data_23 <= io_in_c_bypass_22_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_0_is_stationary_23 <= io_in_c_bypass_22_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_1_data_23 <= io_in_c_bypass_22_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_1_is_stationary_23 <= io_in_c_bypass_22_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_2_data_23 <= io_in_c_bypass_22_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_2_is_stationary_23 <= io_in_c_bypass_22_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_3_data_23 <= io_in_c_bypass_22_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_3_is_stationary_23 <= io_in_c_bypass_22_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_0_data_23 <= io_in_c_bypass_23_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_0_is_stationary_23 <= io_in_c_bypass_23_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_1_data_23 <= io_in_c_bypass_23_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_1_is_stationary_23 <= io_in_c_bypass_23_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_2_data_23 <= io_in_c_bypass_23_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_2_is_stationary_23 <= io_in_c_bypass_23_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_3_data_23 <= io_in_c_bypass_23_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_3_is_stationary_23 <= io_in_c_bypass_23_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_0_data_23 <= io_in_c_bypass_24_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_0_is_stationary_23 <= io_in_c_bypass_24_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_1_data_23 <= io_in_c_bypass_24_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_1_is_stationary_23 <= io_in_c_bypass_24_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_2_data_23 <= io_in_c_bypass_24_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_2_is_stationary_23 <= io_in_c_bypass_24_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_3_data_23 <= io_in_c_bypass_24_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_3_is_stationary_23 <= io_in_c_bypass_24_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_0_data_23 <= io_in_c_bypass_25_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_0_is_stationary_23 <= io_in_c_bypass_25_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_1_data_23 <= io_in_c_bypass_25_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_1_is_stationary_23 <= io_in_c_bypass_25_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_2_data_23 <= io_in_c_bypass_25_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_2_is_stationary_23 <= io_in_c_bypass_25_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_3_data_23 <= io_in_c_bypass_25_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_3_is_stationary_23 <= io_in_c_bypass_25_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_0_data_23 <= io_in_c_bypass_26_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_0_is_stationary_23 <= io_in_c_bypass_26_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_1_data_23 <= io_in_c_bypass_26_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_1_is_stationary_23 <= io_in_c_bypass_26_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_2_data_23 <= io_in_c_bypass_26_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_2_is_stationary_23 <= io_in_c_bypass_26_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_3_data_23 <= io_in_c_bypass_26_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_3_is_stationary_23 <= io_in_c_bypass_26_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_0_data_23 <= io_in_c_bypass_27_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_0_is_stationary_23 <= io_in_c_bypass_27_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_1_data_23 <= io_in_c_bypass_27_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_1_is_stationary_23 <= io_in_c_bypass_27_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_2_data_23 <= io_in_c_bypass_27_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_2_is_stationary_23 <= io_in_c_bypass_27_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_3_data_23 <= io_in_c_bypass_27_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_3_is_stationary_23 <= io_in_c_bypass_27_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_0_data_23 <= io_in_c_bypass_28_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_0_is_stationary_23 <= io_in_c_bypass_28_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_1_data_23 <= io_in_c_bypass_28_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_1_is_stationary_23 <= io_in_c_bypass_28_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_2_data_23 <= io_in_c_bypass_28_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_2_is_stationary_23 <= io_in_c_bypass_28_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_3_data_23 <= io_in_c_bypass_28_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_3_is_stationary_23 <= io_in_c_bypass_28_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_0_data_23 <= io_in_c_bypass_29_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_0_is_stationary_23 <= io_in_c_bypass_29_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_1_data_23 <= io_in_c_bypass_29_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_1_is_stationary_23 <= io_in_c_bypass_29_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_2_data_23 <= io_in_c_bypass_29_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_2_is_stationary_23 <= io_in_c_bypass_29_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_3_data_23 <= io_in_c_bypass_29_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_3_is_stationary_23 <= io_in_c_bypass_29_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_0_data_23 <= io_in_c_bypass_30_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_0_is_stationary_23 <= io_in_c_bypass_30_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_1_data_23 <= io_in_c_bypass_30_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_1_is_stationary_23 <= io_in_c_bypass_30_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_2_data_23 <= io_in_c_bypass_30_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_2_is_stationary_23 <= io_in_c_bypass_30_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_3_data_23 <= io_in_c_bypass_30_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_3_is_stationary_23 <= io_in_c_bypass_30_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_0_data_23 <= io_in_c_bypass_31_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_0_is_stationary_23 <= io_in_c_bypass_31_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_1_data_23 <= io_in_c_bypass_31_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_1_is_stationary_23 <= io_in_c_bypass_31_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_2_data_23 <= io_in_c_bypass_31_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_2_is_stationary_23 <= io_in_c_bypass_31_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_3_data_23 <= io_in_c_bypass_31_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_3_is_stationary_23 <= io_in_c_bypass_31_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_0_data_24 <= io_in_c_bypass_0_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_0_is_stationary_24 <= io_in_c_bypass_0_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_1_data_24 <= io_in_c_bypass_0_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_1_is_stationary_24 <= io_in_c_bypass_0_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_2_data_24 <= io_in_c_bypass_0_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_2_is_stationary_24 <= io_in_c_bypass_0_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_3_data_24 <= io_in_c_bypass_0_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_3_is_stationary_24 <= io_in_c_bypass_0_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_0_data_24 <= io_in_c_bypass_1_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_0_is_stationary_24 <= io_in_c_bypass_1_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_1_data_24 <= io_in_c_bypass_1_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_1_is_stationary_24 <= io_in_c_bypass_1_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_2_data_24 <= io_in_c_bypass_1_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_2_is_stationary_24 <= io_in_c_bypass_1_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_3_data_24 <= io_in_c_bypass_1_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_3_is_stationary_24 <= io_in_c_bypass_1_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_0_data_24 <= io_in_c_bypass_2_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_0_is_stationary_24 <= io_in_c_bypass_2_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_1_data_24 <= io_in_c_bypass_2_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_1_is_stationary_24 <= io_in_c_bypass_2_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_2_data_24 <= io_in_c_bypass_2_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_2_is_stationary_24 <= io_in_c_bypass_2_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_3_data_24 <= io_in_c_bypass_2_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_3_is_stationary_24 <= io_in_c_bypass_2_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_0_data_24 <= io_in_c_bypass_3_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_0_is_stationary_24 <= io_in_c_bypass_3_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_1_data_24 <= io_in_c_bypass_3_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_1_is_stationary_24 <= io_in_c_bypass_3_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_2_data_24 <= io_in_c_bypass_3_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_2_is_stationary_24 <= io_in_c_bypass_3_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_3_data_24 <= io_in_c_bypass_3_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_3_is_stationary_24 <= io_in_c_bypass_3_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_0_data_24 <= io_in_c_bypass_4_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_0_is_stationary_24 <= io_in_c_bypass_4_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_1_data_24 <= io_in_c_bypass_4_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_1_is_stationary_24 <= io_in_c_bypass_4_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_2_data_24 <= io_in_c_bypass_4_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_2_is_stationary_24 <= io_in_c_bypass_4_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_3_data_24 <= io_in_c_bypass_4_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_3_is_stationary_24 <= io_in_c_bypass_4_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_0_data_24 <= io_in_c_bypass_5_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_0_is_stationary_24 <= io_in_c_bypass_5_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_1_data_24 <= io_in_c_bypass_5_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_1_is_stationary_24 <= io_in_c_bypass_5_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_2_data_24 <= io_in_c_bypass_5_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_2_is_stationary_24 <= io_in_c_bypass_5_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_3_data_24 <= io_in_c_bypass_5_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_3_is_stationary_24 <= io_in_c_bypass_5_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_0_data_24 <= io_in_c_bypass_6_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_0_is_stationary_24 <= io_in_c_bypass_6_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_1_data_24 <= io_in_c_bypass_6_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_1_is_stationary_24 <= io_in_c_bypass_6_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_2_data_24 <= io_in_c_bypass_6_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_2_is_stationary_24 <= io_in_c_bypass_6_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_3_data_24 <= io_in_c_bypass_6_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_3_is_stationary_24 <= io_in_c_bypass_6_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_0_data_24 <= io_in_c_bypass_7_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_0_is_stationary_24 <= io_in_c_bypass_7_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_1_data_24 <= io_in_c_bypass_7_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_1_is_stationary_24 <= io_in_c_bypass_7_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_2_data_24 <= io_in_c_bypass_7_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_2_is_stationary_24 <= io_in_c_bypass_7_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_3_data_24 <= io_in_c_bypass_7_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_3_is_stationary_24 <= io_in_c_bypass_7_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_0_data_24 <= io_in_c_bypass_8_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_0_is_stationary_24 <= io_in_c_bypass_8_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_1_data_24 <= io_in_c_bypass_8_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_1_is_stationary_24 <= io_in_c_bypass_8_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_2_data_24 <= io_in_c_bypass_8_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_2_is_stationary_24 <= io_in_c_bypass_8_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_3_data_24 <= io_in_c_bypass_8_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_3_is_stationary_24 <= io_in_c_bypass_8_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_0_data_24 <= io_in_c_bypass_9_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_0_is_stationary_24 <= io_in_c_bypass_9_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_1_data_24 <= io_in_c_bypass_9_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_1_is_stationary_24 <= io_in_c_bypass_9_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_2_data_24 <= io_in_c_bypass_9_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_2_is_stationary_24 <= io_in_c_bypass_9_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_3_data_24 <= io_in_c_bypass_9_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_3_is_stationary_24 <= io_in_c_bypass_9_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_0_data_24 <= io_in_c_bypass_10_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_0_is_stationary_24 <= io_in_c_bypass_10_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_1_data_24 <= io_in_c_bypass_10_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_1_is_stationary_24 <= io_in_c_bypass_10_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_2_data_24 <= io_in_c_bypass_10_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_2_is_stationary_24 <= io_in_c_bypass_10_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_3_data_24 <= io_in_c_bypass_10_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_3_is_stationary_24 <= io_in_c_bypass_10_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_0_data_24 <= io_in_c_bypass_11_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_0_is_stationary_24 <= io_in_c_bypass_11_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_1_data_24 <= io_in_c_bypass_11_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_1_is_stationary_24 <= io_in_c_bypass_11_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_2_data_24 <= io_in_c_bypass_11_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_2_is_stationary_24 <= io_in_c_bypass_11_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_3_data_24 <= io_in_c_bypass_11_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_3_is_stationary_24 <= io_in_c_bypass_11_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_0_data_24 <= io_in_c_bypass_12_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_0_is_stationary_24 <= io_in_c_bypass_12_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_1_data_24 <= io_in_c_bypass_12_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_1_is_stationary_24 <= io_in_c_bypass_12_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_2_data_24 <= io_in_c_bypass_12_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_2_is_stationary_24 <= io_in_c_bypass_12_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_3_data_24 <= io_in_c_bypass_12_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_3_is_stationary_24 <= io_in_c_bypass_12_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_0_data_24 <= io_in_c_bypass_13_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_0_is_stationary_24 <= io_in_c_bypass_13_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_1_data_24 <= io_in_c_bypass_13_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_1_is_stationary_24 <= io_in_c_bypass_13_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_2_data_24 <= io_in_c_bypass_13_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_2_is_stationary_24 <= io_in_c_bypass_13_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_3_data_24 <= io_in_c_bypass_13_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_3_is_stationary_24 <= io_in_c_bypass_13_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_0_data_24 <= io_in_c_bypass_14_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_0_is_stationary_24 <= io_in_c_bypass_14_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_1_data_24 <= io_in_c_bypass_14_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_1_is_stationary_24 <= io_in_c_bypass_14_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_2_data_24 <= io_in_c_bypass_14_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_2_is_stationary_24 <= io_in_c_bypass_14_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_3_data_24 <= io_in_c_bypass_14_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_3_is_stationary_24 <= io_in_c_bypass_14_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_0_data_24 <= io_in_c_bypass_15_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_0_is_stationary_24 <= io_in_c_bypass_15_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_1_data_24 <= io_in_c_bypass_15_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_1_is_stationary_24 <= io_in_c_bypass_15_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_2_data_24 <= io_in_c_bypass_15_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_2_is_stationary_24 <= io_in_c_bypass_15_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_3_data_24 <= io_in_c_bypass_15_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_3_is_stationary_24 <= io_in_c_bypass_15_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_0_data_24 <= io_in_c_bypass_16_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_0_is_stationary_24 <= io_in_c_bypass_16_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_1_data_24 <= io_in_c_bypass_16_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_1_is_stationary_24 <= io_in_c_bypass_16_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_2_data_24 <= io_in_c_bypass_16_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_2_is_stationary_24 <= io_in_c_bypass_16_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_3_data_24 <= io_in_c_bypass_16_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_3_is_stationary_24 <= io_in_c_bypass_16_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_0_data_24 <= io_in_c_bypass_17_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_0_is_stationary_24 <= io_in_c_bypass_17_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_1_data_24 <= io_in_c_bypass_17_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_1_is_stationary_24 <= io_in_c_bypass_17_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_2_data_24 <= io_in_c_bypass_17_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_2_is_stationary_24 <= io_in_c_bypass_17_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_3_data_24 <= io_in_c_bypass_17_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_3_is_stationary_24 <= io_in_c_bypass_17_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_0_data_24 <= io_in_c_bypass_18_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_0_is_stationary_24 <= io_in_c_bypass_18_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_1_data_24 <= io_in_c_bypass_18_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_1_is_stationary_24 <= io_in_c_bypass_18_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_2_data_24 <= io_in_c_bypass_18_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_2_is_stationary_24 <= io_in_c_bypass_18_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_3_data_24 <= io_in_c_bypass_18_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_3_is_stationary_24 <= io_in_c_bypass_18_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_0_data_24 <= io_in_c_bypass_19_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_0_is_stationary_24 <= io_in_c_bypass_19_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_1_data_24 <= io_in_c_bypass_19_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_1_is_stationary_24 <= io_in_c_bypass_19_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_2_data_24 <= io_in_c_bypass_19_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_2_is_stationary_24 <= io_in_c_bypass_19_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_3_data_24 <= io_in_c_bypass_19_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_3_is_stationary_24 <= io_in_c_bypass_19_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_0_data_24 <= io_in_c_bypass_20_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_0_is_stationary_24 <= io_in_c_bypass_20_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_1_data_24 <= io_in_c_bypass_20_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_1_is_stationary_24 <= io_in_c_bypass_20_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_2_data_24 <= io_in_c_bypass_20_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_2_is_stationary_24 <= io_in_c_bypass_20_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_3_data_24 <= io_in_c_bypass_20_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_3_is_stationary_24 <= io_in_c_bypass_20_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_0_data_24 <= io_in_c_bypass_21_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_0_is_stationary_24 <= io_in_c_bypass_21_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_1_data_24 <= io_in_c_bypass_21_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_1_is_stationary_24 <= io_in_c_bypass_21_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_2_data_24 <= io_in_c_bypass_21_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_2_is_stationary_24 <= io_in_c_bypass_21_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_3_data_24 <= io_in_c_bypass_21_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_3_is_stationary_24 <= io_in_c_bypass_21_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_0_data_24 <= io_in_c_bypass_22_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_0_is_stationary_24 <= io_in_c_bypass_22_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_1_data_24 <= io_in_c_bypass_22_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_1_is_stationary_24 <= io_in_c_bypass_22_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_2_data_24 <= io_in_c_bypass_22_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_2_is_stationary_24 <= io_in_c_bypass_22_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_3_data_24 <= io_in_c_bypass_22_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_3_is_stationary_24 <= io_in_c_bypass_22_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_0_data_24 <= io_in_c_bypass_23_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_0_is_stationary_24 <= io_in_c_bypass_23_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_1_data_24 <= io_in_c_bypass_23_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_1_is_stationary_24 <= io_in_c_bypass_23_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_2_data_24 <= io_in_c_bypass_23_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_2_is_stationary_24 <= io_in_c_bypass_23_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_3_data_24 <= io_in_c_bypass_23_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_3_is_stationary_24 <= io_in_c_bypass_23_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_0_data_24 <= io_in_c_bypass_24_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_0_is_stationary_24 <= io_in_c_bypass_24_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_1_data_24 <= io_in_c_bypass_24_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_1_is_stationary_24 <= io_in_c_bypass_24_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_2_data_24 <= io_in_c_bypass_24_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_2_is_stationary_24 <= io_in_c_bypass_24_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_3_data_24 <= io_in_c_bypass_24_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_3_is_stationary_24 <= io_in_c_bypass_24_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_0_data_24 <= io_in_c_bypass_25_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_0_is_stationary_24 <= io_in_c_bypass_25_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_1_data_24 <= io_in_c_bypass_25_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_1_is_stationary_24 <= io_in_c_bypass_25_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_2_data_24 <= io_in_c_bypass_25_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_2_is_stationary_24 <= io_in_c_bypass_25_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_3_data_24 <= io_in_c_bypass_25_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_3_is_stationary_24 <= io_in_c_bypass_25_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_0_data_24 <= io_in_c_bypass_26_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_0_is_stationary_24 <= io_in_c_bypass_26_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_1_data_24 <= io_in_c_bypass_26_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_1_is_stationary_24 <= io_in_c_bypass_26_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_2_data_24 <= io_in_c_bypass_26_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_2_is_stationary_24 <= io_in_c_bypass_26_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_3_data_24 <= io_in_c_bypass_26_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_3_is_stationary_24 <= io_in_c_bypass_26_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_0_data_24 <= io_in_c_bypass_27_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_0_is_stationary_24 <= io_in_c_bypass_27_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_1_data_24 <= io_in_c_bypass_27_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_1_is_stationary_24 <= io_in_c_bypass_27_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_2_data_24 <= io_in_c_bypass_27_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_2_is_stationary_24 <= io_in_c_bypass_27_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_3_data_24 <= io_in_c_bypass_27_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_3_is_stationary_24 <= io_in_c_bypass_27_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_0_data_24 <= io_in_c_bypass_28_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_0_is_stationary_24 <= io_in_c_bypass_28_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_1_data_24 <= io_in_c_bypass_28_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_1_is_stationary_24 <= io_in_c_bypass_28_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_2_data_24 <= io_in_c_bypass_28_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_2_is_stationary_24 <= io_in_c_bypass_28_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_3_data_24 <= io_in_c_bypass_28_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_3_is_stationary_24 <= io_in_c_bypass_28_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_0_data_24 <= io_in_c_bypass_29_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_0_is_stationary_24 <= io_in_c_bypass_29_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_1_data_24 <= io_in_c_bypass_29_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_1_is_stationary_24 <= io_in_c_bypass_29_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_2_data_24 <= io_in_c_bypass_29_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_2_is_stationary_24 <= io_in_c_bypass_29_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_3_data_24 <= io_in_c_bypass_29_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_3_is_stationary_24 <= io_in_c_bypass_29_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_0_data_24 <= io_in_c_bypass_30_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_0_is_stationary_24 <= io_in_c_bypass_30_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_1_data_24 <= io_in_c_bypass_30_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_1_is_stationary_24 <= io_in_c_bypass_30_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_2_data_24 <= io_in_c_bypass_30_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_2_is_stationary_24 <= io_in_c_bypass_30_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_3_data_24 <= io_in_c_bypass_30_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_3_is_stationary_24 <= io_in_c_bypass_30_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_0_data_24 <= io_in_c_bypass_31_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_0_is_stationary_24 <= io_in_c_bypass_31_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_1_data_24 <= io_in_c_bypass_31_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_1_is_stationary_24 <= io_in_c_bypass_31_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_2_data_24 <= io_in_c_bypass_31_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_2_is_stationary_24 <= io_in_c_bypass_31_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_3_data_24 <= io_in_c_bypass_31_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_3_is_stationary_24 <= io_in_c_bypass_31_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_0_data_25 <= io_in_c_bypass_0_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_0_is_stationary_25 <= io_in_c_bypass_0_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_1_data_25 <= io_in_c_bypass_0_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_1_is_stationary_25 <= io_in_c_bypass_0_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_2_data_25 <= io_in_c_bypass_0_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_2_is_stationary_25 <= io_in_c_bypass_0_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_3_data_25 <= io_in_c_bypass_0_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_3_is_stationary_25 <= io_in_c_bypass_0_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_0_data_25 <= io_in_c_bypass_1_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_0_is_stationary_25 <= io_in_c_bypass_1_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_1_data_25 <= io_in_c_bypass_1_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_1_is_stationary_25 <= io_in_c_bypass_1_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_2_data_25 <= io_in_c_bypass_1_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_2_is_stationary_25 <= io_in_c_bypass_1_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_3_data_25 <= io_in_c_bypass_1_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_3_is_stationary_25 <= io_in_c_bypass_1_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_0_data_25 <= io_in_c_bypass_2_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_0_is_stationary_25 <= io_in_c_bypass_2_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_1_data_25 <= io_in_c_bypass_2_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_1_is_stationary_25 <= io_in_c_bypass_2_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_2_data_25 <= io_in_c_bypass_2_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_2_is_stationary_25 <= io_in_c_bypass_2_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_3_data_25 <= io_in_c_bypass_2_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_3_is_stationary_25 <= io_in_c_bypass_2_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_0_data_25 <= io_in_c_bypass_3_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_0_is_stationary_25 <= io_in_c_bypass_3_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_1_data_25 <= io_in_c_bypass_3_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_1_is_stationary_25 <= io_in_c_bypass_3_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_2_data_25 <= io_in_c_bypass_3_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_2_is_stationary_25 <= io_in_c_bypass_3_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_3_data_25 <= io_in_c_bypass_3_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_3_is_stationary_25 <= io_in_c_bypass_3_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_0_data_25 <= io_in_c_bypass_4_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_0_is_stationary_25 <= io_in_c_bypass_4_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_1_data_25 <= io_in_c_bypass_4_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_1_is_stationary_25 <= io_in_c_bypass_4_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_2_data_25 <= io_in_c_bypass_4_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_2_is_stationary_25 <= io_in_c_bypass_4_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_3_data_25 <= io_in_c_bypass_4_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_3_is_stationary_25 <= io_in_c_bypass_4_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_0_data_25 <= io_in_c_bypass_5_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_0_is_stationary_25 <= io_in_c_bypass_5_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_1_data_25 <= io_in_c_bypass_5_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_1_is_stationary_25 <= io_in_c_bypass_5_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_2_data_25 <= io_in_c_bypass_5_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_2_is_stationary_25 <= io_in_c_bypass_5_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_3_data_25 <= io_in_c_bypass_5_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_3_is_stationary_25 <= io_in_c_bypass_5_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_0_data_25 <= io_in_c_bypass_6_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_0_is_stationary_25 <= io_in_c_bypass_6_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_1_data_25 <= io_in_c_bypass_6_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_1_is_stationary_25 <= io_in_c_bypass_6_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_2_data_25 <= io_in_c_bypass_6_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_2_is_stationary_25 <= io_in_c_bypass_6_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_3_data_25 <= io_in_c_bypass_6_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_3_is_stationary_25 <= io_in_c_bypass_6_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_0_data_25 <= io_in_c_bypass_7_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_0_is_stationary_25 <= io_in_c_bypass_7_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_1_data_25 <= io_in_c_bypass_7_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_1_is_stationary_25 <= io_in_c_bypass_7_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_2_data_25 <= io_in_c_bypass_7_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_2_is_stationary_25 <= io_in_c_bypass_7_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_3_data_25 <= io_in_c_bypass_7_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_3_is_stationary_25 <= io_in_c_bypass_7_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_0_data_25 <= io_in_c_bypass_8_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_0_is_stationary_25 <= io_in_c_bypass_8_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_1_data_25 <= io_in_c_bypass_8_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_1_is_stationary_25 <= io_in_c_bypass_8_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_2_data_25 <= io_in_c_bypass_8_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_2_is_stationary_25 <= io_in_c_bypass_8_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_3_data_25 <= io_in_c_bypass_8_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_3_is_stationary_25 <= io_in_c_bypass_8_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_0_data_25 <= io_in_c_bypass_9_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_0_is_stationary_25 <= io_in_c_bypass_9_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_1_data_25 <= io_in_c_bypass_9_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_1_is_stationary_25 <= io_in_c_bypass_9_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_2_data_25 <= io_in_c_bypass_9_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_2_is_stationary_25 <= io_in_c_bypass_9_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_3_data_25 <= io_in_c_bypass_9_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_3_is_stationary_25 <= io_in_c_bypass_9_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_0_data_25 <= io_in_c_bypass_10_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_0_is_stationary_25 <= io_in_c_bypass_10_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_1_data_25 <= io_in_c_bypass_10_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_1_is_stationary_25 <= io_in_c_bypass_10_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_2_data_25 <= io_in_c_bypass_10_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_2_is_stationary_25 <= io_in_c_bypass_10_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_3_data_25 <= io_in_c_bypass_10_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_3_is_stationary_25 <= io_in_c_bypass_10_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_0_data_25 <= io_in_c_bypass_11_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_0_is_stationary_25 <= io_in_c_bypass_11_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_1_data_25 <= io_in_c_bypass_11_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_1_is_stationary_25 <= io_in_c_bypass_11_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_2_data_25 <= io_in_c_bypass_11_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_2_is_stationary_25 <= io_in_c_bypass_11_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_3_data_25 <= io_in_c_bypass_11_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_3_is_stationary_25 <= io_in_c_bypass_11_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_0_data_25 <= io_in_c_bypass_12_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_0_is_stationary_25 <= io_in_c_bypass_12_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_1_data_25 <= io_in_c_bypass_12_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_1_is_stationary_25 <= io_in_c_bypass_12_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_2_data_25 <= io_in_c_bypass_12_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_2_is_stationary_25 <= io_in_c_bypass_12_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_3_data_25 <= io_in_c_bypass_12_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_3_is_stationary_25 <= io_in_c_bypass_12_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_0_data_25 <= io_in_c_bypass_13_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_0_is_stationary_25 <= io_in_c_bypass_13_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_1_data_25 <= io_in_c_bypass_13_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_1_is_stationary_25 <= io_in_c_bypass_13_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_2_data_25 <= io_in_c_bypass_13_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_2_is_stationary_25 <= io_in_c_bypass_13_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_3_data_25 <= io_in_c_bypass_13_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_3_is_stationary_25 <= io_in_c_bypass_13_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_0_data_25 <= io_in_c_bypass_14_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_0_is_stationary_25 <= io_in_c_bypass_14_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_1_data_25 <= io_in_c_bypass_14_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_1_is_stationary_25 <= io_in_c_bypass_14_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_2_data_25 <= io_in_c_bypass_14_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_2_is_stationary_25 <= io_in_c_bypass_14_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_3_data_25 <= io_in_c_bypass_14_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_3_is_stationary_25 <= io_in_c_bypass_14_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_0_data_25 <= io_in_c_bypass_15_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_0_is_stationary_25 <= io_in_c_bypass_15_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_1_data_25 <= io_in_c_bypass_15_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_1_is_stationary_25 <= io_in_c_bypass_15_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_2_data_25 <= io_in_c_bypass_15_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_2_is_stationary_25 <= io_in_c_bypass_15_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_3_data_25 <= io_in_c_bypass_15_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_3_is_stationary_25 <= io_in_c_bypass_15_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_0_data_25 <= io_in_c_bypass_16_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_0_is_stationary_25 <= io_in_c_bypass_16_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_1_data_25 <= io_in_c_bypass_16_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_1_is_stationary_25 <= io_in_c_bypass_16_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_2_data_25 <= io_in_c_bypass_16_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_2_is_stationary_25 <= io_in_c_bypass_16_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_3_data_25 <= io_in_c_bypass_16_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_3_is_stationary_25 <= io_in_c_bypass_16_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_0_data_25 <= io_in_c_bypass_17_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_0_is_stationary_25 <= io_in_c_bypass_17_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_1_data_25 <= io_in_c_bypass_17_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_1_is_stationary_25 <= io_in_c_bypass_17_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_2_data_25 <= io_in_c_bypass_17_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_2_is_stationary_25 <= io_in_c_bypass_17_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_3_data_25 <= io_in_c_bypass_17_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_3_is_stationary_25 <= io_in_c_bypass_17_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_0_data_25 <= io_in_c_bypass_18_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_0_is_stationary_25 <= io_in_c_bypass_18_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_1_data_25 <= io_in_c_bypass_18_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_1_is_stationary_25 <= io_in_c_bypass_18_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_2_data_25 <= io_in_c_bypass_18_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_2_is_stationary_25 <= io_in_c_bypass_18_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_3_data_25 <= io_in_c_bypass_18_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_3_is_stationary_25 <= io_in_c_bypass_18_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_0_data_25 <= io_in_c_bypass_19_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_0_is_stationary_25 <= io_in_c_bypass_19_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_1_data_25 <= io_in_c_bypass_19_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_1_is_stationary_25 <= io_in_c_bypass_19_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_2_data_25 <= io_in_c_bypass_19_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_2_is_stationary_25 <= io_in_c_bypass_19_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_3_data_25 <= io_in_c_bypass_19_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_3_is_stationary_25 <= io_in_c_bypass_19_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_0_data_25 <= io_in_c_bypass_20_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_0_is_stationary_25 <= io_in_c_bypass_20_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_1_data_25 <= io_in_c_bypass_20_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_1_is_stationary_25 <= io_in_c_bypass_20_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_2_data_25 <= io_in_c_bypass_20_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_2_is_stationary_25 <= io_in_c_bypass_20_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_3_data_25 <= io_in_c_bypass_20_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_3_is_stationary_25 <= io_in_c_bypass_20_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_0_data_25 <= io_in_c_bypass_21_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_0_is_stationary_25 <= io_in_c_bypass_21_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_1_data_25 <= io_in_c_bypass_21_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_1_is_stationary_25 <= io_in_c_bypass_21_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_2_data_25 <= io_in_c_bypass_21_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_2_is_stationary_25 <= io_in_c_bypass_21_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_3_data_25 <= io_in_c_bypass_21_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_3_is_stationary_25 <= io_in_c_bypass_21_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_0_data_25 <= io_in_c_bypass_22_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_0_is_stationary_25 <= io_in_c_bypass_22_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_1_data_25 <= io_in_c_bypass_22_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_1_is_stationary_25 <= io_in_c_bypass_22_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_2_data_25 <= io_in_c_bypass_22_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_2_is_stationary_25 <= io_in_c_bypass_22_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_3_data_25 <= io_in_c_bypass_22_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_3_is_stationary_25 <= io_in_c_bypass_22_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_0_data_25 <= io_in_c_bypass_23_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_0_is_stationary_25 <= io_in_c_bypass_23_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_1_data_25 <= io_in_c_bypass_23_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_1_is_stationary_25 <= io_in_c_bypass_23_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_2_data_25 <= io_in_c_bypass_23_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_2_is_stationary_25 <= io_in_c_bypass_23_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_3_data_25 <= io_in_c_bypass_23_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_3_is_stationary_25 <= io_in_c_bypass_23_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_0_data_25 <= io_in_c_bypass_24_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_0_is_stationary_25 <= io_in_c_bypass_24_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_1_data_25 <= io_in_c_bypass_24_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_1_is_stationary_25 <= io_in_c_bypass_24_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_2_data_25 <= io_in_c_bypass_24_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_2_is_stationary_25 <= io_in_c_bypass_24_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_3_data_25 <= io_in_c_bypass_24_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_3_is_stationary_25 <= io_in_c_bypass_24_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_0_data_25 <= io_in_c_bypass_25_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_0_is_stationary_25 <= io_in_c_bypass_25_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_1_data_25 <= io_in_c_bypass_25_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_1_is_stationary_25 <= io_in_c_bypass_25_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_2_data_25 <= io_in_c_bypass_25_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_2_is_stationary_25 <= io_in_c_bypass_25_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_3_data_25 <= io_in_c_bypass_25_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_3_is_stationary_25 <= io_in_c_bypass_25_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_0_data_25 <= io_in_c_bypass_26_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_0_is_stationary_25 <= io_in_c_bypass_26_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_1_data_25 <= io_in_c_bypass_26_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_1_is_stationary_25 <= io_in_c_bypass_26_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_2_data_25 <= io_in_c_bypass_26_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_2_is_stationary_25 <= io_in_c_bypass_26_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_3_data_25 <= io_in_c_bypass_26_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_3_is_stationary_25 <= io_in_c_bypass_26_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_0_data_25 <= io_in_c_bypass_27_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_0_is_stationary_25 <= io_in_c_bypass_27_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_1_data_25 <= io_in_c_bypass_27_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_1_is_stationary_25 <= io_in_c_bypass_27_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_2_data_25 <= io_in_c_bypass_27_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_2_is_stationary_25 <= io_in_c_bypass_27_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_3_data_25 <= io_in_c_bypass_27_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_3_is_stationary_25 <= io_in_c_bypass_27_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_0_data_25 <= io_in_c_bypass_28_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_0_is_stationary_25 <= io_in_c_bypass_28_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_1_data_25 <= io_in_c_bypass_28_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_1_is_stationary_25 <= io_in_c_bypass_28_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_2_data_25 <= io_in_c_bypass_28_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_2_is_stationary_25 <= io_in_c_bypass_28_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_3_data_25 <= io_in_c_bypass_28_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_3_is_stationary_25 <= io_in_c_bypass_28_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_0_data_25 <= io_in_c_bypass_29_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_0_is_stationary_25 <= io_in_c_bypass_29_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_1_data_25 <= io_in_c_bypass_29_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_1_is_stationary_25 <= io_in_c_bypass_29_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_2_data_25 <= io_in_c_bypass_29_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_2_is_stationary_25 <= io_in_c_bypass_29_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_3_data_25 <= io_in_c_bypass_29_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_3_is_stationary_25 <= io_in_c_bypass_29_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_0_data_25 <= io_in_c_bypass_30_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_0_is_stationary_25 <= io_in_c_bypass_30_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_1_data_25 <= io_in_c_bypass_30_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_1_is_stationary_25 <= io_in_c_bypass_30_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_2_data_25 <= io_in_c_bypass_30_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_2_is_stationary_25 <= io_in_c_bypass_30_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_3_data_25 <= io_in_c_bypass_30_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_3_is_stationary_25 <= io_in_c_bypass_30_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_0_data_25 <= io_in_c_bypass_31_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_0_is_stationary_25 <= io_in_c_bypass_31_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_1_data_25 <= io_in_c_bypass_31_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_1_is_stationary_25 <= io_in_c_bypass_31_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_2_data_25 <= io_in_c_bypass_31_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_2_is_stationary_25 <= io_in_c_bypass_31_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_3_data_25 <= io_in_c_bypass_31_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_3_is_stationary_25 <= io_in_c_bypass_31_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_0_data_26 <= io_in_c_bypass_0_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_0_is_stationary_26 <= io_in_c_bypass_0_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_1_data_26 <= io_in_c_bypass_0_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_1_is_stationary_26 <= io_in_c_bypass_0_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_2_data_26 <= io_in_c_bypass_0_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_2_is_stationary_26 <= io_in_c_bypass_0_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_3_data_26 <= io_in_c_bypass_0_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_3_is_stationary_26 <= io_in_c_bypass_0_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_0_data_26 <= io_in_c_bypass_1_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_0_is_stationary_26 <= io_in_c_bypass_1_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_1_data_26 <= io_in_c_bypass_1_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_1_is_stationary_26 <= io_in_c_bypass_1_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_2_data_26 <= io_in_c_bypass_1_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_2_is_stationary_26 <= io_in_c_bypass_1_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_3_data_26 <= io_in_c_bypass_1_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_3_is_stationary_26 <= io_in_c_bypass_1_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_0_data_26 <= io_in_c_bypass_2_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_0_is_stationary_26 <= io_in_c_bypass_2_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_1_data_26 <= io_in_c_bypass_2_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_1_is_stationary_26 <= io_in_c_bypass_2_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_2_data_26 <= io_in_c_bypass_2_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_2_is_stationary_26 <= io_in_c_bypass_2_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_3_data_26 <= io_in_c_bypass_2_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_3_is_stationary_26 <= io_in_c_bypass_2_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_0_data_26 <= io_in_c_bypass_3_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_0_is_stationary_26 <= io_in_c_bypass_3_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_1_data_26 <= io_in_c_bypass_3_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_1_is_stationary_26 <= io_in_c_bypass_3_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_2_data_26 <= io_in_c_bypass_3_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_2_is_stationary_26 <= io_in_c_bypass_3_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_3_data_26 <= io_in_c_bypass_3_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_3_is_stationary_26 <= io_in_c_bypass_3_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_0_data_26 <= io_in_c_bypass_4_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_0_is_stationary_26 <= io_in_c_bypass_4_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_1_data_26 <= io_in_c_bypass_4_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_1_is_stationary_26 <= io_in_c_bypass_4_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_2_data_26 <= io_in_c_bypass_4_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_2_is_stationary_26 <= io_in_c_bypass_4_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_3_data_26 <= io_in_c_bypass_4_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_3_is_stationary_26 <= io_in_c_bypass_4_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_0_data_26 <= io_in_c_bypass_5_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_0_is_stationary_26 <= io_in_c_bypass_5_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_1_data_26 <= io_in_c_bypass_5_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_1_is_stationary_26 <= io_in_c_bypass_5_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_2_data_26 <= io_in_c_bypass_5_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_2_is_stationary_26 <= io_in_c_bypass_5_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_3_data_26 <= io_in_c_bypass_5_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_3_is_stationary_26 <= io_in_c_bypass_5_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_0_data_26 <= io_in_c_bypass_6_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_0_is_stationary_26 <= io_in_c_bypass_6_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_1_data_26 <= io_in_c_bypass_6_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_1_is_stationary_26 <= io_in_c_bypass_6_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_2_data_26 <= io_in_c_bypass_6_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_2_is_stationary_26 <= io_in_c_bypass_6_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_3_data_26 <= io_in_c_bypass_6_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_3_is_stationary_26 <= io_in_c_bypass_6_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_0_data_26 <= io_in_c_bypass_7_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_0_is_stationary_26 <= io_in_c_bypass_7_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_1_data_26 <= io_in_c_bypass_7_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_1_is_stationary_26 <= io_in_c_bypass_7_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_2_data_26 <= io_in_c_bypass_7_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_2_is_stationary_26 <= io_in_c_bypass_7_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_3_data_26 <= io_in_c_bypass_7_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_3_is_stationary_26 <= io_in_c_bypass_7_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_0_data_26 <= io_in_c_bypass_8_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_0_is_stationary_26 <= io_in_c_bypass_8_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_1_data_26 <= io_in_c_bypass_8_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_1_is_stationary_26 <= io_in_c_bypass_8_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_2_data_26 <= io_in_c_bypass_8_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_2_is_stationary_26 <= io_in_c_bypass_8_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_3_data_26 <= io_in_c_bypass_8_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_3_is_stationary_26 <= io_in_c_bypass_8_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_0_data_26 <= io_in_c_bypass_9_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_0_is_stationary_26 <= io_in_c_bypass_9_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_1_data_26 <= io_in_c_bypass_9_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_1_is_stationary_26 <= io_in_c_bypass_9_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_2_data_26 <= io_in_c_bypass_9_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_2_is_stationary_26 <= io_in_c_bypass_9_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_3_data_26 <= io_in_c_bypass_9_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_3_is_stationary_26 <= io_in_c_bypass_9_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_0_data_26 <= io_in_c_bypass_10_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_0_is_stationary_26 <= io_in_c_bypass_10_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_1_data_26 <= io_in_c_bypass_10_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_1_is_stationary_26 <= io_in_c_bypass_10_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_2_data_26 <= io_in_c_bypass_10_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_2_is_stationary_26 <= io_in_c_bypass_10_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_3_data_26 <= io_in_c_bypass_10_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_3_is_stationary_26 <= io_in_c_bypass_10_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_0_data_26 <= io_in_c_bypass_11_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_0_is_stationary_26 <= io_in_c_bypass_11_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_1_data_26 <= io_in_c_bypass_11_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_1_is_stationary_26 <= io_in_c_bypass_11_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_2_data_26 <= io_in_c_bypass_11_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_2_is_stationary_26 <= io_in_c_bypass_11_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_3_data_26 <= io_in_c_bypass_11_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_3_is_stationary_26 <= io_in_c_bypass_11_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_0_data_26 <= io_in_c_bypass_12_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_0_is_stationary_26 <= io_in_c_bypass_12_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_1_data_26 <= io_in_c_bypass_12_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_1_is_stationary_26 <= io_in_c_bypass_12_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_2_data_26 <= io_in_c_bypass_12_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_2_is_stationary_26 <= io_in_c_bypass_12_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_3_data_26 <= io_in_c_bypass_12_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_3_is_stationary_26 <= io_in_c_bypass_12_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_0_data_26 <= io_in_c_bypass_13_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_0_is_stationary_26 <= io_in_c_bypass_13_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_1_data_26 <= io_in_c_bypass_13_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_1_is_stationary_26 <= io_in_c_bypass_13_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_2_data_26 <= io_in_c_bypass_13_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_2_is_stationary_26 <= io_in_c_bypass_13_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_3_data_26 <= io_in_c_bypass_13_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_3_is_stationary_26 <= io_in_c_bypass_13_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_0_data_26 <= io_in_c_bypass_14_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_0_is_stationary_26 <= io_in_c_bypass_14_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_1_data_26 <= io_in_c_bypass_14_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_1_is_stationary_26 <= io_in_c_bypass_14_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_2_data_26 <= io_in_c_bypass_14_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_2_is_stationary_26 <= io_in_c_bypass_14_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_3_data_26 <= io_in_c_bypass_14_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_3_is_stationary_26 <= io_in_c_bypass_14_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_0_data_26 <= io_in_c_bypass_15_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_0_is_stationary_26 <= io_in_c_bypass_15_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_1_data_26 <= io_in_c_bypass_15_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_1_is_stationary_26 <= io_in_c_bypass_15_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_2_data_26 <= io_in_c_bypass_15_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_2_is_stationary_26 <= io_in_c_bypass_15_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_3_data_26 <= io_in_c_bypass_15_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_3_is_stationary_26 <= io_in_c_bypass_15_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_0_data_26 <= io_in_c_bypass_16_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_0_is_stationary_26 <= io_in_c_bypass_16_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_1_data_26 <= io_in_c_bypass_16_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_1_is_stationary_26 <= io_in_c_bypass_16_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_2_data_26 <= io_in_c_bypass_16_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_2_is_stationary_26 <= io_in_c_bypass_16_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_3_data_26 <= io_in_c_bypass_16_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_3_is_stationary_26 <= io_in_c_bypass_16_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_0_data_26 <= io_in_c_bypass_17_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_0_is_stationary_26 <= io_in_c_bypass_17_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_1_data_26 <= io_in_c_bypass_17_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_1_is_stationary_26 <= io_in_c_bypass_17_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_2_data_26 <= io_in_c_bypass_17_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_2_is_stationary_26 <= io_in_c_bypass_17_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_3_data_26 <= io_in_c_bypass_17_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_3_is_stationary_26 <= io_in_c_bypass_17_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_0_data_26 <= io_in_c_bypass_18_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_0_is_stationary_26 <= io_in_c_bypass_18_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_1_data_26 <= io_in_c_bypass_18_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_1_is_stationary_26 <= io_in_c_bypass_18_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_2_data_26 <= io_in_c_bypass_18_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_2_is_stationary_26 <= io_in_c_bypass_18_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_3_data_26 <= io_in_c_bypass_18_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_3_is_stationary_26 <= io_in_c_bypass_18_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_0_data_26 <= io_in_c_bypass_19_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_0_is_stationary_26 <= io_in_c_bypass_19_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_1_data_26 <= io_in_c_bypass_19_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_1_is_stationary_26 <= io_in_c_bypass_19_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_2_data_26 <= io_in_c_bypass_19_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_2_is_stationary_26 <= io_in_c_bypass_19_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_3_data_26 <= io_in_c_bypass_19_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_3_is_stationary_26 <= io_in_c_bypass_19_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_0_data_26 <= io_in_c_bypass_20_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_0_is_stationary_26 <= io_in_c_bypass_20_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_1_data_26 <= io_in_c_bypass_20_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_1_is_stationary_26 <= io_in_c_bypass_20_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_2_data_26 <= io_in_c_bypass_20_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_2_is_stationary_26 <= io_in_c_bypass_20_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_3_data_26 <= io_in_c_bypass_20_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_3_is_stationary_26 <= io_in_c_bypass_20_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_0_data_26 <= io_in_c_bypass_21_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_0_is_stationary_26 <= io_in_c_bypass_21_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_1_data_26 <= io_in_c_bypass_21_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_1_is_stationary_26 <= io_in_c_bypass_21_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_2_data_26 <= io_in_c_bypass_21_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_2_is_stationary_26 <= io_in_c_bypass_21_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_3_data_26 <= io_in_c_bypass_21_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_3_is_stationary_26 <= io_in_c_bypass_21_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_0_data_26 <= io_in_c_bypass_22_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_0_is_stationary_26 <= io_in_c_bypass_22_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_1_data_26 <= io_in_c_bypass_22_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_1_is_stationary_26 <= io_in_c_bypass_22_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_2_data_26 <= io_in_c_bypass_22_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_2_is_stationary_26 <= io_in_c_bypass_22_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_3_data_26 <= io_in_c_bypass_22_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_3_is_stationary_26 <= io_in_c_bypass_22_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_0_data_26 <= io_in_c_bypass_23_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_0_is_stationary_26 <= io_in_c_bypass_23_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_1_data_26 <= io_in_c_bypass_23_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_1_is_stationary_26 <= io_in_c_bypass_23_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_2_data_26 <= io_in_c_bypass_23_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_2_is_stationary_26 <= io_in_c_bypass_23_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_3_data_26 <= io_in_c_bypass_23_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_3_is_stationary_26 <= io_in_c_bypass_23_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_0_data_26 <= io_in_c_bypass_24_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_0_is_stationary_26 <= io_in_c_bypass_24_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_1_data_26 <= io_in_c_bypass_24_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_1_is_stationary_26 <= io_in_c_bypass_24_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_2_data_26 <= io_in_c_bypass_24_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_2_is_stationary_26 <= io_in_c_bypass_24_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_3_data_26 <= io_in_c_bypass_24_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_3_is_stationary_26 <= io_in_c_bypass_24_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_0_data_26 <= io_in_c_bypass_25_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_0_is_stationary_26 <= io_in_c_bypass_25_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_1_data_26 <= io_in_c_bypass_25_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_1_is_stationary_26 <= io_in_c_bypass_25_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_2_data_26 <= io_in_c_bypass_25_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_2_is_stationary_26 <= io_in_c_bypass_25_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_3_data_26 <= io_in_c_bypass_25_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_3_is_stationary_26 <= io_in_c_bypass_25_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_0_data_26 <= io_in_c_bypass_26_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_0_is_stationary_26 <= io_in_c_bypass_26_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_1_data_26 <= io_in_c_bypass_26_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_1_is_stationary_26 <= io_in_c_bypass_26_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_2_data_26 <= io_in_c_bypass_26_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_2_is_stationary_26 <= io_in_c_bypass_26_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_3_data_26 <= io_in_c_bypass_26_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_3_is_stationary_26 <= io_in_c_bypass_26_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_0_data_26 <= io_in_c_bypass_27_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_0_is_stationary_26 <= io_in_c_bypass_27_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_1_data_26 <= io_in_c_bypass_27_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_1_is_stationary_26 <= io_in_c_bypass_27_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_2_data_26 <= io_in_c_bypass_27_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_2_is_stationary_26 <= io_in_c_bypass_27_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_3_data_26 <= io_in_c_bypass_27_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_3_is_stationary_26 <= io_in_c_bypass_27_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_0_data_26 <= io_in_c_bypass_28_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_0_is_stationary_26 <= io_in_c_bypass_28_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_1_data_26 <= io_in_c_bypass_28_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_1_is_stationary_26 <= io_in_c_bypass_28_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_2_data_26 <= io_in_c_bypass_28_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_2_is_stationary_26 <= io_in_c_bypass_28_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_3_data_26 <= io_in_c_bypass_28_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_3_is_stationary_26 <= io_in_c_bypass_28_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_0_data_26 <= io_in_c_bypass_29_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_0_is_stationary_26 <= io_in_c_bypass_29_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_1_data_26 <= io_in_c_bypass_29_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_1_is_stationary_26 <= io_in_c_bypass_29_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_2_data_26 <= io_in_c_bypass_29_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_2_is_stationary_26 <= io_in_c_bypass_29_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_3_data_26 <= io_in_c_bypass_29_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_3_is_stationary_26 <= io_in_c_bypass_29_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_0_data_26 <= io_in_c_bypass_30_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_0_is_stationary_26 <= io_in_c_bypass_30_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_1_data_26 <= io_in_c_bypass_30_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_1_is_stationary_26 <= io_in_c_bypass_30_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_2_data_26 <= io_in_c_bypass_30_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_2_is_stationary_26 <= io_in_c_bypass_30_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_3_data_26 <= io_in_c_bypass_30_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_3_is_stationary_26 <= io_in_c_bypass_30_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_0_data_26 <= io_in_c_bypass_31_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_0_is_stationary_26 <= io_in_c_bypass_31_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_1_data_26 <= io_in_c_bypass_31_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_1_is_stationary_26 <= io_in_c_bypass_31_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_2_data_26 <= io_in_c_bypass_31_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_2_is_stationary_26 <= io_in_c_bypass_31_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_3_data_26 <= io_in_c_bypass_31_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_3_is_stationary_26 <= io_in_c_bypass_31_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_0_data_27 <= io_in_c_bypass_0_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_0_is_stationary_27 <= io_in_c_bypass_0_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_1_data_27 <= io_in_c_bypass_0_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_1_is_stationary_27 <= io_in_c_bypass_0_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_2_data_27 <= io_in_c_bypass_0_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_2_is_stationary_27 <= io_in_c_bypass_0_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_3_data_27 <= io_in_c_bypass_0_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_3_is_stationary_27 <= io_in_c_bypass_0_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_0_data_27 <= io_in_c_bypass_1_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_0_is_stationary_27 <= io_in_c_bypass_1_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_1_data_27 <= io_in_c_bypass_1_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_1_is_stationary_27 <= io_in_c_bypass_1_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_2_data_27 <= io_in_c_bypass_1_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_2_is_stationary_27 <= io_in_c_bypass_1_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_3_data_27 <= io_in_c_bypass_1_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_3_is_stationary_27 <= io_in_c_bypass_1_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_0_data_27 <= io_in_c_bypass_2_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_0_is_stationary_27 <= io_in_c_bypass_2_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_1_data_27 <= io_in_c_bypass_2_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_1_is_stationary_27 <= io_in_c_bypass_2_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_2_data_27 <= io_in_c_bypass_2_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_2_is_stationary_27 <= io_in_c_bypass_2_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_3_data_27 <= io_in_c_bypass_2_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_3_is_stationary_27 <= io_in_c_bypass_2_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_0_data_27 <= io_in_c_bypass_3_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_0_is_stationary_27 <= io_in_c_bypass_3_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_1_data_27 <= io_in_c_bypass_3_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_1_is_stationary_27 <= io_in_c_bypass_3_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_2_data_27 <= io_in_c_bypass_3_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_2_is_stationary_27 <= io_in_c_bypass_3_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_3_data_27 <= io_in_c_bypass_3_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_3_is_stationary_27 <= io_in_c_bypass_3_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_0_data_27 <= io_in_c_bypass_4_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_0_is_stationary_27 <= io_in_c_bypass_4_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_1_data_27 <= io_in_c_bypass_4_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_1_is_stationary_27 <= io_in_c_bypass_4_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_2_data_27 <= io_in_c_bypass_4_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_2_is_stationary_27 <= io_in_c_bypass_4_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_3_data_27 <= io_in_c_bypass_4_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_3_is_stationary_27 <= io_in_c_bypass_4_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_0_data_27 <= io_in_c_bypass_5_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_0_is_stationary_27 <= io_in_c_bypass_5_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_1_data_27 <= io_in_c_bypass_5_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_1_is_stationary_27 <= io_in_c_bypass_5_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_2_data_27 <= io_in_c_bypass_5_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_2_is_stationary_27 <= io_in_c_bypass_5_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_3_data_27 <= io_in_c_bypass_5_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_3_is_stationary_27 <= io_in_c_bypass_5_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_0_data_27 <= io_in_c_bypass_6_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_0_is_stationary_27 <= io_in_c_bypass_6_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_1_data_27 <= io_in_c_bypass_6_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_1_is_stationary_27 <= io_in_c_bypass_6_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_2_data_27 <= io_in_c_bypass_6_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_2_is_stationary_27 <= io_in_c_bypass_6_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_3_data_27 <= io_in_c_bypass_6_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_3_is_stationary_27 <= io_in_c_bypass_6_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_0_data_27 <= io_in_c_bypass_7_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_0_is_stationary_27 <= io_in_c_bypass_7_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_1_data_27 <= io_in_c_bypass_7_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_1_is_stationary_27 <= io_in_c_bypass_7_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_2_data_27 <= io_in_c_bypass_7_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_2_is_stationary_27 <= io_in_c_bypass_7_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_3_data_27 <= io_in_c_bypass_7_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_3_is_stationary_27 <= io_in_c_bypass_7_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_0_data_27 <= io_in_c_bypass_8_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_0_is_stationary_27 <= io_in_c_bypass_8_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_1_data_27 <= io_in_c_bypass_8_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_1_is_stationary_27 <= io_in_c_bypass_8_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_2_data_27 <= io_in_c_bypass_8_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_2_is_stationary_27 <= io_in_c_bypass_8_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_3_data_27 <= io_in_c_bypass_8_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_3_is_stationary_27 <= io_in_c_bypass_8_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_0_data_27 <= io_in_c_bypass_9_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_0_is_stationary_27 <= io_in_c_bypass_9_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_1_data_27 <= io_in_c_bypass_9_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_1_is_stationary_27 <= io_in_c_bypass_9_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_2_data_27 <= io_in_c_bypass_9_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_2_is_stationary_27 <= io_in_c_bypass_9_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_3_data_27 <= io_in_c_bypass_9_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_3_is_stationary_27 <= io_in_c_bypass_9_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_0_data_27 <= io_in_c_bypass_10_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_0_is_stationary_27 <= io_in_c_bypass_10_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_1_data_27 <= io_in_c_bypass_10_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_1_is_stationary_27 <= io_in_c_bypass_10_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_2_data_27 <= io_in_c_bypass_10_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_2_is_stationary_27 <= io_in_c_bypass_10_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_3_data_27 <= io_in_c_bypass_10_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_3_is_stationary_27 <= io_in_c_bypass_10_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_0_data_27 <= io_in_c_bypass_11_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_0_is_stationary_27 <= io_in_c_bypass_11_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_1_data_27 <= io_in_c_bypass_11_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_1_is_stationary_27 <= io_in_c_bypass_11_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_2_data_27 <= io_in_c_bypass_11_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_2_is_stationary_27 <= io_in_c_bypass_11_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_3_data_27 <= io_in_c_bypass_11_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_3_is_stationary_27 <= io_in_c_bypass_11_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_0_data_27 <= io_in_c_bypass_12_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_0_is_stationary_27 <= io_in_c_bypass_12_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_1_data_27 <= io_in_c_bypass_12_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_1_is_stationary_27 <= io_in_c_bypass_12_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_2_data_27 <= io_in_c_bypass_12_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_2_is_stationary_27 <= io_in_c_bypass_12_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_3_data_27 <= io_in_c_bypass_12_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_3_is_stationary_27 <= io_in_c_bypass_12_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_0_data_27 <= io_in_c_bypass_13_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_0_is_stationary_27 <= io_in_c_bypass_13_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_1_data_27 <= io_in_c_bypass_13_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_1_is_stationary_27 <= io_in_c_bypass_13_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_2_data_27 <= io_in_c_bypass_13_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_2_is_stationary_27 <= io_in_c_bypass_13_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_3_data_27 <= io_in_c_bypass_13_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_3_is_stationary_27 <= io_in_c_bypass_13_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_0_data_27 <= io_in_c_bypass_14_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_0_is_stationary_27 <= io_in_c_bypass_14_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_1_data_27 <= io_in_c_bypass_14_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_1_is_stationary_27 <= io_in_c_bypass_14_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_2_data_27 <= io_in_c_bypass_14_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_2_is_stationary_27 <= io_in_c_bypass_14_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_3_data_27 <= io_in_c_bypass_14_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_3_is_stationary_27 <= io_in_c_bypass_14_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_0_data_27 <= io_in_c_bypass_15_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_0_is_stationary_27 <= io_in_c_bypass_15_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_1_data_27 <= io_in_c_bypass_15_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_1_is_stationary_27 <= io_in_c_bypass_15_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_2_data_27 <= io_in_c_bypass_15_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_2_is_stationary_27 <= io_in_c_bypass_15_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_3_data_27 <= io_in_c_bypass_15_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_3_is_stationary_27 <= io_in_c_bypass_15_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_0_data_27 <= io_in_c_bypass_16_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_0_is_stationary_27 <= io_in_c_bypass_16_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_1_data_27 <= io_in_c_bypass_16_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_1_is_stationary_27 <= io_in_c_bypass_16_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_2_data_27 <= io_in_c_bypass_16_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_2_is_stationary_27 <= io_in_c_bypass_16_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_3_data_27 <= io_in_c_bypass_16_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_3_is_stationary_27 <= io_in_c_bypass_16_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_0_data_27 <= io_in_c_bypass_17_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_0_is_stationary_27 <= io_in_c_bypass_17_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_1_data_27 <= io_in_c_bypass_17_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_1_is_stationary_27 <= io_in_c_bypass_17_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_2_data_27 <= io_in_c_bypass_17_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_2_is_stationary_27 <= io_in_c_bypass_17_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_3_data_27 <= io_in_c_bypass_17_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_3_is_stationary_27 <= io_in_c_bypass_17_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_0_data_27 <= io_in_c_bypass_18_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_0_is_stationary_27 <= io_in_c_bypass_18_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_1_data_27 <= io_in_c_bypass_18_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_1_is_stationary_27 <= io_in_c_bypass_18_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_2_data_27 <= io_in_c_bypass_18_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_2_is_stationary_27 <= io_in_c_bypass_18_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_3_data_27 <= io_in_c_bypass_18_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_3_is_stationary_27 <= io_in_c_bypass_18_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_0_data_27 <= io_in_c_bypass_19_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_0_is_stationary_27 <= io_in_c_bypass_19_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_1_data_27 <= io_in_c_bypass_19_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_1_is_stationary_27 <= io_in_c_bypass_19_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_2_data_27 <= io_in_c_bypass_19_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_2_is_stationary_27 <= io_in_c_bypass_19_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_3_data_27 <= io_in_c_bypass_19_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_3_is_stationary_27 <= io_in_c_bypass_19_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_0_data_27 <= io_in_c_bypass_20_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_0_is_stationary_27 <= io_in_c_bypass_20_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_1_data_27 <= io_in_c_bypass_20_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_1_is_stationary_27 <= io_in_c_bypass_20_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_2_data_27 <= io_in_c_bypass_20_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_2_is_stationary_27 <= io_in_c_bypass_20_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_3_data_27 <= io_in_c_bypass_20_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_3_is_stationary_27 <= io_in_c_bypass_20_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_0_data_27 <= io_in_c_bypass_21_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_0_is_stationary_27 <= io_in_c_bypass_21_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_1_data_27 <= io_in_c_bypass_21_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_1_is_stationary_27 <= io_in_c_bypass_21_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_2_data_27 <= io_in_c_bypass_21_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_2_is_stationary_27 <= io_in_c_bypass_21_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_3_data_27 <= io_in_c_bypass_21_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_3_is_stationary_27 <= io_in_c_bypass_21_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_0_data_27 <= io_in_c_bypass_22_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_0_is_stationary_27 <= io_in_c_bypass_22_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_1_data_27 <= io_in_c_bypass_22_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_1_is_stationary_27 <= io_in_c_bypass_22_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_2_data_27 <= io_in_c_bypass_22_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_2_is_stationary_27 <= io_in_c_bypass_22_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_3_data_27 <= io_in_c_bypass_22_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_3_is_stationary_27 <= io_in_c_bypass_22_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_0_data_27 <= io_in_c_bypass_23_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_0_is_stationary_27 <= io_in_c_bypass_23_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_1_data_27 <= io_in_c_bypass_23_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_1_is_stationary_27 <= io_in_c_bypass_23_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_2_data_27 <= io_in_c_bypass_23_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_2_is_stationary_27 <= io_in_c_bypass_23_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_3_data_27 <= io_in_c_bypass_23_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_3_is_stationary_27 <= io_in_c_bypass_23_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_0_data_27 <= io_in_c_bypass_24_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_0_is_stationary_27 <= io_in_c_bypass_24_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_1_data_27 <= io_in_c_bypass_24_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_1_is_stationary_27 <= io_in_c_bypass_24_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_2_data_27 <= io_in_c_bypass_24_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_2_is_stationary_27 <= io_in_c_bypass_24_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_3_data_27 <= io_in_c_bypass_24_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_3_is_stationary_27 <= io_in_c_bypass_24_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_0_data_27 <= io_in_c_bypass_25_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_0_is_stationary_27 <= io_in_c_bypass_25_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_1_data_27 <= io_in_c_bypass_25_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_1_is_stationary_27 <= io_in_c_bypass_25_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_2_data_27 <= io_in_c_bypass_25_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_2_is_stationary_27 <= io_in_c_bypass_25_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_3_data_27 <= io_in_c_bypass_25_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_3_is_stationary_27 <= io_in_c_bypass_25_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_0_data_27 <= io_in_c_bypass_26_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_0_is_stationary_27 <= io_in_c_bypass_26_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_1_data_27 <= io_in_c_bypass_26_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_1_is_stationary_27 <= io_in_c_bypass_26_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_2_data_27 <= io_in_c_bypass_26_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_2_is_stationary_27 <= io_in_c_bypass_26_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_3_data_27 <= io_in_c_bypass_26_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_3_is_stationary_27 <= io_in_c_bypass_26_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_0_data_27 <= io_in_c_bypass_27_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_0_is_stationary_27 <= io_in_c_bypass_27_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_1_data_27 <= io_in_c_bypass_27_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_1_is_stationary_27 <= io_in_c_bypass_27_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_2_data_27 <= io_in_c_bypass_27_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_2_is_stationary_27 <= io_in_c_bypass_27_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_3_data_27 <= io_in_c_bypass_27_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_3_is_stationary_27 <= io_in_c_bypass_27_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_0_data_27 <= io_in_c_bypass_28_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_0_is_stationary_27 <= io_in_c_bypass_28_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_1_data_27 <= io_in_c_bypass_28_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_1_is_stationary_27 <= io_in_c_bypass_28_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_2_data_27 <= io_in_c_bypass_28_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_2_is_stationary_27 <= io_in_c_bypass_28_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_3_data_27 <= io_in_c_bypass_28_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_3_is_stationary_27 <= io_in_c_bypass_28_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_0_data_27 <= io_in_c_bypass_29_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_0_is_stationary_27 <= io_in_c_bypass_29_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_1_data_27 <= io_in_c_bypass_29_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_1_is_stationary_27 <= io_in_c_bypass_29_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_2_data_27 <= io_in_c_bypass_29_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_2_is_stationary_27 <= io_in_c_bypass_29_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_3_data_27 <= io_in_c_bypass_29_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_3_is_stationary_27 <= io_in_c_bypass_29_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_0_data_27 <= io_in_c_bypass_30_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_0_is_stationary_27 <= io_in_c_bypass_30_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_1_data_27 <= io_in_c_bypass_30_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_1_is_stationary_27 <= io_in_c_bypass_30_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_2_data_27 <= io_in_c_bypass_30_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_2_is_stationary_27 <= io_in_c_bypass_30_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_3_data_27 <= io_in_c_bypass_30_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_3_is_stationary_27 <= io_in_c_bypass_30_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_0_data_27 <= io_in_c_bypass_31_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_0_is_stationary_27 <= io_in_c_bypass_31_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_1_data_27 <= io_in_c_bypass_31_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_1_is_stationary_27 <= io_in_c_bypass_31_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_2_data_27 <= io_in_c_bypass_31_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_2_is_stationary_27 <= io_in_c_bypass_31_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_3_data_27 <= io_in_c_bypass_31_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_3_is_stationary_27 <= io_in_c_bypass_31_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_0_data_28 <= io_in_c_bypass_0_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_0_is_stationary_28 <= io_in_c_bypass_0_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_1_data_28 <= io_in_c_bypass_0_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_1_is_stationary_28 <= io_in_c_bypass_0_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_2_data_28 <= io_in_c_bypass_0_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_2_is_stationary_28 <= io_in_c_bypass_0_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_3_data_28 <= io_in_c_bypass_0_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_3_is_stationary_28 <= io_in_c_bypass_0_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_0_data_28 <= io_in_c_bypass_1_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_0_is_stationary_28 <= io_in_c_bypass_1_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_1_data_28 <= io_in_c_bypass_1_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_1_is_stationary_28 <= io_in_c_bypass_1_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_2_data_28 <= io_in_c_bypass_1_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_2_is_stationary_28 <= io_in_c_bypass_1_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_3_data_28 <= io_in_c_bypass_1_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_3_is_stationary_28 <= io_in_c_bypass_1_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_0_data_28 <= io_in_c_bypass_2_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_0_is_stationary_28 <= io_in_c_bypass_2_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_1_data_28 <= io_in_c_bypass_2_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_1_is_stationary_28 <= io_in_c_bypass_2_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_2_data_28 <= io_in_c_bypass_2_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_2_is_stationary_28 <= io_in_c_bypass_2_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_3_data_28 <= io_in_c_bypass_2_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_3_is_stationary_28 <= io_in_c_bypass_2_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_0_data_28 <= io_in_c_bypass_3_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_0_is_stationary_28 <= io_in_c_bypass_3_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_1_data_28 <= io_in_c_bypass_3_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_1_is_stationary_28 <= io_in_c_bypass_3_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_2_data_28 <= io_in_c_bypass_3_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_2_is_stationary_28 <= io_in_c_bypass_3_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_3_data_28 <= io_in_c_bypass_3_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_3_is_stationary_28 <= io_in_c_bypass_3_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_0_data_28 <= io_in_c_bypass_4_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_0_is_stationary_28 <= io_in_c_bypass_4_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_1_data_28 <= io_in_c_bypass_4_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_1_is_stationary_28 <= io_in_c_bypass_4_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_2_data_28 <= io_in_c_bypass_4_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_2_is_stationary_28 <= io_in_c_bypass_4_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_3_data_28 <= io_in_c_bypass_4_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_3_is_stationary_28 <= io_in_c_bypass_4_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_0_data_28 <= io_in_c_bypass_5_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_0_is_stationary_28 <= io_in_c_bypass_5_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_1_data_28 <= io_in_c_bypass_5_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_1_is_stationary_28 <= io_in_c_bypass_5_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_2_data_28 <= io_in_c_bypass_5_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_2_is_stationary_28 <= io_in_c_bypass_5_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_3_data_28 <= io_in_c_bypass_5_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_3_is_stationary_28 <= io_in_c_bypass_5_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_0_data_28 <= io_in_c_bypass_6_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_0_is_stationary_28 <= io_in_c_bypass_6_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_1_data_28 <= io_in_c_bypass_6_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_1_is_stationary_28 <= io_in_c_bypass_6_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_2_data_28 <= io_in_c_bypass_6_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_2_is_stationary_28 <= io_in_c_bypass_6_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_3_data_28 <= io_in_c_bypass_6_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_3_is_stationary_28 <= io_in_c_bypass_6_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_0_data_28 <= io_in_c_bypass_7_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_0_is_stationary_28 <= io_in_c_bypass_7_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_1_data_28 <= io_in_c_bypass_7_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_1_is_stationary_28 <= io_in_c_bypass_7_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_2_data_28 <= io_in_c_bypass_7_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_2_is_stationary_28 <= io_in_c_bypass_7_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_3_data_28 <= io_in_c_bypass_7_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_3_is_stationary_28 <= io_in_c_bypass_7_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_0_data_28 <= io_in_c_bypass_8_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_0_is_stationary_28 <= io_in_c_bypass_8_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_1_data_28 <= io_in_c_bypass_8_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_1_is_stationary_28 <= io_in_c_bypass_8_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_2_data_28 <= io_in_c_bypass_8_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_2_is_stationary_28 <= io_in_c_bypass_8_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_3_data_28 <= io_in_c_bypass_8_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_3_is_stationary_28 <= io_in_c_bypass_8_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_0_data_28 <= io_in_c_bypass_9_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_0_is_stationary_28 <= io_in_c_bypass_9_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_1_data_28 <= io_in_c_bypass_9_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_1_is_stationary_28 <= io_in_c_bypass_9_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_2_data_28 <= io_in_c_bypass_9_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_2_is_stationary_28 <= io_in_c_bypass_9_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_3_data_28 <= io_in_c_bypass_9_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_3_is_stationary_28 <= io_in_c_bypass_9_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_0_data_28 <= io_in_c_bypass_10_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_0_is_stationary_28 <= io_in_c_bypass_10_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_1_data_28 <= io_in_c_bypass_10_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_1_is_stationary_28 <= io_in_c_bypass_10_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_2_data_28 <= io_in_c_bypass_10_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_2_is_stationary_28 <= io_in_c_bypass_10_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_3_data_28 <= io_in_c_bypass_10_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_3_is_stationary_28 <= io_in_c_bypass_10_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_0_data_28 <= io_in_c_bypass_11_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_0_is_stationary_28 <= io_in_c_bypass_11_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_1_data_28 <= io_in_c_bypass_11_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_1_is_stationary_28 <= io_in_c_bypass_11_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_2_data_28 <= io_in_c_bypass_11_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_2_is_stationary_28 <= io_in_c_bypass_11_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_3_data_28 <= io_in_c_bypass_11_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_3_is_stationary_28 <= io_in_c_bypass_11_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_0_data_28 <= io_in_c_bypass_12_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_0_is_stationary_28 <= io_in_c_bypass_12_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_1_data_28 <= io_in_c_bypass_12_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_1_is_stationary_28 <= io_in_c_bypass_12_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_2_data_28 <= io_in_c_bypass_12_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_2_is_stationary_28 <= io_in_c_bypass_12_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_3_data_28 <= io_in_c_bypass_12_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_3_is_stationary_28 <= io_in_c_bypass_12_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_0_data_28 <= io_in_c_bypass_13_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_0_is_stationary_28 <= io_in_c_bypass_13_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_1_data_28 <= io_in_c_bypass_13_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_1_is_stationary_28 <= io_in_c_bypass_13_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_2_data_28 <= io_in_c_bypass_13_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_2_is_stationary_28 <= io_in_c_bypass_13_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_3_data_28 <= io_in_c_bypass_13_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_3_is_stationary_28 <= io_in_c_bypass_13_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_0_data_28 <= io_in_c_bypass_14_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_0_is_stationary_28 <= io_in_c_bypass_14_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_1_data_28 <= io_in_c_bypass_14_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_1_is_stationary_28 <= io_in_c_bypass_14_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_2_data_28 <= io_in_c_bypass_14_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_2_is_stationary_28 <= io_in_c_bypass_14_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_3_data_28 <= io_in_c_bypass_14_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_3_is_stationary_28 <= io_in_c_bypass_14_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_0_data_28 <= io_in_c_bypass_15_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_0_is_stationary_28 <= io_in_c_bypass_15_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_1_data_28 <= io_in_c_bypass_15_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_1_is_stationary_28 <= io_in_c_bypass_15_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_2_data_28 <= io_in_c_bypass_15_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_2_is_stationary_28 <= io_in_c_bypass_15_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_3_data_28 <= io_in_c_bypass_15_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_3_is_stationary_28 <= io_in_c_bypass_15_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_0_data_28 <= io_in_c_bypass_16_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_0_is_stationary_28 <= io_in_c_bypass_16_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_1_data_28 <= io_in_c_bypass_16_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_1_is_stationary_28 <= io_in_c_bypass_16_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_2_data_28 <= io_in_c_bypass_16_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_2_is_stationary_28 <= io_in_c_bypass_16_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_3_data_28 <= io_in_c_bypass_16_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_3_is_stationary_28 <= io_in_c_bypass_16_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_0_data_28 <= io_in_c_bypass_17_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_0_is_stationary_28 <= io_in_c_bypass_17_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_1_data_28 <= io_in_c_bypass_17_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_1_is_stationary_28 <= io_in_c_bypass_17_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_2_data_28 <= io_in_c_bypass_17_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_2_is_stationary_28 <= io_in_c_bypass_17_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_3_data_28 <= io_in_c_bypass_17_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_3_is_stationary_28 <= io_in_c_bypass_17_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_0_data_28 <= io_in_c_bypass_18_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_0_is_stationary_28 <= io_in_c_bypass_18_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_1_data_28 <= io_in_c_bypass_18_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_1_is_stationary_28 <= io_in_c_bypass_18_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_2_data_28 <= io_in_c_bypass_18_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_2_is_stationary_28 <= io_in_c_bypass_18_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_3_data_28 <= io_in_c_bypass_18_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_3_is_stationary_28 <= io_in_c_bypass_18_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_0_data_28 <= io_in_c_bypass_19_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_0_is_stationary_28 <= io_in_c_bypass_19_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_1_data_28 <= io_in_c_bypass_19_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_1_is_stationary_28 <= io_in_c_bypass_19_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_2_data_28 <= io_in_c_bypass_19_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_2_is_stationary_28 <= io_in_c_bypass_19_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_3_data_28 <= io_in_c_bypass_19_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_3_is_stationary_28 <= io_in_c_bypass_19_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_0_data_28 <= io_in_c_bypass_20_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_0_is_stationary_28 <= io_in_c_bypass_20_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_1_data_28 <= io_in_c_bypass_20_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_1_is_stationary_28 <= io_in_c_bypass_20_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_2_data_28 <= io_in_c_bypass_20_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_2_is_stationary_28 <= io_in_c_bypass_20_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_3_data_28 <= io_in_c_bypass_20_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_3_is_stationary_28 <= io_in_c_bypass_20_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_0_data_28 <= io_in_c_bypass_21_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_0_is_stationary_28 <= io_in_c_bypass_21_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_1_data_28 <= io_in_c_bypass_21_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_1_is_stationary_28 <= io_in_c_bypass_21_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_2_data_28 <= io_in_c_bypass_21_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_2_is_stationary_28 <= io_in_c_bypass_21_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_3_data_28 <= io_in_c_bypass_21_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_3_is_stationary_28 <= io_in_c_bypass_21_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_0_data_28 <= io_in_c_bypass_22_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_0_is_stationary_28 <= io_in_c_bypass_22_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_1_data_28 <= io_in_c_bypass_22_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_1_is_stationary_28 <= io_in_c_bypass_22_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_2_data_28 <= io_in_c_bypass_22_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_2_is_stationary_28 <= io_in_c_bypass_22_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_3_data_28 <= io_in_c_bypass_22_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_3_is_stationary_28 <= io_in_c_bypass_22_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_0_data_28 <= io_in_c_bypass_23_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_0_is_stationary_28 <= io_in_c_bypass_23_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_1_data_28 <= io_in_c_bypass_23_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_1_is_stationary_28 <= io_in_c_bypass_23_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_2_data_28 <= io_in_c_bypass_23_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_2_is_stationary_28 <= io_in_c_bypass_23_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_3_data_28 <= io_in_c_bypass_23_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_3_is_stationary_28 <= io_in_c_bypass_23_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_0_data_28 <= io_in_c_bypass_24_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_0_is_stationary_28 <= io_in_c_bypass_24_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_1_data_28 <= io_in_c_bypass_24_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_1_is_stationary_28 <= io_in_c_bypass_24_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_2_data_28 <= io_in_c_bypass_24_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_2_is_stationary_28 <= io_in_c_bypass_24_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_3_data_28 <= io_in_c_bypass_24_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_3_is_stationary_28 <= io_in_c_bypass_24_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_0_data_28 <= io_in_c_bypass_25_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_0_is_stationary_28 <= io_in_c_bypass_25_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_1_data_28 <= io_in_c_bypass_25_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_1_is_stationary_28 <= io_in_c_bypass_25_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_2_data_28 <= io_in_c_bypass_25_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_2_is_stationary_28 <= io_in_c_bypass_25_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_3_data_28 <= io_in_c_bypass_25_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_3_is_stationary_28 <= io_in_c_bypass_25_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_0_data_28 <= io_in_c_bypass_26_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_0_is_stationary_28 <= io_in_c_bypass_26_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_1_data_28 <= io_in_c_bypass_26_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_1_is_stationary_28 <= io_in_c_bypass_26_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_2_data_28 <= io_in_c_bypass_26_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_2_is_stationary_28 <= io_in_c_bypass_26_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_3_data_28 <= io_in_c_bypass_26_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_3_is_stationary_28 <= io_in_c_bypass_26_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_0_data_28 <= io_in_c_bypass_27_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_0_is_stationary_28 <= io_in_c_bypass_27_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_1_data_28 <= io_in_c_bypass_27_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_1_is_stationary_28 <= io_in_c_bypass_27_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_2_data_28 <= io_in_c_bypass_27_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_2_is_stationary_28 <= io_in_c_bypass_27_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_3_data_28 <= io_in_c_bypass_27_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_3_is_stationary_28 <= io_in_c_bypass_27_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_0_data_28 <= io_in_c_bypass_28_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_0_is_stationary_28 <= io_in_c_bypass_28_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_1_data_28 <= io_in_c_bypass_28_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_1_is_stationary_28 <= io_in_c_bypass_28_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_2_data_28 <= io_in_c_bypass_28_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_2_is_stationary_28 <= io_in_c_bypass_28_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_3_data_28 <= io_in_c_bypass_28_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_3_is_stationary_28 <= io_in_c_bypass_28_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_0_data_28 <= io_in_c_bypass_29_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_0_is_stationary_28 <= io_in_c_bypass_29_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_1_data_28 <= io_in_c_bypass_29_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_1_is_stationary_28 <= io_in_c_bypass_29_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_2_data_28 <= io_in_c_bypass_29_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_2_is_stationary_28 <= io_in_c_bypass_29_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_3_data_28 <= io_in_c_bypass_29_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_3_is_stationary_28 <= io_in_c_bypass_29_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_0_data_28 <= io_in_c_bypass_30_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_0_is_stationary_28 <= io_in_c_bypass_30_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_1_data_28 <= io_in_c_bypass_30_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_1_is_stationary_28 <= io_in_c_bypass_30_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_2_data_28 <= io_in_c_bypass_30_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_2_is_stationary_28 <= io_in_c_bypass_30_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_3_data_28 <= io_in_c_bypass_30_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_3_is_stationary_28 <= io_in_c_bypass_30_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_0_data_28 <= io_in_c_bypass_31_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_0_is_stationary_28 <= io_in_c_bypass_31_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_1_data_28 <= io_in_c_bypass_31_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_1_is_stationary_28 <= io_in_c_bypass_31_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_2_data_28 <= io_in_c_bypass_31_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_2_is_stationary_28 <= io_in_c_bypass_31_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_3_data_28 <= io_in_c_bypass_31_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_3_is_stationary_28 <= io_in_c_bypass_31_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_0_data_29 <= io_in_c_bypass_0_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_0_is_stationary_29 <= io_in_c_bypass_0_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_1_data_29 <= io_in_c_bypass_0_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_1_is_stationary_29 <= io_in_c_bypass_0_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_2_data_29 <= io_in_c_bypass_0_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_2_is_stationary_29 <= io_in_c_bypass_0_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_3_data_29 <= io_in_c_bypass_0_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_3_is_stationary_29 <= io_in_c_bypass_0_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_0_data_29 <= io_in_c_bypass_1_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_0_is_stationary_29 <= io_in_c_bypass_1_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_1_data_29 <= io_in_c_bypass_1_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_1_is_stationary_29 <= io_in_c_bypass_1_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_2_data_29 <= io_in_c_bypass_1_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_2_is_stationary_29 <= io_in_c_bypass_1_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_3_data_29 <= io_in_c_bypass_1_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_3_is_stationary_29 <= io_in_c_bypass_1_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_0_data_29 <= io_in_c_bypass_2_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_0_is_stationary_29 <= io_in_c_bypass_2_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_1_data_29 <= io_in_c_bypass_2_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_1_is_stationary_29 <= io_in_c_bypass_2_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_2_data_29 <= io_in_c_bypass_2_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_2_is_stationary_29 <= io_in_c_bypass_2_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_3_data_29 <= io_in_c_bypass_2_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_3_is_stationary_29 <= io_in_c_bypass_2_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_0_data_29 <= io_in_c_bypass_3_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_0_is_stationary_29 <= io_in_c_bypass_3_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_1_data_29 <= io_in_c_bypass_3_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_1_is_stationary_29 <= io_in_c_bypass_3_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_2_data_29 <= io_in_c_bypass_3_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_2_is_stationary_29 <= io_in_c_bypass_3_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_3_data_29 <= io_in_c_bypass_3_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_3_is_stationary_29 <= io_in_c_bypass_3_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_0_data_29 <= io_in_c_bypass_4_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_0_is_stationary_29 <= io_in_c_bypass_4_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_1_data_29 <= io_in_c_bypass_4_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_1_is_stationary_29 <= io_in_c_bypass_4_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_2_data_29 <= io_in_c_bypass_4_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_2_is_stationary_29 <= io_in_c_bypass_4_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_3_data_29 <= io_in_c_bypass_4_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_3_is_stationary_29 <= io_in_c_bypass_4_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_0_data_29 <= io_in_c_bypass_5_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_0_is_stationary_29 <= io_in_c_bypass_5_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_1_data_29 <= io_in_c_bypass_5_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_1_is_stationary_29 <= io_in_c_bypass_5_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_2_data_29 <= io_in_c_bypass_5_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_2_is_stationary_29 <= io_in_c_bypass_5_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_3_data_29 <= io_in_c_bypass_5_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_3_is_stationary_29 <= io_in_c_bypass_5_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_0_data_29 <= io_in_c_bypass_6_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_0_is_stationary_29 <= io_in_c_bypass_6_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_1_data_29 <= io_in_c_bypass_6_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_1_is_stationary_29 <= io_in_c_bypass_6_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_2_data_29 <= io_in_c_bypass_6_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_2_is_stationary_29 <= io_in_c_bypass_6_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_3_data_29 <= io_in_c_bypass_6_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_3_is_stationary_29 <= io_in_c_bypass_6_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_0_data_29 <= io_in_c_bypass_7_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_0_is_stationary_29 <= io_in_c_bypass_7_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_1_data_29 <= io_in_c_bypass_7_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_1_is_stationary_29 <= io_in_c_bypass_7_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_2_data_29 <= io_in_c_bypass_7_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_2_is_stationary_29 <= io_in_c_bypass_7_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_3_data_29 <= io_in_c_bypass_7_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_3_is_stationary_29 <= io_in_c_bypass_7_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_0_data_29 <= io_in_c_bypass_8_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_0_is_stationary_29 <= io_in_c_bypass_8_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_1_data_29 <= io_in_c_bypass_8_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_1_is_stationary_29 <= io_in_c_bypass_8_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_2_data_29 <= io_in_c_bypass_8_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_2_is_stationary_29 <= io_in_c_bypass_8_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_3_data_29 <= io_in_c_bypass_8_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_3_is_stationary_29 <= io_in_c_bypass_8_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_0_data_29 <= io_in_c_bypass_9_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_0_is_stationary_29 <= io_in_c_bypass_9_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_1_data_29 <= io_in_c_bypass_9_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_1_is_stationary_29 <= io_in_c_bypass_9_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_2_data_29 <= io_in_c_bypass_9_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_2_is_stationary_29 <= io_in_c_bypass_9_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_3_data_29 <= io_in_c_bypass_9_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_3_is_stationary_29 <= io_in_c_bypass_9_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_0_data_29 <= io_in_c_bypass_10_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_0_is_stationary_29 <= io_in_c_bypass_10_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_1_data_29 <= io_in_c_bypass_10_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_1_is_stationary_29 <= io_in_c_bypass_10_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_2_data_29 <= io_in_c_bypass_10_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_2_is_stationary_29 <= io_in_c_bypass_10_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_3_data_29 <= io_in_c_bypass_10_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_3_is_stationary_29 <= io_in_c_bypass_10_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_0_data_29 <= io_in_c_bypass_11_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_0_is_stationary_29 <= io_in_c_bypass_11_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_1_data_29 <= io_in_c_bypass_11_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_1_is_stationary_29 <= io_in_c_bypass_11_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_2_data_29 <= io_in_c_bypass_11_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_2_is_stationary_29 <= io_in_c_bypass_11_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_3_data_29 <= io_in_c_bypass_11_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_3_is_stationary_29 <= io_in_c_bypass_11_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_0_data_29 <= io_in_c_bypass_12_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_0_is_stationary_29 <= io_in_c_bypass_12_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_1_data_29 <= io_in_c_bypass_12_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_1_is_stationary_29 <= io_in_c_bypass_12_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_2_data_29 <= io_in_c_bypass_12_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_2_is_stationary_29 <= io_in_c_bypass_12_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_3_data_29 <= io_in_c_bypass_12_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_3_is_stationary_29 <= io_in_c_bypass_12_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_0_data_29 <= io_in_c_bypass_13_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_0_is_stationary_29 <= io_in_c_bypass_13_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_1_data_29 <= io_in_c_bypass_13_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_1_is_stationary_29 <= io_in_c_bypass_13_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_2_data_29 <= io_in_c_bypass_13_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_2_is_stationary_29 <= io_in_c_bypass_13_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_3_data_29 <= io_in_c_bypass_13_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_3_is_stationary_29 <= io_in_c_bypass_13_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_0_data_29 <= io_in_c_bypass_14_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_0_is_stationary_29 <= io_in_c_bypass_14_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_1_data_29 <= io_in_c_bypass_14_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_1_is_stationary_29 <= io_in_c_bypass_14_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_2_data_29 <= io_in_c_bypass_14_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_2_is_stationary_29 <= io_in_c_bypass_14_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_3_data_29 <= io_in_c_bypass_14_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_3_is_stationary_29 <= io_in_c_bypass_14_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_0_data_29 <= io_in_c_bypass_15_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_0_is_stationary_29 <= io_in_c_bypass_15_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_1_data_29 <= io_in_c_bypass_15_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_1_is_stationary_29 <= io_in_c_bypass_15_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_2_data_29 <= io_in_c_bypass_15_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_2_is_stationary_29 <= io_in_c_bypass_15_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_3_data_29 <= io_in_c_bypass_15_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_3_is_stationary_29 <= io_in_c_bypass_15_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_0_data_29 <= io_in_c_bypass_16_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_0_is_stationary_29 <= io_in_c_bypass_16_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_1_data_29 <= io_in_c_bypass_16_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_1_is_stationary_29 <= io_in_c_bypass_16_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_2_data_29 <= io_in_c_bypass_16_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_2_is_stationary_29 <= io_in_c_bypass_16_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_3_data_29 <= io_in_c_bypass_16_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_3_is_stationary_29 <= io_in_c_bypass_16_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_0_data_29 <= io_in_c_bypass_17_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_0_is_stationary_29 <= io_in_c_bypass_17_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_1_data_29 <= io_in_c_bypass_17_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_1_is_stationary_29 <= io_in_c_bypass_17_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_2_data_29 <= io_in_c_bypass_17_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_2_is_stationary_29 <= io_in_c_bypass_17_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_3_data_29 <= io_in_c_bypass_17_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_3_is_stationary_29 <= io_in_c_bypass_17_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_0_data_29 <= io_in_c_bypass_18_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_0_is_stationary_29 <= io_in_c_bypass_18_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_1_data_29 <= io_in_c_bypass_18_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_1_is_stationary_29 <= io_in_c_bypass_18_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_2_data_29 <= io_in_c_bypass_18_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_2_is_stationary_29 <= io_in_c_bypass_18_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_3_data_29 <= io_in_c_bypass_18_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_3_is_stationary_29 <= io_in_c_bypass_18_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_0_data_29 <= io_in_c_bypass_19_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_0_is_stationary_29 <= io_in_c_bypass_19_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_1_data_29 <= io_in_c_bypass_19_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_1_is_stationary_29 <= io_in_c_bypass_19_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_2_data_29 <= io_in_c_bypass_19_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_2_is_stationary_29 <= io_in_c_bypass_19_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_3_data_29 <= io_in_c_bypass_19_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_3_is_stationary_29 <= io_in_c_bypass_19_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_0_data_29 <= io_in_c_bypass_20_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_0_is_stationary_29 <= io_in_c_bypass_20_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_1_data_29 <= io_in_c_bypass_20_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_1_is_stationary_29 <= io_in_c_bypass_20_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_2_data_29 <= io_in_c_bypass_20_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_2_is_stationary_29 <= io_in_c_bypass_20_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_3_data_29 <= io_in_c_bypass_20_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_3_is_stationary_29 <= io_in_c_bypass_20_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_0_data_29 <= io_in_c_bypass_21_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_0_is_stationary_29 <= io_in_c_bypass_21_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_1_data_29 <= io_in_c_bypass_21_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_1_is_stationary_29 <= io_in_c_bypass_21_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_2_data_29 <= io_in_c_bypass_21_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_2_is_stationary_29 <= io_in_c_bypass_21_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_3_data_29 <= io_in_c_bypass_21_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_3_is_stationary_29 <= io_in_c_bypass_21_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_0_data_29 <= io_in_c_bypass_22_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_0_is_stationary_29 <= io_in_c_bypass_22_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_1_data_29 <= io_in_c_bypass_22_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_1_is_stationary_29 <= io_in_c_bypass_22_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_2_data_29 <= io_in_c_bypass_22_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_2_is_stationary_29 <= io_in_c_bypass_22_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_3_data_29 <= io_in_c_bypass_22_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_3_is_stationary_29 <= io_in_c_bypass_22_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_0_data_29 <= io_in_c_bypass_23_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_0_is_stationary_29 <= io_in_c_bypass_23_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_1_data_29 <= io_in_c_bypass_23_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_1_is_stationary_29 <= io_in_c_bypass_23_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_2_data_29 <= io_in_c_bypass_23_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_2_is_stationary_29 <= io_in_c_bypass_23_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_3_data_29 <= io_in_c_bypass_23_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_3_is_stationary_29 <= io_in_c_bypass_23_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_0_data_29 <= io_in_c_bypass_24_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_0_is_stationary_29 <= io_in_c_bypass_24_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_1_data_29 <= io_in_c_bypass_24_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_1_is_stationary_29 <= io_in_c_bypass_24_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_2_data_29 <= io_in_c_bypass_24_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_2_is_stationary_29 <= io_in_c_bypass_24_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_3_data_29 <= io_in_c_bypass_24_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_3_is_stationary_29 <= io_in_c_bypass_24_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_0_data_29 <= io_in_c_bypass_25_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_0_is_stationary_29 <= io_in_c_bypass_25_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_1_data_29 <= io_in_c_bypass_25_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_1_is_stationary_29 <= io_in_c_bypass_25_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_2_data_29 <= io_in_c_bypass_25_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_2_is_stationary_29 <= io_in_c_bypass_25_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_3_data_29 <= io_in_c_bypass_25_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_3_is_stationary_29 <= io_in_c_bypass_25_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_0_data_29 <= io_in_c_bypass_26_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_0_is_stationary_29 <= io_in_c_bypass_26_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_1_data_29 <= io_in_c_bypass_26_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_1_is_stationary_29 <= io_in_c_bypass_26_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_2_data_29 <= io_in_c_bypass_26_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_2_is_stationary_29 <= io_in_c_bypass_26_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_3_data_29 <= io_in_c_bypass_26_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_3_is_stationary_29 <= io_in_c_bypass_26_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_0_data_29 <= io_in_c_bypass_27_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_0_is_stationary_29 <= io_in_c_bypass_27_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_1_data_29 <= io_in_c_bypass_27_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_1_is_stationary_29 <= io_in_c_bypass_27_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_2_data_29 <= io_in_c_bypass_27_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_2_is_stationary_29 <= io_in_c_bypass_27_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_3_data_29 <= io_in_c_bypass_27_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_3_is_stationary_29 <= io_in_c_bypass_27_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_0_data_29 <= io_in_c_bypass_28_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_0_is_stationary_29 <= io_in_c_bypass_28_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_1_data_29 <= io_in_c_bypass_28_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_1_is_stationary_29 <= io_in_c_bypass_28_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_2_data_29 <= io_in_c_bypass_28_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_2_is_stationary_29 <= io_in_c_bypass_28_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_3_data_29 <= io_in_c_bypass_28_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_3_is_stationary_29 <= io_in_c_bypass_28_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_0_data_29 <= io_in_c_bypass_29_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_0_is_stationary_29 <= io_in_c_bypass_29_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_1_data_29 <= io_in_c_bypass_29_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_1_is_stationary_29 <= io_in_c_bypass_29_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_2_data_29 <= io_in_c_bypass_29_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_2_is_stationary_29 <= io_in_c_bypass_29_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_3_data_29 <= io_in_c_bypass_29_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_3_is_stationary_29 <= io_in_c_bypass_29_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_0_data_29 <= io_in_c_bypass_30_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_0_is_stationary_29 <= io_in_c_bypass_30_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_1_data_29 <= io_in_c_bypass_30_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_1_is_stationary_29 <= io_in_c_bypass_30_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_2_data_29 <= io_in_c_bypass_30_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_2_is_stationary_29 <= io_in_c_bypass_30_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_3_data_29 <= io_in_c_bypass_30_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_3_is_stationary_29 <= io_in_c_bypass_30_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_0_data_29 <= io_in_c_bypass_31_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_0_is_stationary_29 <= io_in_c_bypass_31_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_1_data_29 <= io_in_c_bypass_31_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_1_is_stationary_29 <= io_in_c_bypass_31_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_2_data_29 <= io_in_c_bypass_31_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_2_is_stationary_29 <= io_in_c_bypass_31_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_3_data_29 <= io_in_c_bypass_31_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_3_is_stationary_29 <= io_in_c_bypass_31_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_0_data_30 <= io_in_c_bypass_0_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_0_is_stationary_30 <= io_in_c_bypass_0_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_1_data_30 <= io_in_c_bypass_0_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_1_is_stationary_30 <= io_in_c_bypass_0_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_2_data_30 <= io_in_c_bypass_0_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_2_is_stationary_30 <= io_in_c_bypass_0_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_3_data_30 <= io_in_c_bypass_0_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_3_is_stationary_30 <= io_in_c_bypass_0_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_0_data_30 <= io_in_c_bypass_1_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_0_is_stationary_30 <= io_in_c_bypass_1_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_1_data_30 <= io_in_c_bypass_1_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_1_is_stationary_30 <= io_in_c_bypass_1_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_2_data_30 <= io_in_c_bypass_1_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_2_is_stationary_30 <= io_in_c_bypass_1_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_3_data_30 <= io_in_c_bypass_1_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_3_is_stationary_30 <= io_in_c_bypass_1_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_0_data_30 <= io_in_c_bypass_2_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_0_is_stationary_30 <= io_in_c_bypass_2_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_1_data_30 <= io_in_c_bypass_2_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_1_is_stationary_30 <= io_in_c_bypass_2_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_2_data_30 <= io_in_c_bypass_2_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_2_is_stationary_30 <= io_in_c_bypass_2_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_3_data_30 <= io_in_c_bypass_2_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_2_3_is_stationary_30 <= io_in_c_bypass_2_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_0_data_30 <= io_in_c_bypass_3_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_0_is_stationary_30 <= io_in_c_bypass_3_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_1_data_30 <= io_in_c_bypass_3_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_1_is_stationary_30 <= io_in_c_bypass_3_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_2_data_30 <= io_in_c_bypass_3_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_2_is_stationary_30 <= io_in_c_bypass_3_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_3_data_30 <= io_in_c_bypass_3_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_3_3_is_stationary_30 <= io_in_c_bypass_3_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_0_data_30 <= io_in_c_bypass_4_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_0_is_stationary_30 <= io_in_c_bypass_4_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_1_data_30 <= io_in_c_bypass_4_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_1_is_stationary_30 <= io_in_c_bypass_4_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_2_data_30 <= io_in_c_bypass_4_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_2_is_stationary_30 <= io_in_c_bypass_4_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_3_data_30 <= io_in_c_bypass_4_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_4_3_is_stationary_30 <= io_in_c_bypass_4_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_0_data_30 <= io_in_c_bypass_5_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_0_is_stationary_30 <= io_in_c_bypass_5_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_1_data_30 <= io_in_c_bypass_5_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_1_is_stationary_30 <= io_in_c_bypass_5_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_2_data_30 <= io_in_c_bypass_5_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_2_is_stationary_30 <= io_in_c_bypass_5_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_3_data_30 <= io_in_c_bypass_5_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_5_3_is_stationary_30 <= io_in_c_bypass_5_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_0_data_30 <= io_in_c_bypass_6_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_0_is_stationary_30 <= io_in_c_bypass_6_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_1_data_30 <= io_in_c_bypass_6_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_1_is_stationary_30 <= io_in_c_bypass_6_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_2_data_30 <= io_in_c_bypass_6_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_2_is_stationary_30 <= io_in_c_bypass_6_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_3_data_30 <= io_in_c_bypass_6_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_6_3_is_stationary_30 <= io_in_c_bypass_6_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_0_data_30 <= io_in_c_bypass_7_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_0_is_stationary_30 <= io_in_c_bypass_7_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_1_data_30 <= io_in_c_bypass_7_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_1_is_stationary_30 <= io_in_c_bypass_7_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_2_data_30 <= io_in_c_bypass_7_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_2_is_stationary_30 <= io_in_c_bypass_7_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_3_data_30 <= io_in_c_bypass_7_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_7_3_is_stationary_30 <= io_in_c_bypass_7_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_0_data_30 <= io_in_c_bypass_8_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_0_is_stationary_30 <= io_in_c_bypass_8_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_1_data_30 <= io_in_c_bypass_8_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_1_is_stationary_30 <= io_in_c_bypass_8_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_2_data_30 <= io_in_c_bypass_8_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_2_is_stationary_30 <= io_in_c_bypass_8_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_3_data_30 <= io_in_c_bypass_8_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_8_3_is_stationary_30 <= io_in_c_bypass_8_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_0_data_30 <= io_in_c_bypass_9_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_0_is_stationary_30 <= io_in_c_bypass_9_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_1_data_30 <= io_in_c_bypass_9_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_1_is_stationary_30 <= io_in_c_bypass_9_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_2_data_30 <= io_in_c_bypass_9_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_2_is_stationary_30 <= io_in_c_bypass_9_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_3_data_30 <= io_in_c_bypass_9_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_9_3_is_stationary_30 <= io_in_c_bypass_9_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_0_data_30 <= io_in_c_bypass_10_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_0_is_stationary_30 <= io_in_c_bypass_10_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_1_data_30 <= io_in_c_bypass_10_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_1_is_stationary_30 <= io_in_c_bypass_10_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_2_data_30 <= io_in_c_bypass_10_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_2_is_stationary_30 <= io_in_c_bypass_10_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_3_data_30 <= io_in_c_bypass_10_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_10_3_is_stationary_30 <= io_in_c_bypass_10_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_0_data_30 <= io_in_c_bypass_11_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_0_is_stationary_30 <= io_in_c_bypass_11_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_1_data_30 <= io_in_c_bypass_11_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_1_is_stationary_30 <= io_in_c_bypass_11_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_2_data_30 <= io_in_c_bypass_11_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_2_is_stationary_30 <= io_in_c_bypass_11_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_3_data_30 <= io_in_c_bypass_11_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_11_3_is_stationary_30 <= io_in_c_bypass_11_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_0_data_30 <= io_in_c_bypass_12_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_0_is_stationary_30 <= io_in_c_bypass_12_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_1_data_30 <= io_in_c_bypass_12_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_1_is_stationary_30 <= io_in_c_bypass_12_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_2_data_30 <= io_in_c_bypass_12_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_2_is_stationary_30 <= io_in_c_bypass_12_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_3_data_30 <= io_in_c_bypass_12_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_12_3_is_stationary_30 <= io_in_c_bypass_12_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_0_data_30 <= io_in_c_bypass_13_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_0_is_stationary_30 <= io_in_c_bypass_13_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_1_data_30 <= io_in_c_bypass_13_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_1_is_stationary_30 <= io_in_c_bypass_13_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_2_data_30 <= io_in_c_bypass_13_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_2_is_stationary_30 <= io_in_c_bypass_13_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_3_data_30 <= io_in_c_bypass_13_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_13_3_is_stationary_30 <= io_in_c_bypass_13_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_0_data_30 <= io_in_c_bypass_14_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_0_is_stationary_30 <= io_in_c_bypass_14_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_1_data_30 <= io_in_c_bypass_14_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_1_is_stationary_30 <= io_in_c_bypass_14_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_2_data_30 <= io_in_c_bypass_14_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_2_is_stationary_30 <= io_in_c_bypass_14_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_3_data_30 <= io_in_c_bypass_14_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_14_3_is_stationary_30 <= io_in_c_bypass_14_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_0_data_30 <= io_in_c_bypass_15_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_0_is_stationary_30 <= io_in_c_bypass_15_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_1_data_30 <= io_in_c_bypass_15_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_1_is_stationary_30 <= io_in_c_bypass_15_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_2_data_30 <= io_in_c_bypass_15_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_2_is_stationary_30 <= io_in_c_bypass_15_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_3_data_30 <= io_in_c_bypass_15_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_15_3_is_stationary_30 <= io_in_c_bypass_15_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_0_data_30 <= io_in_c_bypass_16_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_0_is_stationary_30 <= io_in_c_bypass_16_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_1_data_30 <= io_in_c_bypass_16_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_1_is_stationary_30 <= io_in_c_bypass_16_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_2_data_30 <= io_in_c_bypass_16_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_2_is_stationary_30 <= io_in_c_bypass_16_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_3_data_30 <= io_in_c_bypass_16_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_16_3_is_stationary_30 <= io_in_c_bypass_16_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_0_data_30 <= io_in_c_bypass_17_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_0_is_stationary_30 <= io_in_c_bypass_17_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_1_data_30 <= io_in_c_bypass_17_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_1_is_stationary_30 <= io_in_c_bypass_17_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_2_data_30 <= io_in_c_bypass_17_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_2_is_stationary_30 <= io_in_c_bypass_17_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_3_data_30 <= io_in_c_bypass_17_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_17_3_is_stationary_30 <= io_in_c_bypass_17_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_0_data_30 <= io_in_c_bypass_18_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_0_is_stationary_30 <= io_in_c_bypass_18_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_1_data_30 <= io_in_c_bypass_18_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_1_is_stationary_30 <= io_in_c_bypass_18_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_2_data_30 <= io_in_c_bypass_18_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_2_is_stationary_30 <= io_in_c_bypass_18_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_3_data_30 <= io_in_c_bypass_18_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_18_3_is_stationary_30 <= io_in_c_bypass_18_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_0_data_30 <= io_in_c_bypass_19_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_0_is_stationary_30 <= io_in_c_bypass_19_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_1_data_30 <= io_in_c_bypass_19_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_1_is_stationary_30 <= io_in_c_bypass_19_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_2_data_30 <= io_in_c_bypass_19_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_2_is_stationary_30 <= io_in_c_bypass_19_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_3_data_30 <= io_in_c_bypass_19_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_19_3_is_stationary_30 <= io_in_c_bypass_19_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_0_data_30 <= io_in_c_bypass_20_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_0_is_stationary_30 <= io_in_c_bypass_20_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_1_data_30 <= io_in_c_bypass_20_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_1_is_stationary_30 <= io_in_c_bypass_20_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_2_data_30 <= io_in_c_bypass_20_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_2_is_stationary_30 <= io_in_c_bypass_20_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_3_data_30 <= io_in_c_bypass_20_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_20_3_is_stationary_30 <= io_in_c_bypass_20_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_0_data_30 <= io_in_c_bypass_21_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_0_is_stationary_30 <= io_in_c_bypass_21_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_1_data_30 <= io_in_c_bypass_21_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_1_is_stationary_30 <= io_in_c_bypass_21_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_2_data_30 <= io_in_c_bypass_21_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_2_is_stationary_30 <= io_in_c_bypass_21_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_3_data_30 <= io_in_c_bypass_21_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_21_3_is_stationary_30 <= io_in_c_bypass_21_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_0_data_30 <= io_in_c_bypass_22_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_0_is_stationary_30 <= io_in_c_bypass_22_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_1_data_30 <= io_in_c_bypass_22_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_1_is_stationary_30 <= io_in_c_bypass_22_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_2_data_30 <= io_in_c_bypass_22_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_2_is_stationary_30 <= io_in_c_bypass_22_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_3_data_30 <= io_in_c_bypass_22_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_22_3_is_stationary_30 <= io_in_c_bypass_22_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_0_data_30 <= io_in_c_bypass_23_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_0_is_stationary_30 <= io_in_c_bypass_23_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_1_data_30 <= io_in_c_bypass_23_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_1_is_stationary_30 <= io_in_c_bypass_23_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_2_data_30 <= io_in_c_bypass_23_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_2_is_stationary_30 <= io_in_c_bypass_23_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_3_data_30 <= io_in_c_bypass_23_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_23_3_is_stationary_30 <= io_in_c_bypass_23_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_0_data_30 <= io_in_c_bypass_24_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_0_is_stationary_30 <= io_in_c_bypass_24_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_1_data_30 <= io_in_c_bypass_24_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_1_is_stationary_30 <= io_in_c_bypass_24_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_2_data_30 <= io_in_c_bypass_24_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_2_is_stationary_30 <= io_in_c_bypass_24_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_3_data_30 <= io_in_c_bypass_24_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_24_3_is_stationary_30 <= io_in_c_bypass_24_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_0_data_30 <= io_in_c_bypass_25_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_0_is_stationary_30 <= io_in_c_bypass_25_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_1_data_30 <= io_in_c_bypass_25_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_1_is_stationary_30 <= io_in_c_bypass_25_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_2_data_30 <= io_in_c_bypass_25_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_2_is_stationary_30 <= io_in_c_bypass_25_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_3_data_30 <= io_in_c_bypass_25_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_25_3_is_stationary_30 <= io_in_c_bypass_25_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_0_data_30 <= io_in_c_bypass_26_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_0_is_stationary_30 <= io_in_c_bypass_26_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_1_data_30 <= io_in_c_bypass_26_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_1_is_stationary_30 <= io_in_c_bypass_26_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_2_data_30 <= io_in_c_bypass_26_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_2_is_stationary_30 <= io_in_c_bypass_26_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_3_data_30 <= io_in_c_bypass_26_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_26_3_is_stationary_30 <= io_in_c_bypass_26_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_0_data_30 <= io_in_c_bypass_27_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_0_is_stationary_30 <= io_in_c_bypass_27_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_1_data_30 <= io_in_c_bypass_27_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_1_is_stationary_30 <= io_in_c_bypass_27_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_2_data_30 <= io_in_c_bypass_27_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_2_is_stationary_30 <= io_in_c_bypass_27_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_3_data_30 <= io_in_c_bypass_27_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_27_3_is_stationary_30 <= io_in_c_bypass_27_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_0_data_30 <= io_in_c_bypass_28_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_0_is_stationary_30 <= io_in_c_bypass_28_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_1_data_30 <= io_in_c_bypass_28_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_1_is_stationary_30 <= io_in_c_bypass_28_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_2_data_30 <= io_in_c_bypass_28_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_2_is_stationary_30 <= io_in_c_bypass_28_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_3_data_30 <= io_in_c_bypass_28_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_28_3_is_stationary_30 <= io_in_c_bypass_28_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_0_data_30 <= io_in_c_bypass_29_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_0_is_stationary_30 <= io_in_c_bypass_29_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_1_data_30 <= io_in_c_bypass_29_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_1_is_stationary_30 <= io_in_c_bypass_29_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_2_data_30 <= io_in_c_bypass_29_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_2_is_stationary_30 <= io_in_c_bypass_29_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_3_data_30 <= io_in_c_bypass_29_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_29_3_is_stationary_30 <= io_in_c_bypass_29_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_0_data_30 <= io_in_c_bypass_30_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_0_is_stationary_30 <= io_in_c_bypass_30_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_1_data_30 <= io_in_c_bypass_30_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_1_is_stationary_30 <= io_in_c_bypass_30_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_2_data_30 <= io_in_c_bypass_30_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_2_is_stationary_30 <= io_in_c_bypass_30_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_3_data_30 <= io_in_c_bypass_30_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_30_3_is_stationary_30 <= io_in_c_bypass_30_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_0_data_30 <= io_in_c_bypass_31_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_0_is_stationary_30 <= io_in_c_bypass_31_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_1_data_30 <= io_in_c_bypass_31_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_1_is_stationary_30 <= io_in_c_bypass_31_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_2_data_30 <= io_in_c_bypass_31_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_2_is_stationary_30 <= io_in_c_bypass_31_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_3_data_30 <= io_in_c_bypass_31_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_31_3_is_stationary_30 <= io_in_c_bypass_31_3_is_stationary; // @[Reg.scala 39:30]
    io_in_r_input_from_bypass_regNext_0 <= io_in_r_input_from_bypass_0; // @[Reg.scala 39:30]
    io_in_r_input_from_bypass_regNext_1 <= io_in_r_input_from_bypass_1; // @[Reg.scala 39:30]
    io_in_r_input_from_bypass_regNext_2 <= io_in_r_input_from_bypass_2; // @[Reg.scala 39:30]
    io_in_r_input_from_bypass_regNext_3 <= io_in_r_input_from_bypass_3; // @[Reg.scala 39:30]
    io_in_r_input_from_bypass_regNext_4 <= io_in_r_input_from_bypass_4; // @[Reg.scala 39:30]
    io_in_r_input_from_bypass_regNext_5 <= io_in_r_input_from_bypass_5; // @[Reg.scala 39:30]
    io_in_r_input_from_bypass_regNext_6 <= io_in_r_input_from_bypass_6; // @[Reg.scala 39:30]
    io_in_r_input_from_bypass_regNext_7 <= io_in_r_input_from_bypass_7; // @[Reg.scala 39:30]
    io_in_r_input_from_bypass_regNext_8 <= io_in_r_input_from_bypass_8; // @[Reg.scala 39:30]
    io_in_r_input_from_bypass_regNext_9 <= io_in_r_input_from_bypass_9; // @[Reg.scala 39:30]
    io_in_r_input_from_bypass_regNext_10 <= io_in_r_input_from_bypass_10; // @[Reg.scala 39:30]
    io_in_r_input_from_bypass_regNext_11 <= io_in_r_input_from_bypass_11; // @[Reg.scala 39:30]
    io_in_r_input_from_bypass_regNext_12 <= io_in_r_input_from_bypass_12; // @[Reg.scala 39:30]
    io_in_r_input_from_bypass_regNext_13 <= io_in_r_input_from_bypass_13; // @[Reg.scala 39:30]
    io_in_r_input_from_bypass_regNext_14 <= io_in_r_input_from_bypass_14; // @[Reg.scala 39:30]
    io_in_r_input_from_bypass_regNext_15 <= io_in_r_input_from_bypass_15; // @[Reg.scala 39:30]
    io_in_r_input_from_bypass_regNext_16 <= io_in_r_input_from_bypass_16; // @[Reg.scala 39:30]
    io_in_r_input_from_bypass_regNext_17 <= io_in_r_input_from_bypass_17; // @[Reg.scala 39:30]
    io_in_r_input_from_bypass_regNext_18 <= io_in_r_input_from_bypass_18; // @[Reg.scala 39:30]
    io_in_r_input_from_bypass_regNext_19 <= io_in_r_input_from_bypass_19; // @[Reg.scala 39:30]
    io_in_r_input_from_bypass_regNext_20 <= io_in_r_input_from_bypass_20; // @[Reg.scala 39:30]
    io_in_r_input_from_bypass_regNext_21 <= io_in_r_input_from_bypass_21; // @[Reg.scala 39:30]
    io_in_r_input_from_bypass_regNext_22 <= io_in_r_input_from_bypass_22; // @[Reg.scala 39:30]
    io_in_r_input_from_bypass_regNext_23 <= io_in_r_input_from_bypass_23; // @[Reg.scala 39:30]
    io_in_r_input_from_bypass_regNext_24 <= io_in_r_input_from_bypass_24; // @[Reg.scala 39:30]
    io_in_r_input_from_bypass_regNext_25 <= io_in_r_input_from_bypass_25; // @[Reg.scala 39:30]
    io_in_r_input_from_bypass_regNext_26 <= io_in_r_input_from_bypass_26; // @[Reg.scala 39:30]
    io_in_r_input_from_bypass_regNext_27 <= io_in_r_input_from_bypass_27; // @[Reg.scala 39:30]
    io_in_r_input_from_bypass_regNext_28 <= io_in_r_input_from_bypass_28; // @[Reg.scala 39:30]
    io_in_r_input_from_bypass_regNext_29 <= io_in_r_input_from_bypass_29; // @[Reg.scala 39:30]
    io_in_r_input_from_bypass_regNext_30 <= io_in_r_input_from_bypass_30; // @[Reg.scala 39:30]
    io_in_r_input_from_bypass_regNext_31 <= io_in_r_input_from_bypass_31; // @[Reg.scala 39:30]
    io_in_c_input_from_bypass_regNext_0 <= io_in_c_input_from_bypass_0; // @[Reg.scala 39:30]
    io_in_c_input_from_bypass_regNext_1 <= io_in_c_input_from_bypass_1; // @[Reg.scala 39:30]
    io_in_c_input_from_bypass_regNext_2 <= io_in_c_input_from_bypass_2; // @[Reg.scala 39:30]
    io_in_c_input_from_bypass_regNext_3 <= io_in_c_input_from_bypass_3; // @[Reg.scala 39:30]
    io_in_c_input_from_bypass_regNext_4 <= io_in_c_input_from_bypass_4; // @[Reg.scala 39:30]
    io_in_c_input_from_bypass_regNext_5 <= io_in_c_input_from_bypass_5; // @[Reg.scala 39:30]
    io_in_c_input_from_bypass_regNext_6 <= io_in_c_input_from_bypass_6; // @[Reg.scala 39:30]
    io_in_c_input_from_bypass_regNext_7 <= io_in_c_input_from_bypass_7; // @[Reg.scala 39:30]
    io_in_c_input_from_bypass_regNext_8 <= io_in_c_input_from_bypass_8; // @[Reg.scala 39:30]
    io_in_c_input_from_bypass_regNext_9 <= io_in_c_input_from_bypass_9; // @[Reg.scala 39:30]
    io_in_c_input_from_bypass_regNext_10 <= io_in_c_input_from_bypass_10; // @[Reg.scala 39:30]
    io_in_c_input_from_bypass_regNext_11 <= io_in_c_input_from_bypass_11; // @[Reg.scala 39:30]
    io_in_c_input_from_bypass_regNext_12 <= io_in_c_input_from_bypass_12; // @[Reg.scala 39:30]
    io_in_c_input_from_bypass_regNext_13 <= io_in_c_input_from_bypass_13; // @[Reg.scala 39:30]
    io_in_c_input_from_bypass_regNext_14 <= io_in_c_input_from_bypass_14; // @[Reg.scala 39:30]
    io_in_c_input_from_bypass_regNext_15 <= io_in_c_input_from_bypass_15; // @[Reg.scala 39:30]
    io_in_c_input_from_bypass_regNext_16 <= io_in_c_input_from_bypass_16; // @[Reg.scala 39:30]
    io_in_c_input_from_bypass_regNext_17 <= io_in_c_input_from_bypass_17; // @[Reg.scala 39:30]
    io_in_c_input_from_bypass_regNext_18 <= io_in_c_input_from_bypass_18; // @[Reg.scala 39:30]
    io_in_c_input_from_bypass_regNext_19 <= io_in_c_input_from_bypass_19; // @[Reg.scala 39:30]
    io_in_c_input_from_bypass_regNext_20 <= io_in_c_input_from_bypass_20; // @[Reg.scala 39:30]
    io_in_c_input_from_bypass_regNext_21 <= io_in_c_input_from_bypass_21; // @[Reg.scala 39:30]
    io_in_c_input_from_bypass_regNext_22 <= io_in_c_input_from_bypass_22; // @[Reg.scala 39:30]
    io_in_c_input_from_bypass_regNext_23 <= io_in_c_input_from_bypass_23; // @[Reg.scala 39:30]
    io_in_c_input_from_bypass_regNext_24 <= io_in_c_input_from_bypass_24; // @[Reg.scala 39:30]
    io_in_c_input_from_bypass_regNext_25 <= io_in_c_input_from_bypass_25; // @[Reg.scala 39:30]
    io_in_c_input_from_bypass_regNext_26 <= io_in_c_input_from_bypass_26; // @[Reg.scala 39:30]
    io_in_c_input_from_bypass_regNext_27 <= io_in_c_input_from_bypass_27; // @[Reg.scala 39:30]
    io_in_c_input_from_bypass_regNext_28 <= io_in_c_input_from_bypass_28; // @[Reg.scala 39:30]
    io_in_c_input_from_bypass_regNext_29 <= io_in_c_input_from_bypass_29; // @[Reg.scala 39:30]
    io_in_c_input_from_bypass_regNext_30 <= io_in_c_input_from_bypass_30; // @[Reg.scala 39:30]
    io_in_c_input_from_bypass_regNext_31 <= io_in_c_input_from_bypass_31; // @[Reg.scala 39:30]
  end


endmodule

//PEWSOS_15 replaced by PEWSOS_15

//PEWSOS_15 replaced by PEWSOS_15

//PEWSOS_15 replaced by PEWSOS_15

//PEWSOS_15 replaced by PEWSOS_15

//PEWSOS_15 replaced by PEWSOS_15

//PEWSOS_15 replaced by PEWSOS_15

//PEWSOS_15 replaced by PEWSOS_15

//PEWSOS_15 replaced by PEWSOS_15

//PEWSOS_15 replaced by PEWSOS_15

//PEWSOS_15 replaced by PEWSOS_15

//PEWSOS_15 replaced by PEWSOS_15

//PEWSOS_15 replaced by PEWSOS_15

//PEWSOS_15 replaced by PEWSOS_15

//PEWSOS_15 replaced by PEWSOS_15

//PEWSOS_15 replaced by PEWSOS_15

module PEWSOS_15 (
  input      [15:0]   io_in_r_data,
  input               io_in_r_load_store,
  input               io_in_r_df_is_ws,
  input               io_in_r_stall,
  output     [15:0]   io_out_r_data,
  output              io_out_r_load_store,
  output              io_out_r_df_is_ws,
  output              io_out_r_stall,
  input      [15:0]   io_in_c_data,
  input               io_in_c_is_stationary,
  output     [15:0]   io_out_c_data,
  output              io_out_c_is_stationary,
  input               clk,
  input               reset
);

  wire       [15:0]   mac_16_io_psum;
  wire       [15:0]   mac_16_io_weight;
  wire       [15:0]   mac_16_io_result;
  wire                not_stall;
  wire       [15:0]   mac_result;
  reg        [15:0]   stationary;
  reg                 stationary_en;
  wire                when_PEWSOS_l68;
  reg        [15:0]   stationary_reg;
  reg                 io_in_r_stall_regNext;
  reg        [15:0]   io_in_r_data_regNextWhen;
  reg                 io_in_r_load_store_regNextWhen;
  reg                 io_in_r_df_is_ws_regNextWhen;
  reg        [15:0]   out_c_data;
  reg                 out_c_is_stationary;
  wire                when_PEWSOS_l87;
  wire                when_PEWSOS_l95;
  reg        [15:0]   out_c_data_regNextWhen;
  reg                 out_c_is_stationary_regNextWhen;

  Mac_15 mac_16 (
    .io_psum            (mac_16_io_psum[15:0]  ), //i
    .io_weight          (mac_16_io_weight[15:0]), //i
    .io_inputActivation (io_in_r_data[15:0]    ), //i
    .io_result          (mac_16_io_result[15:0])  //o
  );
  assign not_stall = (! io_in_r_stall); // @[BaseType.scala 299:24]
  always @(*) begin
    if(io_in_r_df_is_ws) begin
      stationary = io_in_c_data; // @[PEWSOS.scala 57:16]
    end else begin
      if(io_in_c_is_stationary) begin
        stationary = 16'h0; // @[PEWSOS.scala 61:18]
      end else begin
        stationary = mac_result; // @[PEWSOS.scala 64:18]
      end
    end
  end

  always @(*) begin
    if(io_in_r_df_is_ws) begin
      stationary_en = io_in_r_load_store; // @[PEWSOS.scala 58:19]
    end else begin
      if(io_in_c_is_stationary) begin
        stationary_en = io_in_r_load_store; // @[PEWSOS.scala 62:21]
      end else begin
        stationary_en = 1'b1; // @[PEWSOS.scala 65:21]
      end
    end
  end

  assign when_PEWSOS_l68 = (stationary_en && not_stall); // @[BaseType.scala 305:24]
  assign mac_16_io_psum = (io_in_r_df_is_ws ? io_in_c_data : stationary_reg); // @[PEWSOS.scala 72:15]
  assign mac_16_io_weight = (io_in_r_df_is_ws ? stationary_reg : io_in_c_data); // @[PEWSOS.scala 73:17]
  assign mac_result = mac_16_io_result; // @[PEWSOS.scala 75:14]
  assign io_out_r_stall = io_in_r_stall_regNext; // @[PEWSOS.scala 78:18]
  assign io_out_r_data = io_in_r_data_regNextWhen; // @[PEWSOS.scala 79:17]
  assign io_out_r_load_store = io_in_r_load_store_regNextWhen; // @[PEWSOS.scala 80:23]
  assign io_out_r_df_is_ws = io_in_r_df_is_ws_regNextWhen; // @[PEWSOS.scala 81:21]
  assign when_PEWSOS_l87 = (io_in_c_is_stationary && (! io_in_r_load_store)); // @[BaseType.scala 305:24]
  always @(*) begin
    if(io_in_r_df_is_ws) begin
      if(when_PEWSOS_l87) begin
        out_c_data = io_in_c_data; // @[PEWSOS.scala 88:18]
      end else begin
        out_c_data = mac_result; // @[PEWSOS.scala 91:18]
      end
    end else begin
      if(when_PEWSOS_l95) begin
        out_c_data = io_in_c_data; // @[PEWSOS.scala 96:18]
      end else begin
        if(io_in_r_load_store) begin
          out_c_data = stationary_reg; // @[PEWSOS.scala 99:18]
        end else begin
          out_c_data = io_in_c_data; // @[PEWSOS.scala 102:18]
        end
      end
    end
  end

  always @(*) begin
    if(io_in_r_df_is_ws) begin
      if(when_PEWSOS_l87) begin
        out_c_is_stationary = 1'b1; // @[PEWSOS.scala 89:27]
      end else begin
        out_c_is_stationary = 1'b0; // @[PEWSOS.scala 92:27]
      end
    end else begin
      if(when_PEWSOS_l95) begin
        out_c_is_stationary = 1'b1; // @[PEWSOS.scala 97:27]
      end else begin
        if(io_in_r_load_store) begin
          out_c_is_stationary = 1'b1; // @[PEWSOS.scala 100:27]
        end else begin
          out_c_is_stationary = 1'b0; // @[PEWSOS.scala 103:27]
        end
      end
    end
  end

  assign when_PEWSOS_l95 = (io_in_c_is_stationary && (! io_in_r_load_store)); // @[BaseType.scala 305:24]
  assign io_out_c_data = out_c_data_regNextWhen; // @[PEWSOS.scala 106:17]
  assign io_out_c_is_stationary = out_c_is_stationary_regNextWhen; // @[PEWSOS.scala 107:26]
  always @(posedge clk) begin
    if(when_PEWSOS_l68) begin
      stationary_reg <= stationary; // @[PEWSOS.scala 68:35]
    end
    io_in_r_stall_regNext <= io_in_r_stall; // @[Reg.scala 39:30]
    if(not_stall) begin
      io_in_r_data_regNextWhen <= io_in_r_data; // @[PEWSOS.scala 79:31]
    end
    if(not_stall) begin
      io_in_r_load_store_regNextWhen <= io_in_r_load_store; // @[PEWSOS.scala 80:37]
    end
    if(not_stall) begin
      io_in_r_df_is_ws_regNextWhen <= io_in_r_df_is_ws; // @[PEWSOS.scala 81:35]
    end
    if(not_stall) begin
      out_c_data_regNextWhen <= out_c_data; // @[PEWSOS.scala 106:31]
    end
    if(not_stall) begin
      out_c_is_stationary_regNextWhen <= out_c_is_stationary; // @[PEWSOS.scala 107:40]
    end
  end


endmodule

//Mac_15 replaced by Mac_15

//Mac_15 replaced by Mac_15

//Mac_15 replaced by Mac_15

//Mac_15 replaced by Mac_15

//Mac_15 replaced by Mac_15

//Mac_15 replaced by Mac_15

//Mac_15 replaced by Mac_15

//Mac_15 replaced by Mac_15

//Mac_15 replaced by Mac_15

//Mac_15 replaced by Mac_15

//Mac_15 replaced by Mac_15

//Mac_15 replaced by Mac_15

//Mac_15 replaced by Mac_15

//Mac_15 replaced by Mac_15

//Mac_15 replaced by Mac_15

module Mac_15 (
  input      [15:0]   io_psum,
  input      [15:0]   io_weight,
  input      [15:0]   io_inputActivation,
  output     [15:0]   io_result
);

  wire       [31:0]   _zz_io_result;
  wire       [31:0]   _zz_io_result_1;
  wire       [31:0]   _zz_io_result_2;

  assign _zz_io_result = ($signed(_zz_io_result_1) + $signed(_zz_io_result_2));
  assign _zz_io_result_1 = ($signed(io_inputActivation) * $signed(io_weight));
  assign _zz_io_result_2 = {{16{io_psum[15]}}, io_psum};
  assign io_result = _zz_io_result[15:0]; // @[Mac.scala 14:31]

endmodule
