// Generator : SpinalHDL v1.8.0    git head : 4e3563a282582b41f4eaafc503787757251d23ea
// Component : ArrayTPU
// Git hash  : 880d730121882c0a9e393151e88289ab6120d150

`timescale 1ns/1ps

module ArrayTPU (
  input      [15:0]   io_in_r_0_data,
  input               io_in_r_0_stop_weight,
  input               io_in_r_0_stall,
  input      [15:0]   io_in_r_1_data,
  input               io_in_r_1_stop_weight,
  input               io_in_r_1_stall,
  input      [15:0]   io_in_r_2_data,
  input               io_in_r_2_stop_weight,
  input               io_in_r_2_stall,
  input      [15:0]   io_in_r_3_data,
  input               io_in_r_3_stop_weight,
  input               io_in_r_3_stall,
  input      [15:0]   io_in_r_4_data,
  input               io_in_r_4_stop_weight,
  input               io_in_r_4_stall,
  input      [15:0]   io_in_r_5_data,
  input               io_in_r_5_stop_weight,
  input               io_in_r_5_stall,
  input      [15:0]   io_in_r_6_data,
  input               io_in_r_6_stop_weight,
  input               io_in_r_6_stall,
  input      [15:0]   io_in_r_7_data,
  input               io_in_r_7_stop_weight,
  input               io_in_r_7_stall,
  input      [15:0]   io_in_r_8_data,
  input               io_in_r_8_stop_weight,
  input               io_in_r_8_stall,
  input      [15:0]   io_in_r_9_data,
  input               io_in_r_9_stop_weight,
  input               io_in_r_9_stall,
  input      [15:0]   io_in_r_10_data,
  input               io_in_r_10_stop_weight,
  input               io_in_r_10_stall,
  input      [15:0]   io_in_r_11_data,
  input               io_in_r_11_stop_weight,
  input               io_in_r_11_stall,
  input      [15:0]   io_in_r_12_data,
  input               io_in_r_12_stop_weight,
  input               io_in_r_12_stall,
  input      [15:0]   io_in_r_13_data,
  input               io_in_r_13_stop_weight,
  input               io_in_r_13_stall,
  input      [15:0]   io_in_r_14_data,
  input               io_in_r_14_stop_weight,
  input               io_in_r_14_stall,
  input      [15:0]   io_in_r_15_data,
  input               io_in_r_15_stop_weight,
  input               io_in_r_15_stall,
  input      [15:0]   io_in_r_16_data,
  input               io_in_r_16_stop_weight,
  input               io_in_r_16_stall,
  input      [15:0]   io_in_r_17_data,
  input               io_in_r_17_stop_weight,
  input               io_in_r_17_stall,
  input      [15:0]   io_in_r_18_data,
  input               io_in_r_18_stop_weight,
  input               io_in_r_18_stall,
  input      [15:0]   io_in_r_19_data,
  input               io_in_r_19_stop_weight,
  input               io_in_r_19_stall,
  input      [15:0]   io_in_r_20_data,
  input               io_in_r_20_stop_weight,
  input               io_in_r_20_stall,
  input      [15:0]   io_in_r_21_data,
  input               io_in_r_21_stop_weight,
  input               io_in_r_21_stall,
  input      [15:0]   io_in_r_22_data,
  input               io_in_r_22_stop_weight,
  input               io_in_r_22_stall,
  input      [15:0]   io_in_r_23_data,
  input               io_in_r_23_stop_weight,
  input               io_in_r_23_stall,
  input      [15:0]   io_in_r_24_data,
  input               io_in_r_24_stop_weight,
  input               io_in_r_24_stall,
  input      [15:0]   io_in_r_25_data,
  input               io_in_r_25_stop_weight,
  input               io_in_r_25_stall,
  input      [15:0]   io_in_r_26_data,
  input               io_in_r_26_stop_weight,
  input               io_in_r_26_stall,
  input      [15:0]   io_in_r_27_data,
  input               io_in_r_27_stop_weight,
  input               io_in_r_27_stall,
  input      [15:0]   io_in_r_28_data,
  input               io_in_r_28_stop_weight,
  input               io_in_r_28_stall,
  input      [15:0]   io_in_r_29_data,
  input               io_in_r_29_stop_weight,
  input               io_in_r_29_stall,
  input      [15:0]   io_in_r_30_data,
  input               io_in_r_30_stop_weight,
  input               io_in_r_30_stall,
  input      [15:0]   io_in_r_31_data,
  input               io_in_r_31_stop_weight,
  input               io_in_r_31_stall,
  output     [15:0]   io_out_r_0_data,
  output              io_out_r_0_stop_weight,
  output              io_out_r_0_stall,
  output     [15:0]   io_out_r_1_data,
  output              io_out_r_1_stop_weight,
  output              io_out_r_1_stall,
  output     [15:0]   io_out_r_2_data,
  output              io_out_r_2_stop_weight,
  output              io_out_r_2_stall,
  output     [15:0]   io_out_r_3_data,
  output              io_out_r_3_stop_weight,
  output              io_out_r_3_stall,
  output     [15:0]   io_out_r_4_data,
  output              io_out_r_4_stop_weight,
  output              io_out_r_4_stall,
  output     [15:0]   io_out_r_5_data,
  output              io_out_r_5_stop_weight,
  output              io_out_r_5_stall,
  output     [15:0]   io_out_r_6_data,
  output              io_out_r_6_stop_weight,
  output              io_out_r_6_stall,
  output     [15:0]   io_out_r_7_data,
  output              io_out_r_7_stop_weight,
  output              io_out_r_7_stall,
  output     [15:0]   io_out_r_8_data,
  output              io_out_r_8_stop_weight,
  output              io_out_r_8_stall,
  output     [15:0]   io_out_r_9_data,
  output              io_out_r_9_stop_weight,
  output              io_out_r_9_stall,
  output     [15:0]   io_out_r_10_data,
  output              io_out_r_10_stop_weight,
  output              io_out_r_10_stall,
  output     [15:0]   io_out_r_11_data,
  output              io_out_r_11_stop_weight,
  output              io_out_r_11_stall,
  output     [15:0]   io_out_r_12_data,
  output              io_out_r_12_stop_weight,
  output              io_out_r_12_stall,
  output     [15:0]   io_out_r_13_data,
  output              io_out_r_13_stop_weight,
  output              io_out_r_13_stall,
  output     [15:0]   io_out_r_14_data,
  output              io_out_r_14_stop_weight,
  output              io_out_r_14_stall,
  output     [15:0]   io_out_r_15_data,
  output              io_out_r_15_stop_weight,
  output              io_out_r_15_stall,
  output     [15:0]   io_out_r_16_data,
  output              io_out_r_16_stop_weight,
  output              io_out_r_16_stall,
  output     [15:0]   io_out_r_17_data,
  output              io_out_r_17_stop_weight,
  output              io_out_r_17_stall,
  output     [15:0]   io_out_r_18_data,
  output              io_out_r_18_stop_weight,
  output              io_out_r_18_stall,
  output     [15:0]   io_out_r_19_data,
  output              io_out_r_19_stop_weight,
  output              io_out_r_19_stall,
  output     [15:0]   io_out_r_20_data,
  output              io_out_r_20_stop_weight,
  output              io_out_r_20_stall,
  output     [15:0]   io_out_r_21_data,
  output              io_out_r_21_stop_weight,
  output              io_out_r_21_stall,
  output     [15:0]   io_out_r_22_data,
  output              io_out_r_22_stop_weight,
  output              io_out_r_22_stall,
  output     [15:0]   io_out_r_23_data,
  output              io_out_r_23_stop_weight,
  output              io_out_r_23_stall,
  output     [15:0]   io_out_r_24_data,
  output              io_out_r_24_stop_weight,
  output              io_out_r_24_stall,
  output     [15:0]   io_out_r_25_data,
  output              io_out_r_25_stop_weight,
  output              io_out_r_25_stall,
  output     [15:0]   io_out_r_26_data,
  output              io_out_r_26_stop_weight,
  output              io_out_r_26_stall,
  output     [15:0]   io_out_r_27_data,
  output              io_out_r_27_stop_weight,
  output              io_out_r_27_stall,
  output     [15:0]   io_out_r_28_data,
  output              io_out_r_28_stop_weight,
  output              io_out_r_28_stall,
  output     [15:0]   io_out_r_29_data,
  output              io_out_r_29_stop_weight,
  output              io_out_r_29_stall,
  output     [15:0]   io_out_r_30_data,
  output              io_out_r_30_stop_weight,
  output              io_out_r_30_stall,
  output     [15:0]   io_out_r_31_data,
  output              io_out_r_31_stop_weight,
  output              io_out_r_31_stall,
  input      [15:0]   io_in_c_0_data,
  input               io_in_c_0_is_weight,
  input      [15:0]   io_in_c_1_data,
  input               io_in_c_1_is_weight,
  input      [15:0]   io_in_c_2_data,
  input               io_in_c_2_is_weight,
  input      [15:0]   io_in_c_3_data,
  input               io_in_c_3_is_weight,
  input      [15:0]   io_in_c_4_data,
  input               io_in_c_4_is_weight,
  input      [15:0]   io_in_c_5_data,
  input               io_in_c_5_is_weight,
  input      [15:0]   io_in_c_6_data,
  input               io_in_c_6_is_weight,
  input      [15:0]   io_in_c_7_data,
  input               io_in_c_7_is_weight,
  input      [15:0]   io_in_c_8_data,
  input               io_in_c_8_is_weight,
  input      [15:0]   io_in_c_9_data,
  input               io_in_c_9_is_weight,
  input      [15:0]   io_in_c_10_data,
  input               io_in_c_10_is_weight,
  input      [15:0]   io_in_c_11_data,
  input               io_in_c_11_is_weight,
  input      [15:0]   io_in_c_12_data,
  input               io_in_c_12_is_weight,
  input      [15:0]   io_in_c_13_data,
  input               io_in_c_13_is_weight,
  input      [15:0]   io_in_c_14_data,
  input               io_in_c_14_is_weight,
  input      [15:0]   io_in_c_15_data,
  input               io_in_c_15_is_weight,
  input      [15:0]   io_in_c_16_data,
  input               io_in_c_16_is_weight,
  input      [15:0]   io_in_c_17_data,
  input               io_in_c_17_is_weight,
  input      [15:0]   io_in_c_18_data,
  input               io_in_c_18_is_weight,
  input      [15:0]   io_in_c_19_data,
  input               io_in_c_19_is_weight,
  input      [15:0]   io_in_c_20_data,
  input               io_in_c_20_is_weight,
  input      [15:0]   io_in_c_21_data,
  input               io_in_c_21_is_weight,
  input      [15:0]   io_in_c_22_data,
  input               io_in_c_22_is_weight,
  input      [15:0]   io_in_c_23_data,
  input               io_in_c_23_is_weight,
  input      [15:0]   io_in_c_24_data,
  input               io_in_c_24_is_weight,
  input      [15:0]   io_in_c_25_data,
  input               io_in_c_25_is_weight,
  input      [15:0]   io_in_c_26_data,
  input               io_in_c_26_is_weight,
  input      [15:0]   io_in_c_27_data,
  input               io_in_c_27_is_weight,
  input      [15:0]   io_in_c_28_data,
  input               io_in_c_28_is_weight,
  input      [15:0]   io_in_c_29_data,
  input               io_in_c_29_is_weight,
  input      [15:0]   io_in_c_30_data,
  input               io_in_c_30_is_weight,
  input      [15:0]   io_in_c_31_data,
  input               io_in_c_31_is_weight,
  output     [15:0]   io_out_c_0_data,
  output              io_out_c_0_is_weight,
  output     [15:0]   io_out_c_1_data,
  output              io_out_c_1_is_weight,
  output     [15:0]   io_out_c_2_data,
  output              io_out_c_2_is_weight,
  output     [15:0]   io_out_c_3_data,
  output              io_out_c_3_is_weight,
  output     [15:0]   io_out_c_4_data,
  output              io_out_c_4_is_weight,
  output     [15:0]   io_out_c_5_data,
  output              io_out_c_5_is_weight,
  output     [15:0]   io_out_c_6_data,
  output              io_out_c_6_is_weight,
  output     [15:0]   io_out_c_7_data,
  output              io_out_c_7_is_weight,
  output     [15:0]   io_out_c_8_data,
  output              io_out_c_8_is_weight,
  output     [15:0]   io_out_c_9_data,
  output              io_out_c_9_is_weight,
  output     [15:0]   io_out_c_10_data,
  output              io_out_c_10_is_weight,
  output     [15:0]   io_out_c_11_data,
  output              io_out_c_11_is_weight,
  output     [15:0]   io_out_c_12_data,
  output              io_out_c_12_is_weight,
  output     [15:0]   io_out_c_13_data,
  output              io_out_c_13_is_weight,
  output     [15:0]   io_out_c_14_data,
  output              io_out_c_14_is_weight,
  output     [15:0]   io_out_c_15_data,
  output              io_out_c_15_is_weight,
  output     [15:0]   io_out_c_16_data,
  output              io_out_c_16_is_weight,
  output     [15:0]   io_out_c_17_data,
  output              io_out_c_17_is_weight,
  output     [15:0]   io_out_c_18_data,
  output              io_out_c_18_is_weight,
  output     [15:0]   io_out_c_19_data,
  output              io_out_c_19_is_weight,
  output     [15:0]   io_out_c_20_data,
  output              io_out_c_20_is_weight,
  output     [15:0]   io_out_c_21_data,
  output              io_out_c_21_is_weight,
  output     [15:0]   io_out_c_22_data,
  output              io_out_c_22_is_weight,
  output     [15:0]   io_out_c_23_data,
  output              io_out_c_23_is_weight,
  output     [15:0]   io_out_c_24_data,
  output              io_out_c_24_is_weight,
  output     [15:0]   io_out_c_25_data,
  output              io_out_c_25_is_weight,
  output     [15:0]   io_out_c_26_data,
  output              io_out_c_26_is_weight,
  output     [15:0]   io_out_c_27_data,
  output              io_out_c_27_is_weight,
  output     [15:0]   io_out_c_28_data,
  output              io_out_c_28_is_weight,
  output     [15:0]   io_out_c_29_data,
  output              io_out_c_29_is_weight,
  output     [15:0]   io_out_c_30_data,
  output              io_out_c_30_is_weight,
  output     [15:0]   io_out_c_31_data,
  output              io_out_c_31_is_weight,
  input               clk,
  input               reset
);

  wire       [15:0]   pe_mat_0_0_io_out_r_data;
  wire                pe_mat_0_0_io_out_r_stop_weight;
  wire                pe_mat_0_0_io_out_r_stall;
  wire       [15:0]   pe_mat_0_0_io_out_c_data;
  wire                pe_mat_0_0_io_out_c_is_weight;
  wire       [15:0]   pe_mat_0_1_io_out_r_data;
  wire                pe_mat_0_1_io_out_r_stop_weight;
  wire                pe_mat_0_1_io_out_r_stall;
  wire       [15:0]   pe_mat_0_1_io_out_c_data;
  wire                pe_mat_0_1_io_out_c_is_weight;
  wire       [15:0]   pe_mat_0_2_io_out_r_data;
  wire                pe_mat_0_2_io_out_r_stop_weight;
  wire                pe_mat_0_2_io_out_r_stall;
  wire       [15:0]   pe_mat_0_2_io_out_c_data;
  wire                pe_mat_0_2_io_out_c_is_weight;
  wire       [15:0]   pe_mat_0_3_io_out_r_data;
  wire                pe_mat_0_3_io_out_r_stop_weight;
  wire                pe_mat_0_3_io_out_r_stall;
  wire       [15:0]   pe_mat_0_3_io_out_c_data;
  wire                pe_mat_0_3_io_out_c_is_weight;
  wire       [15:0]   pe_mat_0_4_io_out_r_data;
  wire                pe_mat_0_4_io_out_r_stop_weight;
  wire                pe_mat_0_4_io_out_r_stall;
  wire       [15:0]   pe_mat_0_4_io_out_c_data;
  wire                pe_mat_0_4_io_out_c_is_weight;
  wire       [15:0]   pe_mat_0_5_io_out_r_data;
  wire                pe_mat_0_5_io_out_r_stop_weight;
  wire                pe_mat_0_5_io_out_r_stall;
  wire       [15:0]   pe_mat_0_5_io_out_c_data;
  wire                pe_mat_0_5_io_out_c_is_weight;
  wire       [15:0]   pe_mat_0_6_io_out_r_data;
  wire                pe_mat_0_6_io_out_r_stop_weight;
  wire                pe_mat_0_6_io_out_r_stall;
  wire       [15:0]   pe_mat_0_6_io_out_c_data;
  wire                pe_mat_0_6_io_out_c_is_weight;
  wire       [15:0]   pe_mat_0_7_io_out_r_data;
  wire                pe_mat_0_7_io_out_r_stop_weight;
  wire                pe_mat_0_7_io_out_r_stall;
  wire       [15:0]   pe_mat_0_7_io_out_c_data;
  wire                pe_mat_0_7_io_out_c_is_weight;
  wire       [15:0]   pe_mat_0_8_io_out_r_data;
  wire                pe_mat_0_8_io_out_r_stop_weight;
  wire                pe_mat_0_8_io_out_r_stall;
  wire       [15:0]   pe_mat_0_8_io_out_c_data;
  wire                pe_mat_0_8_io_out_c_is_weight;
  wire       [15:0]   pe_mat_0_9_io_out_r_data;
  wire                pe_mat_0_9_io_out_r_stop_weight;
  wire                pe_mat_0_9_io_out_r_stall;
  wire       [15:0]   pe_mat_0_9_io_out_c_data;
  wire                pe_mat_0_9_io_out_c_is_weight;
  wire       [15:0]   pe_mat_0_10_io_out_r_data;
  wire                pe_mat_0_10_io_out_r_stop_weight;
  wire                pe_mat_0_10_io_out_r_stall;
  wire       [15:0]   pe_mat_0_10_io_out_c_data;
  wire                pe_mat_0_10_io_out_c_is_weight;
  wire       [15:0]   pe_mat_0_11_io_out_r_data;
  wire                pe_mat_0_11_io_out_r_stop_weight;
  wire                pe_mat_0_11_io_out_r_stall;
  wire       [15:0]   pe_mat_0_11_io_out_c_data;
  wire                pe_mat_0_11_io_out_c_is_weight;
  wire       [15:0]   pe_mat_0_12_io_out_r_data;
  wire                pe_mat_0_12_io_out_r_stop_weight;
  wire                pe_mat_0_12_io_out_r_stall;
  wire       [15:0]   pe_mat_0_12_io_out_c_data;
  wire                pe_mat_0_12_io_out_c_is_weight;
  wire       [15:0]   pe_mat_0_13_io_out_r_data;
  wire                pe_mat_0_13_io_out_r_stop_weight;
  wire                pe_mat_0_13_io_out_r_stall;
  wire       [15:0]   pe_mat_0_13_io_out_c_data;
  wire                pe_mat_0_13_io_out_c_is_weight;
  wire       [15:0]   pe_mat_0_14_io_out_r_data;
  wire                pe_mat_0_14_io_out_r_stop_weight;
  wire                pe_mat_0_14_io_out_r_stall;
  wire       [15:0]   pe_mat_0_14_io_out_c_data;
  wire                pe_mat_0_14_io_out_c_is_weight;
  wire       [15:0]   pe_mat_0_15_io_out_r_data;
  wire                pe_mat_0_15_io_out_r_stop_weight;
  wire                pe_mat_0_15_io_out_r_stall;
  wire       [15:0]   pe_mat_0_15_io_out_c_data;
  wire                pe_mat_0_15_io_out_c_is_weight;
  wire       [15:0]   pe_mat_0_16_io_out_r_data;
  wire                pe_mat_0_16_io_out_r_stop_weight;
  wire                pe_mat_0_16_io_out_r_stall;
  wire       [15:0]   pe_mat_0_16_io_out_c_data;
  wire                pe_mat_0_16_io_out_c_is_weight;
  wire       [15:0]   pe_mat_0_17_io_out_r_data;
  wire                pe_mat_0_17_io_out_r_stop_weight;
  wire                pe_mat_0_17_io_out_r_stall;
  wire       [15:0]   pe_mat_0_17_io_out_c_data;
  wire                pe_mat_0_17_io_out_c_is_weight;
  wire       [15:0]   pe_mat_0_18_io_out_r_data;
  wire                pe_mat_0_18_io_out_r_stop_weight;
  wire                pe_mat_0_18_io_out_r_stall;
  wire       [15:0]   pe_mat_0_18_io_out_c_data;
  wire                pe_mat_0_18_io_out_c_is_weight;
  wire       [15:0]   pe_mat_0_19_io_out_r_data;
  wire                pe_mat_0_19_io_out_r_stop_weight;
  wire                pe_mat_0_19_io_out_r_stall;
  wire       [15:0]   pe_mat_0_19_io_out_c_data;
  wire                pe_mat_0_19_io_out_c_is_weight;
  wire       [15:0]   pe_mat_0_20_io_out_r_data;
  wire                pe_mat_0_20_io_out_r_stop_weight;
  wire                pe_mat_0_20_io_out_r_stall;
  wire       [15:0]   pe_mat_0_20_io_out_c_data;
  wire                pe_mat_0_20_io_out_c_is_weight;
  wire       [15:0]   pe_mat_0_21_io_out_r_data;
  wire                pe_mat_0_21_io_out_r_stop_weight;
  wire                pe_mat_0_21_io_out_r_stall;
  wire       [15:0]   pe_mat_0_21_io_out_c_data;
  wire                pe_mat_0_21_io_out_c_is_weight;
  wire       [15:0]   pe_mat_0_22_io_out_r_data;
  wire                pe_mat_0_22_io_out_r_stop_weight;
  wire                pe_mat_0_22_io_out_r_stall;
  wire       [15:0]   pe_mat_0_22_io_out_c_data;
  wire                pe_mat_0_22_io_out_c_is_weight;
  wire       [15:0]   pe_mat_0_23_io_out_r_data;
  wire                pe_mat_0_23_io_out_r_stop_weight;
  wire                pe_mat_0_23_io_out_r_stall;
  wire       [15:0]   pe_mat_0_23_io_out_c_data;
  wire                pe_mat_0_23_io_out_c_is_weight;
  wire       [15:0]   pe_mat_0_24_io_out_r_data;
  wire                pe_mat_0_24_io_out_r_stop_weight;
  wire                pe_mat_0_24_io_out_r_stall;
  wire       [15:0]   pe_mat_0_24_io_out_c_data;
  wire                pe_mat_0_24_io_out_c_is_weight;
  wire       [15:0]   pe_mat_0_25_io_out_r_data;
  wire                pe_mat_0_25_io_out_r_stop_weight;
  wire                pe_mat_0_25_io_out_r_stall;
  wire       [15:0]   pe_mat_0_25_io_out_c_data;
  wire                pe_mat_0_25_io_out_c_is_weight;
  wire       [15:0]   pe_mat_0_26_io_out_r_data;
  wire                pe_mat_0_26_io_out_r_stop_weight;
  wire                pe_mat_0_26_io_out_r_stall;
  wire       [15:0]   pe_mat_0_26_io_out_c_data;
  wire                pe_mat_0_26_io_out_c_is_weight;
  wire       [15:0]   pe_mat_0_27_io_out_r_data;
  wire                pe_mat_0_27_io_out_r_stop_weight;
  wire                pe_mat_0_27_io_out_r_stall;
  wire       [15:0]   pe_mat_0_27_io_out_c_data;
  wire                pe_mat_0_27_io_out_c_is_weight;
  wire       [15:0]   pe_mat_0_28_io_out_r_data;
  wire                pe_mat_0_28_io_out_r_stop_weight;
  wire                pe_mat_0_28_io_out_r_stall;
  wire       [15:0]   pe_mat_0_28_io_out_c_data;
  wire                pe_mat_0_28_io_out_c_is_weight;
  wire       [15:0]   pe_mat_0_29_io_out_r_data;
  wire                pe_mat_0_29_io_out_r_stop_weight;
  wire                pe_mat_0_29_io_out_r_stall;
  wire       [15:0]   pe_mat_0_29_io_out_c_data;
  wire                pe_mat_0_29_io_out_c_is_weight;
  wire       [15:0]   pe_mat_0_30_io_out_r_data;
  wire                pe_mat_0_30_io_out_r_stop_weight;
  wire                pe_mat_0_30_io_out_r_stall;
  wire       [15:0]   pe_mat_0_30_io_out_c_data;
  wire                pe_mat_0_30_io_out_c_is_weight;
  wire       [15:0]   pe_mat_0_31_io_out_r_data;
  wire                pe_mat_0_31_io_out_r_stop_weight;
  wire                pe_mat_0_31_io_out_r_stall;
  wire       [15:0]   pe_mat_0_31_io_out_c_data;
  wire                pe_mat_0_31_io_out_c_is_weight;
  wire       [15:0]   pe_mat_1_0_io_out_r_data;
  wire                pe_mat_1_0_io_out_r_stop_weight;
  wire                pe_mat_1_0_io_out_r_stall;
  wire       [15:0]   pe_mat_1_0_io_out_c_data;
  wire                pe_mat_1_0_io_out_c_is_weight;
  wire       [15:0]   pe_mat_1_1_io_out_r_data;
  wire                pe_mat_1_1_io_out_r_stop_weight;
  wire                pe_mat_1_1_io_out_r_stall;
  wire       [15:0]   pe_mat_1_1_io_out_c_data;
  wire                pe_mat_1_1_io_out_c_is_weight;
  wire       [15:0]   pe_mat_1_2_io_out_r_data;
  wire                pe_mat_1_2_io_out_r_stop_weight;
  wire                pe_mat_1_2_io_out_r_stall;
  wire       [15:0]   pe_mat_1_2_io_out_c_data;
  wire                pe_mat_1_2_io_out_c_is_weight;
  wire       [15:0]   pe_mat_1_3_io_out_r_data;
  wire                pe_mat_1_3_io_out_r_stop_weight;
  wire                pe_mat_1_3_io_out_r_stall;
  wire       [15:0]   pe_mat_1_3_io_out_c_data;
  wire                pe_mat_1_3_io_out_c_is_weight;
  wire       [15:0]   pe_mat_1_4_io_out_r_data;
  wire                pe_mat_1_4_io_out_r_stop_weight;
  wire                pe_mat_1_4_io_out_r_stall;
  wire       [15:0]   pe_mat_1_4_io_out_c_data;
  wire                pe_mat_1_4_io_out_c_is_weight;
  wire       [15:0]   pe_mat_1_5_io_out_r_data;
  wire                pe_mat_1_5_io_out_r_stop_weight;
  wire                pe_mat_1_5_io_out_r_stall;
  wire       [15:0]   pe_mat_1_5_io_out_c_data;
  wire                pe_mat_1_5_io_out_c_is_weight;
  wire       [15:0]   pe_mat_1_6_io_out_r_data;
  wire                pe_mat_1_6_io_out_r_stop_weight;
  wire                pe_mat_1_6_io_out_r_stall;
  wire       [15:0]   pe_mat_1_6_io_out_c_data;
  wire                pe_mat_1_6_io_out_c_is_weight;
  wire       [15:0]   pe_mat_1_7_io_out_r_data;
  wire                pe_mat_1_7_io_out_r_stop_weight;
  wire                pe_mat_1_7_io_out_r_stall;
  wire       [15:0]   pe_mat_1_7_io_out_c_data;
  wire                pe_mat_1_7_io_out_c_is_weight;
  wire       [15:0]   pe_mat_1_8_io_out_r_data;
  wire                pe_mat_1_8_io_out_r_stop_weight;
  wire                pe_mat_1_8_io_out_r_stall;
  wire       [15:0]   pe_mat_1_8_io_out_c_data;
  wire                pe_mat_1_8_io_out_c_is_weight;
  wire       [15:0]   pe_mat_1_9_io_out_r_data;
  wire                pe_mat_1_9_io_out_r_stop_weight;
  wire                pe_mat_1_9_io_out_r_stall;
  wire       [15:0]   pe_mat_1_9_io_out_c_data;
  wire                pe_mat_1_9_io_out_c_is_weight;
  wire       [15:0]   pe_mat_1_10_io_out_r_data;
  wire                pe_mat_1_10_io_out_r_stop_weight;
  wire                pe_mat_1_10_io_out_r_stall;
  wire       [15:0]   pe_mat_1_10_io_out_c_data;
  wire                pe_mat_1_10_io_out_c_is_weight;
  wire       [15:0]   pe_mat_1_11_io_out_r_data;
  wire                pe_mat_1_11_io_out_r_stop_weight;
  wire                pe_mat_1_11_io_out_r_stall;
  wire       [15:0]   pe_mat_1_11_io_out_c_data;
  wire                pe_mat_1_11_io_out_c_is_weight;
  wire       [15:0]   pe_mat_1_12_io_out_r_data;
  wire                pe_mat_1_12_io_out_r_stop_weight;
  wire                pe_mat_1_12_io_out_r_stall;
  wire       [15:0]   pe_mat_1_12_io_out_c_data;
  wire                pe_mat_1_12_io_out_c_is_weight;
  wire       [15:0]   pe_mat_1_13_io_out_r_data;
  wire                pe_mat_1_13_io_out_r_stop_weight;
  wire                pe_mat_1_13_io_out_r_stall;
  wire       [15:0]   pe_mat_1_13_io_out_c_data;
  wire                pe_mat_1_13_io_out_c_is_weight;
  wire       [15:0]   pe_mat_1_14_io_out_r_data;
  wire                pe_mat_1_14_io_out_r_stop_weight;
  wire                pe_mat_1_14_io_out_r_stall;
  wire       [15:0]   pe_mat_1_14_io_out_c_data;
  wire                pe_mat_1_14_io_out_c_is_weight;
  wire       [15:0]   pe_mat_1_15_io_out_r_data;
  wire                pe_mat_1_15_io_out_r_stop_weight;
  wire                pe_mat_1_15_io_out_r_stall;
  wire       [15:0]   pe_mat_1_15_io_out_c_data;
  wire                pe_mat_1_15_io_out_c_is_weight;
  wire       [15:0]   pe_mat_1_16_io_out_r_data;
  wire                pe_mat_1_16_io_out_r_stop_weight;
  wire                pe_mat_1_16_io_out_r_stall;
  wire       [15:0]   pe_mat_1_16_io_out_c_data;
  wire                pe_mat_1_16_io_out_c_is_weight;
  wire       [15:0]   pe_mat_1_17_io_out_r_data;
  wire                pe_mat_1_17_io_out_r_stop_weight;
  wire                pe_mat_1_17_io_out_r_stall;
  wire       [15:0]   pe_mat_1_17_io_out_c_data;
  wire                pe_mat_1_17_io_out_c_is_weight;
  wire       [15:0]   pe_mat_1_18_io_out_r_data;
  wire                pe_mat_1_18_io_out_r_stop_weight;
  wire                pe_mat_1_18_io_out_r_stall;
  wire       [15:0]   pe_mat_1_18_io_out_c_data;
  wire                pe_mat_1_18_io_out_c_is_weight;
  wire       [15:0]   pe_mat_1_19_io_out_r_data;
  wire                pe_mat_1_19_io_out_r_stop_weight;
  wire                pe_mat_1_19_io_out_r_stall;
  wire       [15:0]   pe_mat_1_19_io_out_c_data;
  wire                pe_mat_1_19_io_out_c_is_weight;
  wire       [15:0]   pe_mat_1_20_io_out_r_data;
  wire                pe_mat_1_20_io_out_r_stop_weight;
  wire                pe_mat_1_20_io_out_r_stall;
  wire       [15:0]   pe_mat_1_20_io_out_c_data;
  wire                pe_mat_1_20_io_out_c_is_weight;
  wire       [15:0]   pe_mat_1_21_io_out_r_data;
  wire                pe_mat_1_21_io_out_r_stop_weight;
  wire                pe_mat_1_21_io_out_r_stall;
  wire       [15:0]   pe_mat_1_21_io_out_c_data;
  wire                pe_mat_1_21_io_out_c_is_weight;
  wire       [15:0]   pe_mat_1_22_io_out_r_data;
  wire                pe_mat_1_22_io_out_r_stop_weight;
  wire                pe_mat_1_22_io_out_r_stall;
  wire       [15:0]   pe_mat_1_22_io_out_c_data;
  wire                pe_mat_1_22_io_out_c_is_weight;
  wire       [15:0]   pe_mat_1_23_io_out_r_data;
  wire                pe_mat_1_23_io_out_r_stop_weight;
  wire                pe_mat_1_23_io_out_r_stall;
  wire       [15:0]   pe_mat_1_23_io_out_c_data;
  wire                pe_mat_1_23_io_out_c_is_weight;
  wire       [15:0]   pe_mat_1_24_io_out_r_data;
  wire                pe_mat_1_24_io_out_r_stop_weight;
  wire                pe_mat_1_24_io_out_r_stall;
  wire       [15:0]   pe_mat_1_24_io_out_c_data;
  wire                pe_mat_1_24_io_out_c_is_weight;
  wire       [15:0]   pe_mat_1_25_io_out_r_data;
  wire                pe_mat_1_25_io_out_r_stop_weight;
  wire                pe_mat_1_25_io_out_r_stall;
  wire       [15:0]   pe_mat_1_25_io_out_c_data;
  wire                pe_mat_1_25_io_out_c_is_weight;
  wire       [15:0]   pe_mat_1_26_io_out_r_data;
  wire                pe_mat_1_26_io_out_r_stop_weight;
  wire                pe_mat_1_26_io_out_r_stall;
  wire       [15:0]   pe_mat_1_26_io_out_c_data;
  wire                pe_mat_1_26_io_out_c_is_weight;
  wire       [15:0]   pe_mat_1_27_io_out_r_data;
  wire                pe_mat_1_27_io_out_r_stop_weight;
  wire                pe_mat_1_27_io_out_r_stall;
  wire       [15:0]   pe_mat_1_27_io_out_c_data;
  wire                pe_mat_1_27_io_out_c_is_weight;
  wire       [15:0]   pe_mat_1_28_io_out_r_data;
  wire                pe_mat_1_28_io_out_r_stop_weight;
  wire                pe_mat_1_28_io_out_r_stall;
  wire       [15:0]   pe_mat_1_28_io_out_c_data;
  wire                pe_mat_1_28_io_out_c_is_weight;
  wire       [15:0]   pe_mat_1_29_io_out_r_data;
  wire                pe_mat_1_29_io_out_r_stop_weight;
  wire                pe_mat_1_29_io_out_r_stall;
  wire       [15:0]   pe_mat_1_29_io_out_c_data;
  wire                pe_mat_1_29_io_out_c_is_weight;
  wire       [15:0]   pe_mat_1_30_io_out_r_data;
  wire                pe_mat_1_30_io_out_r_stop_weight;
  wire                pe_mat_1_30_io_out_r_stall;
  wire       [15:0]   pe_mat_1_30_io_out_c_data;
  wire                pe_mat_1_30_io_out_c_is_weight;
  wire       [15:0]   pe_mat_1_31_io_out_r_data;
  wire                pe_mat_1_31_io_out_r_stop_weight;
  wire                pe_mat_1_31_io_out_r_stall;
  wire       [15:0]   pe_mat_1_31_io_out_c_data;
  wire                pe_mat_1_31_io_out_c_is_weight;
  wire       [15:0]   pe_mat_2_0_io_out_r_data;
  wire                pe_mat_2_0_io_out_r_stop_weight;
  wire                pe_mat_2_0_io_out_r_stall;
  wire       [15:0]   pe_mat_2_0_io_out_c_data;
  wire                pe_mat_2_0_io_out_c_is_weight;
  wire       [15:0]   pe_mat_2_1_io_out_r_data;
  wire                pe_mat_2_1_io_out_r_stop_weight;
  wire                pe_mat_2_1_io_out_r_stall;
  wire       [15:0]   pe_mat_2_1_io_out_c_data;
  wire                pe_mat_2_1_io_out_c_is_weight;
  wire       [15:0]   pe_mat_2_2_io_out_r_data;
  wire                pe_mat_2_2_io_out_r_stop_weight;
  wire                pe_mat_2_2_io_out_r_stall;
  wire       [15:0]   pe_mat_2_2_io_out_c_data;
  wire                pe_mat_2_2_io_out_c_is_weight;
  wire       [15:0]   pe_mat_2_3_io_out_r_data;
  wire                pe_mat_2_3_io_out_r_stop_weight;
  wire                pe_mat_2_3_io_out_r_stall;
  wire       [15:0]   pe_mat_2_3_io_out_c_data;
  wire                pe_mat_2_3_io_out_c_is_weight;
  wire       [15:0]   pe_mat_2_4_io_out_r_data;
  wire                pe_mat_2_4_io_out_r_stop_weight;
  wire                pe_mat_2_4_io_out_r_stall;
  wire       [15:0]   pe_mat_2_4_io_out_c_data;
  wire                pe_mat_2_4_io_out_c_is_weight;
  wire       [15:0]   pe_mat_2_5_io_out_r_data;
  wire                pe_mat_2_5_io_out_r_stop_weight;
  wire                pe_mat_2_5_io_out_r_stall;
  wire       [15:0]   pe_mat_2_5_io_out_c_data;
  wire                pe_mat_2_5_io_out_c_is_weight;
  wire       [15:0]   pe_mat_2_6_io_out_r_data;
  wire                pe_mat_2_6_io_out_r_stop_weight;
  wire                pe_mat_2_6_io_out_r_stall;
  wire       [15:0]   pe_mat_2_6_io_out_c_data;
  wire                pe_mat_2_6_io_out_c_is_weight;
  wire       [15:0]   pe_mat_2_7_io_out_r_data;
  wire                pe_mat_2_7_io_out_r_stop_weight;
  wire                pe_mat_2_7_io_out_r_stall;
  wire       [15:0]   pe_mat_2_7_io_out_c_data;
  wire                pe_mat_2_7_io_out_c_is_weight;
  wire       [15:0]   pe_mat_2_8_io_out_r_data;
  wire                pe_mat_2_8_io_out_r_stop_weight;
  wire                pe_mat_2_8_io_out_r_stall;
  wire       [15:0]   pe_mat_2_8_io_out_c_data;
  wire                pe_mat_2_8_io_out_c_is_weight;
  wire       [15:0]   pe_mat_2_9_io_out_r_data;
  wire                pe_mat_2_9_io_out_r_stop_weight;
  wire                pe_mat_2_9_io_out_r_stall;
  wire       [15:0]   pe_mat_2_9_io_out_c_data;
  wire                pe_mat_2_9_io_out_c_is_weight;
  wire       [15:0]   pe_mat_2_10_io_out_r_data;
  wire                pe_mat_2_10_io_out_r_stop_weight;
  wire                pe_mat_2_10_io_out_r_stall;
  wire       [15:0]   pe_mat_2_10_io_out_c_data;
  wire                pe_mat_2_10_io_out_c_is_weight;
  wire       [15:0]   pe_mat_2_11_io_out_r_data;
  wire                pe_mat_2_11_io_out_r_stop_weight;
  wire                pe_mat_2_11_io_out_r_stall;
  wire       [15:0]   pe_mat_2_11_io_out_c_data;
  wire                pe_mat_2_11_io_out_c_is_weight;
  wire       [15:0]   pe_mat_2_12_io_out_r_data;
  wire                pe_mat_2_12_io_out_r_stop_weight;
  wire                pe_mat_2_12_io_out_r_stall;
  wire       [15:0]   pe_mat_2_12_io_out_c_data;
  wire                pe_mat_2_12_io_out_c_is_weight;
  wire       [15:0]   pe_mat_2_13_io_out_r_data;
  wire                pe_mat_2_13_io_out_r_stop_weight;
  wire                pe_mat_2_13_io_out_r_stall;
  wire       [15:0]   pe_mat_2_13_io_out_c_data;
  wire                pe_mat_2_13_io_out_c_is_weight;
  wire       [15:0]   pe_mat_2_14_io_out_r_data;
  wire                pe_mat_2_14_io_out_r_stop_weight;
  wire                pe_mat_2_14_io_out_r_stall;
  wire       [15:0]   pe_mat_2_14_io_out_c_data;
  wire                pe_mat_2_14_io_out_c_is_weight;
  wire       [15:0]   pe_mat_2_15_io_out_r_data;
  wire                pe_mat_2_15_io_out_r_stop_weight;
  wire                pe_mat_2_15_io_out_r_stall;
  wire       [15:0]   pe_mat_2_15_io_out_c_data;
  wire                pe_mat_2_15_io_out_c_is_weight;
  wire       [15:0]   pe_mat_2_16_io_out_r_data;
  wire                pe_mat_2_16_io_out_r_stop_weight;
  wire                pe_mat_2_16_io_out_r_stall;
  wire       [15:0]   pe_mat_2_16_io_out_c_data;
  wire                pe_mat_2_16_io_out_c_is_weight;
  wire       [15:0]   pe_mat_2_17_io_out_r_data;
  wire                pe_mat_2_17_io_out_r_stop_weight;
  wire                pe_mat_2_17_io_out_r_stall;
  wire       [15:0]   pe_mat_2_17_io_out_c_data;
  wire                pe_mat_2_17_io_out_c_is_weight;
  wire       [15:0]   pe_mat_2_18_io_out_r_data;
  wire                pe_mat_2_18_io_out_r_stop_weight;
  wire                pe_mat_2_18_io_out_r_stall;
  wire       [15:0]   pe_mat_2_18_io_out_c_data;
  wire                pe_mat_2_18_io_out_c_is_weight;
  wire       [15:0]   pe_mat_2_19_io_out_r_data;
  wire                pe_mat_2_19_io_out_r_stop_weight;
  wire                pe_mat_2_19_io_out_r_stall;
  wire       [15:0]   pe_mat_2_19_io_out_c_data;
  wire                pe_mat_2_19_io_out_c_is_weight;
  wire       [15:0]   pe_mat_2_20_io_out_r_data;
  wire                pe_mat_2_20_io_out_r_stop_weight;
  wire                pe_mat_2_20_io_out_r_stall;
  wire       [15:0]   pe_mat_2_20_io_out_c_data;
  wire                pe_mat_2_20_io_out_c_is_weight;
  wire       [15:0]   pe_mat_2_21_io_out_r_data;
  wire                pe_mat_2_21_io_out_r_stop_weight;
  wire                pe_mat_2_21_io_out_r_stall;
  wire       [15:0]   pe_mat_2_21_io_out_c_data;
  wire                pe_mat_2_21_io_out_c_is_weight;
  wire       [15:0]   pe_mat_2_22_io_out_r_data;
  wire                pe_mat_2_22_io_out_r_stop_weight;
  wire                pe_mat_2_22_io_out_r_stall;
  wire       [15:0]   pe_mat_2_22_io_out_c_data;
  wire                pe_mat_2_22_io_out_c_is_weight;
  wire       [15:0]   pe_mat_2_23_io_out_r_data;
  wire                pe_mat_2_23_io_out_r_stop_weight;
  wire                pe_mat_2_23_io_out_r_stall;
  wire       [15:0]   pe_mat_2_23_io_out_c_data;
  wire                pe_mat_2_23_io_out_c_is_weight;
  wire       [15:0]   pe_mat_2_24_io_out_r_data;
  wire                pe_mat_2_24_io_out_r_stop_weight;
  wire                pe_mat_2_24_io_out_r_stall;
  wire       [15:0]   pe_mat_2_24_io_out_c_data;
  wire                pe_mat_2_24_io_out_c_is_weight;
  wire       [15:0]   pe_mat_2_25_io_out_r_data;
  wire                pe_mat_2_25_io_out_r_stop_weight;
  wire                pe_mat_2_25_io_out_r_stall;
  wire       [15:0]   pe_mat_2_25_io_out_c_data;
  wire                pe_mat_2_25_io_out_c_is_weight;
  wire       [15:0]   pe_mat_2_26_io_out_r_data;
  wire                pe_mat_2_26_io_out_r_stop_weight;
  wire                pe_mat_2_26_io_out_r_stall;
  wire       [15:0]   pe_mat_2_26_io_out_c_data;
  wire                pe_mat_2_26_io_out_c_is_weight;
  wire       [15:0]   pe_mat_2_27_io_out_r_data;
  wire                pe_mat_2_27_io_out_r_stop_weight;
  wire                pe_mat_2_27_io_out_r_stall;
  wire       [15:0]   pe_mat_2_27_io_out_c_data;
  wire                pe_mat_2_27_io_out_c_is_weight;
  wire       [15:0]   pe_mat_2_28_io_out_r_data;
  wire                pe_mat_2_28_io_out_r_stop_weight;
  wire                pe_mat_2_28_io_out_r_stall;
  wire       [15:0]   pe_mat_2_28_io_out_c_data;
  wire                pe_mat_2_28_io_out_c_is_weight;
  wire       [15:0]   pe_mat_2_29_io_out_r_data;
  wire                pe_mat_2_29_io_out_r_stop_weight;
  wire                pe_mat_2_29_io_out_r_stall;
  wire       [15:0]   pe_mat_2_29_io_out_c_data;
  wire                pe_mat_2_29_io_out_c_is_weight;
  wire       [15:0]   pe_mat_2_30_io_out_r_data;
  wire                pe_mat_2_30_io_out_r_stop_weight;
  wire                pe_mat_2_30_io_out_r_stall;
  wire       [15:0]   pe_mat_2_30_io_out_c_data;
  wire                pe_mat_2_30_io_out_c_is_weight;
  wire       [15:0]   pe_mat_2_31_io_out_r_data;
  wire                pe_mat_2_31_io_out_r_stop_weight;
  wire                pe_mat_2_31_io_out_r_stall;
  wire       [15:0]   pe_mat_2_31_io_out_c_data;
  wire                pe_mat_2_31_io_out_c_is_weight;
  wire       [15:0]   pe_mat_3_0_io_out_r_data;
  wire                pe_mat_3_0_io_out_r_stop_weight;
  wire                pe_mat_3_0_io_out_r_stall;
  wire       [15:0]   pe_mat_3_0_io_out_c_data;
  wire                pe_mat_3_0_io_out_c_is_weight;
  wire       [15:0]   pe_mat_3_1_io_out_r_data;
  wire                pe_mat_3_1_io_out_r_stop_weight;
  wire                pe_mat_3_1_io_out_r_stall;
  wire       [15:0]   pe_mat_3_1_io_out_c_data;
  wire                pe_mat_3_1_io_out_c_is_weight;
  wire       [15:0]   pe_mat_3_2_io_out_r_data;
  wire                pe_mat_3_2_io_out_r_stop_weight;
  wire                pe_mat_3_2_io_out_r_stall;
  wire       [15:0]   pe_mat_3_2_io_out_c_data;
  wire                pe_mat_3_2_io_out_c_is_weight;
  wire       [15:0]   pe_mat_3_3_io_out_r_data;
  wire                pe_mat_3_3_io_out_r_stop_weight;
  wire                pe_mat_3_3_io_out_r_stall;
  wire       [15:0]   pe_mat_3_3_io_out_c_data;
  wire                pe_mat_3_3_io_out_c_is_weight;
  wire       [15:0]   pe_mat_3_4_io_out_r_data;
  wire                pe_mat_3_4_io_out_r_stop_weight;
  wire                pe_mat_3_4_io_out_r_stall;
  wire       [15:0]   pe_mat_3_4_io_out_c_data;
  wire                pe_mat_3_4_io_out_c_is_weight;
  wire       [15:0]   pe_mat_3_5_io_out_r_data;
  wire                pe_mat_3_5_io_out_r_stop_weight;
  wire                pe_mat_3_5_io_out_r_stall;
  wire       [15:0]   pe_mat_3_5_io_out_c_data;
  wire                pe_mat_3_5_io_out_c_is_weight;
  wire       [15:0]   pe_mat_3_6_io_out_r_data;
  wire                pe_mat_3_6_io_out_r_stop_weight;
  wire                pe_mat_3_6_io_out_r_stall;
  wire       [15:0]   pe_mat_3_6_io_out_c_data;
  wire                pe_mat_3_6_io_out_c_is_weight;
  wire       [15:0]   pe_mat_3_7_io_out_r_data;
  wire                pe_mat_3_7_io_out_r_stop_weight;
  wire                pe_mat_3_7_io_out_r_stall;
  wire       [15:0]   pe_mat_3_7_io_out_c_data;
  wire                pe_mat_3_7_io_out_c_is_weight;
  wire       [15:0]   pe_mat_3_8_io_out_r_data;
  wire                pe_mat_3_8_io_out_r_stop_weight;
  wire                pe_mat_3_8_io_out_r_stall;
  wire       [15:0]   pe_mat_3_8_io_out_c_data;
  wire                pe_mat_3_8_io_out_c_is_weight;
  wire       [15:0]   pe_mat_3_9_io_out_r_data;
  wire                pe_mat_3_9_io_out_r_stop_weight;
  wire                pe_mat_3_9_io_out_r_stall;
  wire       [15:0]   pe_mat_3_9_io_out_c_data;
  wire                pe_mat_3_9_io_out_c_is_weight;
  wire       [15:0]   pe_mat_3_10_io_out_r_data;
  wire                pe_mat_3_10_io_out_r_stop_weight;
  wire                pe_mat_3_10_io_out_r_stall;
  wire       [15:0]   pe_mat_3_10_io_out_c_data;
  wire                pe_mat_3_10_io_out_c_is_weight;
  wire       [15:0]   pe_mat_3_11_io_out_r_data;
  wire                pe_mat_3_11_io_out_r_stop_weight;
  wire                pe_mat_3_11_io_out_r_stall;
  wire       [15:0]   pe_mat_3_11_io_out_c_data;
  wire                pe_mat_3_11_io_out_c_is_weight;
  wire       [15:0]   pe_mat_3_12_io_out_r_data;
  wire                pe_mat_3_12_io_out_r_stop_weight;
  wire                pe_mat_3_12_io_out_r_stall;
  wire       [15:0]   pe_mat_3_12_io_out_c_data;
  wire                pe_mat_3_12_io_out_c_is_weight;
  wire       [15:0]   pe_mat_3_13_io_out_r_data;
  wire                pe_mat_3_13_io_out_r_stop_weight;
  wire                pe_mat_3_13_io_out_r_stall;
  wire       [15:0]   pe_mat_3_13_io_out_c_data;
  wire                pe_mat_3_13_io_out_c_is_weight;
  wire       [15:0]   pe_mat_3_14_io_out_r_data;
  wire                pe_mat_3_14_io_out_r_stop_weight;
  wire                pe_mat_3_14_io_out_r_stall;
  wire       [15:0]   pe_mat_3_14_io_out_c_data;
  wire                pe_mat_3_14_io_out_c_is_weight;
  wire       [15:0]   pe_mat_3_15_io_out_r_data;
  wire                pe_mat_3_15_io_out_r_stop_weight;
  wire                pe_mat_3_15_io_out_r_stall;
  wire       [15:0]   pe_mat_3_15_io_out_c_data;
  wire                pe_mat_3_15_io_out_c_is_weight;
  wire       [15:0]   pe_mat_3_16_io_out_r_data;
  wire                pe_mat_3_16_io_out_r_stop_weight;
  wire                pe_mat_3_16_io_out_r_stall;
  wire       [15:0]   pe_mat_3_16_io_out_c_data;
  wire                pe_mat_3_16_io_out_c_is_weight;
  wire       [15:0]   pe_mat_3_17_io_out_r_data;
  wire                pe_mat_3_17_io_out_r_stop_weight;
  wire                pe_mat_3_17_io_out_r_stall;
  wire       [15:0]   pe_mat_3_17_io_out_c_data;
  wire                pe_mat_3_17_io_out_c_is_weight;
  wire       [15:0]   pe_mat_3_18_io_out_r_data;
  wire                pe_mat_3_18_io_out_r_stop_weight;
  wire                pe_mat_3_18_io_out_r_stall;
  wire       [15:0]   pe_mat_3_18_io_out_c_data;
  wire                pe_mat_3_18_io_out_c_is_weight;
  wire       [15:0]   pe_mat_3_19_io_out_r_data;
  wire                pe_mat_3_19_io_out_r_stop_weight;
  wire                pe_mat_3_19_io_out_r_stall;
  wire       [15:0]   pe_mat_3_19_io_out_c_data;
  wire                pe_mat_3_19_io_out_c_is_weight;
  wire       [15:0]   pe_mat_3_20_io_out_r_data;
  wire                pe_mat_3_20_io_out_r_stop_weight;
  wire                pe_mat_3_20_io_out_r_stall;
  wire       [15:0]   pe_mat_3_20_io_out_c_data;
  wire                pe_mat_3_20_io_out_c_is_weight;
  wire       [15:0]   pe_mat_3_21_io_out_r_data;
  wire                pe_mat_3_21_io_out_r_stop_weight;
  wire                pe_mat_3_21_io_out_r_stall;
  wire       [15:0]   pe_mat_3_21_io_out_c_data;
  wire                pe_mat_3_21_io_out_c_is_weight;
  wire       [15:0]   pe_mat_3_22_io_out_r_data;
  wire                pe_mat_3_22_io_out_r_stop_weight;
  wire                pe_mat_3_22_io_out_r_stall;
  wire       [15:0]   pe_mat_3_22_io_out_c_data;
  wire                pe_mat_3_22_io_out_c_is_weight;
  wire       [15:0]   pe_mat_3_23_io_out_r_data;
  wire                pe_mat_3_23_io_out_r_stop_weight;
  wire                pe_mat_3_23_io_out_r_stall;
  wire       [15:0]   pe_mat_3_23_io_out_c_data;
  wire                pe_mat_3_23_io_out_c_is_weight;
  wire       [15:0]   pe_mat_3_24_io_out_r_data;
  wire                pe_mat_3_24_io_out_r_stop_weight;
  wire                pe_mat_3_24_io_out_r_stall;
  wire       [15:0]   pe_mat_3_24_io_out_c_data;
  wire                pe_mat_3_24_io_out_c_is_weight;
  wire       [15:0]   pe_mat_3_25_io_out_r_data;
  wire                pe_mat_3_25_io_out_r_stop_weight;
  wire                pe_mat_3_25_io_out_r_stall;
  wire       [15:0]   pe_mat_3_25_io_out_c_data;
  wire                pe_mat_3_25_io_out_c_is_weight;
  wire       [15:0]   pe_mat_3_26_io_out_r_data;
  wire                pe_mat_3_26_io_out_r_stop_weight;
  wire                pe_mat_3_26_io_out_r_stall;
  wire       [15:0]   pe_mat_3_26_io_out_c_data;
  wire                pe_mat_3_26_io_out_c_is_weight;
  wire       [15:0]   pe_mat_3_27_io_out_r_data;
  wire                pe_mat_3_27_io_out_r_stop_weight;
  wire                pe_mat_3_27_io_out_r_stall;
  wire       [15:0]   pe_mat_3_27_io_out_c_data;
  wire                pe_mat_3_27_io_out_c_is_weight;
  wire       [15:0]   pe_mat_3_28_io_out_r_data;
  wire                pe_mat_3_28_io_out_r_stop_weight;
  wire                pe_mat_3_28_io_out_r_stall;
  wire       [15:0]   pe_mat_3_28_io_out_c_data;
  wire                pe_mat_3_28_io_out_c_is_weight;
  wire       [15:0]   pe_mat_3_29_io_out_r_data;
  wire                pe_mat_3_29_io_out_r_stop_weight;
  wire                pe_mat_3_29_io_out_r_stall;
  wire       [15:0]   pe_mat_3_29_io_out_c_data;
  wire                pe_mat_3_29_io_out_c_is_weight;
  wire       [15:0]   pe_mat_3_30_io_out_r_data;
  wire                pe_mat_3_30_io_out_r_stop_weight;
  wire                pe_mat_3_30_io_out_r_stall;
  wire       [15:0]   pe_mat_3_30_io_out_c_data;
  wire                pe_mat_3_30_io_out_c_is_weight;
  wire       [15:0]   pe_mat_3_31_io_out_r_data;
  wire                pe_mat_3_31_io_out_r_stop_weight;
  wire                pe_mat_3_31_io_out_r_stall;
  wire       [15:0]   pe_mat_3_31_io_out_c_data;
  wire                pe_mat_3_31_io_out_c_is_weight;
  wire       [15:0]   pe_mat_4_0_io_out_r_data;
  wire                pe_mat_4_0_io_out_r_stop_weight;
  wire                pe_mat_4_0_io_out_r_stall;
  wire       [15:0]   pe_mat_4_0_io_out_c_data;
  wire                pe_mat_4_0_io_out_c_is_weight;
  wire       [15:0]   pe_mat_4_1_io_out_r_data;
  wire                pe_mat_4_1_io_out_r_stop_weight;
  wire                pe_mat_4_1_io_out_r_stall;
  wire       [15:0]   pe_mat_4_1_io_out_c_data;
  wire                pe_mat_4_1_io_out_c_is_weight;
  wire       [15:0]   pe_mat_4_2_io_out_r_data;
  wire                pe_mat_4_2_io_out_r_stop_weight;
  wire                pe_mat_4_2_io_out_r_stall;
  wire       [15:0]   pe_mat_4_2_io_out_c_data;
  wire                pe_mat_4_2_io_out_c_is_weight;
  wire       [15:0]   pe_mat_4_3_io_out_r_data;
  wire                pe_mat_4_3_io_out_r_stop_weight;
  wire                pe_mat_4_3_io_out_r_stall;
  wire       [15:0]   pe_mat_4_3_io_out_c_data;
  wire                pe_mat_4_3_io_out_c_is_weight;
  wire       [15:0]   pe_mat_4_4_io_out_r_data;
  wire                pe_mat_4_4_io_out_r_stop_weight;
  wire                pe_mat_4_4_io_out_r_stall;
  wire       [15:0]   pe_mat_4_4_io_out_c_data;
  wire                pe_mat_4_4_io_out_c_is_weight;
  wire       [15:0]   pe_mat_4_5_io_out_r_data;
  wire                pe_mat_4_5_io_out_r_stop_weight;
  wire                pe_mat_4_5_io_out_r_stall;
  wire       [15:0]   pe_mat_4_5_io_out_c_data;
  wire                pe_mat_4_5_io_out_c_is_weight;
  wire       [15:0]   pe_mat_4_6_io_out_r_data;
  wire                pe_mat_4_6_io_out_r_stop_weight;
  wire                pe_mat_4_6_io_out_r_stall;
  wire       [15:0]   pe_mat_4_6_io_out_c_data;
  wire                pe_mat_4_6_io_out_c_is_weight;
  wire       [15:0]   pe_mat_4_7_io_out_r_data;
  wire                pe_mat_4_7_io_out_r_stop_weight;
  wire                pe_mat_4_7_io_out_r_stall;
  wire       [15:0]   pe_mat_4_7_io_out_c_data;
  wire                pe_mat_4_7_io_out_c_is_weight;
  wire       [15:0]   pe_mat_4_8_io_out_r_data;
  wire                pe_mat_4_8_io_out_r_stop_weight;
  wire                pe_mat_4_8_io_out_r_stall;
  wire       [15:0]   pe_mat_4_8_io_out_c_data;
  wire                pe_mat_4_8_io_out_c_is_weight;
  wire       [15:0]   pe_mat_4_9_io_out_r_data;
  wire                pe_mat_4_9_io_out_r_stop_weight;
  wire                pe_mat_4_9_io_out_r_stall;
  wire       [15:0]   pe_mat_4_9_io_out_c_data;
  wire                pe_mat_4_9_io_out_c_is_weight;
  wire       [15:0]   pe_mat_4_10_io_out_r_data;
  wire                pe_mat_4_10_io_out_r_stop_weight;
  wire                pe_mat_4_10_io_out_r_stall;
  wire       [15:0]   pe_mat_4_10_io_out_c_data;
  wire                pe_mat_4_10_io_out_c_is_weight;
  wire       [15:0]   pe_mat_4_11_io_out_r_data;
  wire                pe_mat_4_11_io_out_r_stop_weight;
  wire                pe_mat_4_11_io_out_r_stall;
  wire       [15:0]   pe_mat_4_11_io_out_c_data;
  wire                pe_mat_4_11_io_out_c_is_weight;
  wire       [15:0]   pe_mat_4_12_io_out_r_data;
  wire                pe_mat_4_12_io_out_r_stop_weight;
  wire                pe_mat_4_12_io_out_r_stall;
  wire       [15:0]   pe_mat_4_12_io_out_c_data;
  wire                pe_mat_4_12_io_out_c_is_weight;
  wire       [15:0]   pe_mat_4_13_io_out_r_data;
  wire                pe_mat_4_13_io_out_r_stop_weight;
  wire                pe_mat_4_13_io_out_r_stall;
  wire       [15:0]   pe_mat_4_13_io_out_c_data;
  wire                pe_mat_4_13_io_out_c_is_weight;
  wire       [15:0]   pe_mat_4_14_io_out_r_data;
  wire                pe_mat_4_14_io_out_r_stop_weight;
  wire                pe_mat_4_14_io_out_r_stall;
  wire       [15:0]   pe_mat_4_14_io_out_c_data;
  wire                pe_mat_4_14_io_out_c_is_weight;
  wire       [15:0]   pe_mat_4_15_io_out_r_data;
  wire                pe_mat_4_15_io_out_r_stop_weight;
  wire                pe_mat_4_15_io_out_r_stall;
  wire       [15:0]   pe_mat_4_15_io_out_c_data;
  wire                pe_mat_4_15_io_out_c_is_weight;
  wire       [15:0]   pe_mat_4_16_io_out_r_data;
  wire                pe_mat_4_16_io_out_r_stop_weight;
  wire                pe_mat_4_16_io_out_r_stall;
  wire       [15:0]   pe_mat_4_16_io_out_c_data;
  wire                pe_mat_4_16_io_out_c_is_weight;
  wire       [15:0]   pe_mat_4_17_io_out_r_data;
  wire                pe_mat_4_17_io_out_r_stop_weight;
  wire                pe_mat_4_17_io_out_r_stall;
  wire       [15:0]   pe_mat_4_17_io_out_c_data;
  wire                pe_mat_4_17_io_out_c_is_weight;
  wire       [15:0]   pe_mat_4_18_io_out_r_data;
  wire                pe_mat_4_18_io_out_r_stop_weight;
  wire                pe_mat_4_18_io_out_r_stall;
  wire       [15:0]   pe_mat_4_18_io_out_c_data;
  wire                pe_mat_4_18_io_out_c_is_weight;
  wire       [15:0]   pe_mat_4_19_io_out_r_data;
  wire                pe_mat_4_19_io_out_r_stop_weight;
  wire                pe_mat_4_19_io_out_r_stall;
  wire       [15:0]   pe_mat_4_19_io_out_c_data;
  wire                pe_mat_4_19_io_out_c_is_weight;
  wire       [15:0]   pe_mat_4_20_io_out_r_data;
  wire                pe_mat_4_20_io_out_r_stop_weight;
  wire                pe_mat_4_20_io_out_r_stall;
  wire       [15:0]   pe_mat_4_20_io_out_c_data;
  wire                pe_mat_4_20_io_out_c_is_weight;
  wire       [15:0]   pe_mat_4_21_io_out_r_data;
  wire                pe_mat_4_21_io_out_r_stop_weight;
  wire                pe_mat_4_21_io_out_r_stall;
  wire       [15:0]   pe_mat_4_21_io_out_c_data;
  wire                pe_mat_4_21_io_out_c_is_weight;
  wire       [15:0]   pe_mat_4_22_io_out_r_data;
  wire                pe_mat_4_22_io_out_r_stop_weight;
  wire                pe_mat_4_22_io_out_r_stall;
  wire       [15:0]   pe_mat_4_22_io_out_c_data;
  wire                pe_mat_4_22_io_out_c_is_weight;
  wire       [15:0]   pe_mat_4_23_io_out_r_data;
  wire                pe_mat_4_23_io_out_r_stop_weight;
  wire                pe_mat_4_23_io_out_r_stall;
  wire       [15:0]   pe_mat_4_23_io_out_c_data;
  wire                pe_mat_4_23_io_out_c_is_weight;
  wire       [15:0]   pe_mat_4_24_io_out_r_data;
  wire                pe_mat_4_24_io_out_r_stop_weight;
  wire                pe_mat_4_24_io_out_r_stall;
  wire       [15:0]   pe_mat_4_24_io_out_c_data;
  wire                pe_mat_4_24_io_out_c_is_weight;
  wire       [15:0]   pe_mat_4_25_io_out_r_data;
  wire                pe_mat_4_25_io_out_r_stop_weight;
  wire                pe_mat_4_25_io_out_r_stall;
  wire       [15:0]   pe_mat_4_25_io_out_c_data;
  wire                pe_mat_4_25_io_out_c_is_weight;
  wire       [15:0]   pe_mat_4_26_io_out_r_data;
  wire                pe_mat_4_26_io_out_r_stop_weight;
  wire                pe_mat_4_26_io_out_r_stall;
  wire       [15:0]   pe_mat_4_26_io_out_c_data;
  wire                pe_mat_4_26_io_out_c_is_weight;
  wire       [15:0]   pe_mat_4_27_io_out_r_data;
  wire                pe_mat_4_27_io_out_r_stop_weight;
  wire                pe_mat_4_27_io_out_r_stall;
  wire       [15:0]   pe_mat_4_27_io_out_c_data;
  wire                pe_mat_4_27_io_out_c_is_weight;
  wire       [15:0]   pe_mat_4_28_io_out_r_data;
  wire                pe_mat_4_28_io_out_r_stop_weight;
  wire                pe_mat_4_28_io_out_r_stall;
  wire       [15:0]   pe_mat_4_28_io_out_c_data;
  wire                pe_mat_4_28_io_out_c_is_weight;
  wire       [15:0]   pe_mat_4_29_io_out_r_data;
  wire                pe_mat_4_29_io_out_r_stop_weight;
  wire                pe_mat_4_29_io_out_r_stall;
  wire       [15:0]   pe_mat_4_29_io_out_c_data;
  wire                pe_mat_4_29_io_out_c_is_weight;
  wire       [15:0]   pe_mat_4_30_io_out_r_data;
  wire                pe_mat_4_30_io_out_r_stop_weight;
  wire                pe_mat_4_30_io_out_r_stall;
  wire       [15:0]   pe_mat_4_30_io_out_c_data;
  wire                pe_mat_4_30_io_out_c_is_weight;
  wire       [15:0]   pe_mat_4_31_io_out_r_data;
  wire                pe_mat_4_31_io_out_r_stop_weight;
  wire                pe_mat_4_31_io_out_r_stall;
  wire       [15:0]   pe_mat_4_31_io_out_c_data;
  wire                pe_mat_4_31_io_out_c_is_weight;
  wire       [15:0]   pe_mat_5_0_io_out_r_data;
  wire                pe_mat_5_0_io_out_r_stop_weight;
  wire                pe_mat_5_0_io_out_r_stall;
  wire       [15:0]   pe_mat_5_0_io_out_c_data;
  wire                pe_mat_5_0_io_out_c_is_weight;
  wire       [15:0]   pe_mat_5_1_io_out_r_data;
  wire                pe_mat_5_1_io_out_r_stop_weight;
  wire                pe_mat_5_1_io_out_r_stall;
  wire       [15:0]   pe_mat_5_1_io_out_c_data;
  wire                pe_mat_5_1_io_out_c_is_weight;
  wire       [15:0]   pe_mat_5_2_io_out_r_data;
  wire                pe_mat_5_2_io_out_r_stop_weight;
  wire                pe_mat_5_2_io_out_r_stall;
  wire       [15:0]   pe_mat_5_2_io_out_c_data;
  wire                pe_mat_5_2_io_out_c_is_weight;
  wire       [15:0]   pe_mat_5_3_io_out_r_data;
  wire                pe_mat_5_3_io_out_r_stop_weight;
  wire                pe_mat_5_3_io_out_r_stall;
  wire       [15:0]   pe_mat_5_3_io_out_c_data;
  wire                pe_mat_5_3_io_out_c_is_weight;
  wire       [15:0]   pe_mat_5_4_io_out_r_data;
  wire                pe_mat_5_4_io_out_r_stop_weight;
  wire                pe_mat_5_4_io_out_r_stall;
  wire       [15:0]   pe_mat_5_4_io_out_c_data;
  wire                pe_mat_5_4_io_out_c_is_weight;
  wire       [15:0]   pe_mat_5_5_io_out_r_data;
  wire                pe_mat_5_5_io_out_r_stop_weight;
  wire                pe_mat_5_5_io_out_r_stall;
  wire       [15:0]   pe_mat_5_5_io_out_c_data;
  wire                pe_mat_5_5_io_out_c_is_weight;
  wire       [15:0]   pe_mat_5_6_io_out_r_data;
  wire                pe_mat_5_6_io_out_r_stop_weight;
  wire                pe_mat_5_6_io_out_r_stall;
  wire       [15:0]   pe_mat_5_6_io_out_c_data;
  wire                pe_mat_5_6_io_out_c_is_weight;
  wire       [15:0]   pe_mat_5_7_io_out_r_data;
  wire                pe_mat_5_7_io_out_r_stop_weight;
  wire                pe_mat_5_7_io_out_r_stall;
  wire       [15:0]   pe_mat_5_7_io_out_c_data;
  wire                pe_mat_5_7_io_out_c_is_weight;
  wire       [15:0]   pe_mat_5_8_io_out_r_data;
  wire                pe_mat_5_8_io_out_r_stop_weight;
  wire                pe_mat_5_8_io_out_r_stall;
  wire       [15:0]   pe_mat_5_8_io_out_c_data;
  wire                pe_mat_5_8_io_out_c_is_weight;
  wire       [15:0]   pe_mat_5_9_io_out_r_data;
  wire                pe_mat_5_9_io_out_r_stop_weight;
  wire                pe_mat_5_9_io_out_r_stall;
  wire       [15:0]   pe_mat_5_9_io_out_c_data;
  wire                pe_mat_5_9_io_out_c_is_weight;
  wire       [15:0]   pe_mat_5_10_io_out_r_data;
  wire                pe_mat_5_10_io_out_r_stop_weight;
  wire                pe_mat_5_10_io_out_r_stall;
  wire       [15:0]   pe_mat_5_10_io_out_c_data;
  wire                pe_mat_5_10_io_out_c_is_weight;
  wire       [15:0]   pe_mat_5_11_io_out_r_data;
  wire                pe_mat_5_11_io_out_r_stop_weight;
  wire                pe_mat_5_11_io_out_r_stall;
  wire       [15:0]   pe_mat_5_11_io_out_c_data;
  wire                pe_mat_5_11_io_out_c_is_weight;
  wire       [15:0]   pe_mat_5_12_io_out_r_data;
  wire                pe_mat_5_12_io_out_r_stop_weight;
  wire                pe_mat_5_12_io_out_r_stall;
  wire       [15:0]   pe_mat_5_12_io_out_c_data;
  wire                pe_mat_5_12_io_out_c_is_weight;
  wire       [15:0]   pe_mat_5_13_io_out_r_data;
  wire                pe_mat_5_13_io_out_r_stop_weight;
  wire                pe_mat_5_13_io_out_r_stall;
  wire       [15:0]   pe_mat_5_13_io_out_c_data;
  wire                pe_mat_5_13_io_out_c_is_weight;
  wire       [15:0]   pe_mat_5_14_io_out_r_data;
  wire                pe_mat_5_14_io_out_r_stop_weight;
  wire                pe_mat_5_14_io_out_r_stall;
  wire       [15:0]   pe_mat_5_14_io_out_c_data;
  wire                pe_mat_5_14_io_out_c_is_weight;
  wire       [15:0]   pe_mat_5_15_io_out_r_data;
  wire                pe_mat_5_15_io_out_r_stop_weight;
  wire                pe_mat_5_15_io_out_r_stall;
  wire       [15:0]   pe_mat_5_15_io_out_c_data;
  wire                pe_mat_5_15_io_out_c_is_weight;
  wire       [15:0]   pe_mat_5_16_io_out_r_data;
  wire                pe_mat_5_16_io_out_r_stop_weight;
  wire                pe_mat_5_16_io_out_r_stall;
  wire       [15:0]   pe_mat_5_16_io_out_c_data;
  wire                pe_mat_5_16_io_out_c_is_weight;
  wire       [15:0]   pe_mat_5_17_io_out_r_data;
  wire                pe_mat_5_17_io_out_r_stop_weight;
  wire                pe_mat_5_17_io_out_r_stall;
  wire       [15:0]   pe_mat_5_17_io_out_c_data;
  wire                pe_mat_5_17_io_out_c_is_weight;
  wire       [15:0]   pe_mat_5_18_io_out_r_data;
  wire                pe_mat_5_18_io_out_r_stop_weight;
  wire                pe_mat_5_18_io_out_r_stall;
  wire       [15:0]   pe_mat_5_18_io_out_c_data;
  wire                pe_mat_5_18_io_out_c_is_weight;
  wire       [15:0]   pe_mat_5_19_io_out_r_data;
  wire                pe_mat_5_19_io_out_r_stop_weight;
  wire                pe_mat_5_19_io_out_r_stall;
  wire       [15:0]   pe_mat_5_19_io_out_c_data;
  wire                pe_mat_5_19_io_out_c_is_weight;
  wire       [15:0]   pe_mat_5_20_io_out_r_data;
  wire                pe_mat_5_20_io_out_r_stop_weight;
  wire                pe_mat_5_20_io_out_r_stall;
  wire       [15:0]   pe_mat_5_20_io_out_c_data;
  wire                pe_mat_5_20_io_out_c_is_weight;
  wire       [15:0]   pe_mat_5_21_io_out_r_data;
  wire                pe_mat_5_21_io_out_r_stop_weight;
  wire                pe_mat_5_21_io_out_r_stall;
  wire       [15:0]   pe_mat_5_21_io_out_c_data;
  wire                pe_mat_5_21_io_out_c_is_weight;
  wire       [15:0]   pe_mat_5_22_io_out_r_data;
  wire                pe_mat_5_22_io_out_r_stop_weight;
  wire                pe_mat_5_22_io_out_r_stall;
  wire       [15:0]   pe_mat_5_22_io_out_c_data;
  wire                pe_mat_5_22_io_out_c_is_weight;
  wire       [15:0]   pe_mat_5_23_io_out_r_data;
  wire                pe_mat_5_23_io_out_r_stop_weight;
  wire                pe_mat_5_23_io_out_r_stall;
  wire       [15:0]   pe_mat_5_23_io_out_c_data;
  wire                pe_mat_5_23_io_out_c_is_weight;
  wire       [15:0]   pe_mat_5_24_io_out_r_data;
  wire                pe_mat_5_24_io_out_r_stop_weight;
  wire                pe_mat_5_24_io_out_r_stall;
  wire       [15:0]   pe_mat_5_24_io_out_c_data;
  wire                pe_mat_5_24_io_out_c_is_weight;
  wire       [15:0]   pe_mat_5_25_io_out_r_data;
  wire                pe_mat_5_25_io_out_r_stop_weight;
  wire                pe_mat_5_25_io_out_r_stall;
  wire       [15:0]   pe_mat_5_25_io_out_c_data;
  wire                pe_mat_5_25_io_out_c_is_weight;
  wire       [15:0]   pe_mat_5_26_io_out_r_data;
  wire                pe_mat_5_26_io_out_r_stop_weight;
  wire                pe_mat_5_26_io_out_r_stall;
  wire       [15:0]   pe_mat_5_26_io_out_c_data;
  wire                pe_mat_5_26_io_out_c_is_weight;
  wire       [15:0]   pe_mat_5_27_io_out_r_data;
  wire                pe_mat_5_27_io_out_r_stop_weight;
  wire                pe_mat_5_27_io_out_r_stall;
  wire       [15:0]   pe_mat_5_27_io_out_c_data;
  wire                pe_mat_5_27_io_out_c_is_weight;
  wire       [15:0]   pe_mat_5_28_io_out_r_data;
  wire                pe_mat_5_28_io_out_r_stop_weight;
  wire                pe_mat_5_28_io_out_r_stall;
  wire       [15:0]   pe_mat_5_28_io_out_c_data;
  wire                pe_mat_5_28_io_out_c_is_weight;
  wire       [15:0]   pe_mat_5_29_io_out_r_data;
  wire                pe_mat_5_29_io_out_r_stop_weight;
  wire                pe_mat_5_29_io_out_r_stall;
  wire       [15:0]   pe_mat_5_29_io_out_c_data;
  wire                pe_mat_5_29_io_out_c_is_weight;
  wire       [15:0]   pe_mat_5_30_io_out_r_data;
  wire                pe_mat_5_30_io_out_r_stop_weight;
  wire                pe_mat_5_30_io_out_r_stall;
  wire       [15:0]   pe_mat_5_30_io_out_c_data;
  wire                pe_mat_5_30_io_out_c_is_weight;
  wire       [15:0]   pe_mat_5_31_io_out_r_data;
  wire                pe_mat_5_31_io_out_r_stop_weight;
  wire                pe_mat_5_31_io_out_r_stall;
  wire       [15:0]   pe_mat_5_31_io_out_c_data;
  wire                pe_mat_5_31_io_out_c_is_weight;
  wire       [15:0]   pe_mat_6_0_io_out_r_data;
  wire                pe_mat_6_0_io_out_r_stop_weight;
  wire                pe_mat_6_0_io_out_r_stall;
  wire       [15:0]   pe_mat_6_0_io_out_c_data;
  wire                pe_mat_6_0_io_out_c_is_weight;
  wire       [15:0]   pe_mat_6_1_io_out_r_data;
  wire                pe_mat_6_1_io_out_r_stop_weight;
  wire                pe_mat_6_1_io_out_r_stall;
  wire       [15:0]   pe_mat_6_1_io_out_c_data;
  wire                pe_mat_6_1_io_out_c_is_weight;
  wire       [15:0]   pe_mat_6_2_io_out_r_data;
  wire                pe_mat_6_2_io_out_r_stop_weight;
  wire                pe_mat_6_2_io_out_r_stall;
  wire       [15:0]   pe_mat_6_2_io_out_c_data;
  wire                pe_mat_6_2_io_out_c_is_weight;
  wire       [15:0]   pe_mat_6_3_io_out_r_data;
  wire                pe_mat_6_3_io_out_r_stop_weight;
  wire                pe_mat_6_3_io_out_r_stall;
  wire       [15:0]   pe_mat_6_3_io_out_c_data;
  wire                pe_mat_6_3_io_out_c_is_weight;
  wire       [15:0]   pe_mat_6_4_io_out_r_data;
  wire                pe_mat_6_4_io_out_r_stop_weight;
  wire                pe_mat_6_4_io_out_r_stall;
  wire       [15:0]   pe_mat_6_4_io_out_c_data;
  wire                pe_mat_6_4_io_out_c_is_weight;
  wire       [15:0]   pe_mat_6_5_io_out_r_data;
  wire                pe_mat_6_5_io_out_r_stop_weight;
  wire                pe_mat_6_5_io_out_r_stall;
  wire       [15:0]   pe_mat_6_5_io_out_c_data;
  wire                pe_mat_6_5_io_out_c_is_weight;
  wire       [15:0]   pe_mat_6_6_io_out_r_data;
  wire                pe_mat_6_6_io_out_r_stop_weight;
  wire                pe_mat_6_6_io_out_r_stall;
  wire       [15:0]   pe_mat_6_6_io_out_c_data;
  wire                pe_mat_6_6_io_out_c_is_weight;
  wire       [15:0]   pe_mat_6_7_io_out_r_data;
  wire                pe_mat_6_7_io_out_r_stop_weight;
  wire                pe_mat_6_7_io_out_r_stall;
  wire       [15:0]   pe_mat_6_7_io_out_c_data;
  wire                pe_mat_6_7_io_out_c_is_weight;
  wire       [15:0]   pe_mat_6_8_io_out_r_data;
  wire                pe_mat_6_8_io_out_r_stop_weight;
  wire                pe_mat_6_8_io_out_r_stall;
  wire       [15:0]   pe_mat_6_8_io_out_c_data;
  wire                pe_mat_6_8_io_out_c_is_weight;
  wire       [15:0]   pe_mat_6_9_io_out_r_data;
  wire                pe_mat_6_9_io_out_r_stop_weight;
  wire                pe_mat_6_9_io_out_r_stall;
  wire       [15:0]   pe_mat_6_9_io_out_c_data;
  wire                pe_mat_6_9_io_out_c_is_weight;
  wire       [15:0]   pe_mat_6_10_io_out_r_data;
  wire                pe_mat_6_10_io_out_r_stop_weight;
  wire                pe_mat_6_10_io_out_r_stall;
  wire       [15:0]   pe_mat_6_10_io_out_c_data;
  wire                pe_mat_6_10_io_out_c_is_weight;
  wire       [15:0]   pe_mat_6_11_io_out_r_data;
  wire                pe_mat_6_11_io_out_r_stop_weight;
  wire                pe_mat_6_11_io_out_r_stall;
  wire       [15:0]   pe_mat_6_11_io_out_c_data;
  wire                pe_mat_6_11_io_out_c_is_weight;
  wire       [15:0]   pe_mat_6_12_io_out_r_data;
  wire                pe_mat_6_12_io_out_r_stop_weight;
  wire                pe_mat_6_12_io_out_r_stall;
  wire       [15:0]   pe_mat_6_12_io_out_c_data;
  wire                pe_mat_6_12_io_out_c_is_weight;
  wire       [15:0]   pe_mat_6_13_io_out_r_data;
  wire                pe_mat_6_13_io_out_r_stop_weight;
  wire                pe_mat_6_13_io_out_r_stall;
  wire       [15:0]   pe_mat_6_13_io_out_c_data;
  wire                pe_mat_6_13_io_out_c_is_weight;
  wire       [15:0]   pe_mat_6_14_io_out_r_data;
  wire                pe_mat_6_14_io_out_r_stop_weight;
  wire                pe_mat_6_14_io_out_r_stall;
  wire       [15:0]   pe_mat_6_14_io_out_c_data;
  wire                pe_mat_6_14_io_out_c_is_weight;
  wire       [15:0]   pe_mat_6_15_io_out_r_data;
  wire                pe_mat_6_15_io_out_r_stop_weight;
  wire                pe_mat_6_15_io_out_r_stall;
  wire       [15:0]   pe_mat_6_15_io_out_c_data;
  wire                pe_mat_6_15_io_out_c_is_weight;
  wire       [15:0]   pe_mat_6_16_io_out_r_data;
  wire                pe_mat_6_16_io_out_r_stop_weight;
  wire                pe_mat_6_16_io_out_r_stall;
  wire       [15:0]   pe_mat_6_16_io_out_c_data;
  wire                pe_mat_6_16_io_out_c_is_weight;
  wire       [15:0]   pe_mat_6_17_io_out_r_data;
  wire                pe_mat_6_17_io_out_r_stop_weight;
  wire                pe_mat_6_17_io_out_r_stall;
  wire       [15:0]   pe_mat_6_17_io_out_c_data;
  wire                pe_mat_6_17_io_out_c_is_weight;
  wire       [15:0]   pe_mat_6_18_io_out_r_data;
  wire                pe_mat_6_18_io_out_r_stop_weight;
  wire                pe_mat_6_18_io_out_r_stall;
  wire       [15:0]   pe_mat_6_18_io_out_c_data;
  wire                pe_mat_6_18_io_out_c_is_weight;
  wire       [15:0]   pe_mat_6_19_io_out_r_data;
  wire                pe_mat_6_19_io_out_r_stop_weight;
  wire                pe_mat_6_19_io_out_r_stall;
  wire       [15:0]   pe_mat_6_19_io_out_c_data;
  wire                pe_mat_6_19_io_out_c_is_weight;
  wire       [15:0]   pe_mat_6_20_io_out_r_data;
  wire                pe_mat_6_20_io_out_r_stop_weight;
  wire                pe_mat_6_20_io_out_r_stall;
  wire       [15:0]   pe_mat_6_20_io_out_c_data;
  wire                pe_mat_6_20_io_out_c_is_weight;
  wire       [15:0]   pe_mat_6_21_io_out_r_data;
  wire                pe_mat_6_21_io_out_r_stop_weight;
  wire                pe_mat_6_21_io_out_r_stall;
  wire       [15:0]   pe_mat_6_21_io_out_c_data;
  wire                pe_mat_6_21_io_out_c_is_weight;
  wire       [15:0]   pe_mat_6_22_io_out_r_data;
  wire                pe_mat_6_22_io_out_r_stop_weight;
  wire                pe_mat_6_22_io_out_r_stall;
  wire       [15:0]   pe_mat_6_22_io_out_c_data;
  wire                pe_mat_6_22_io_out_c_is_weight;
  wire       [15:0]   pe_mat_6_23_io_out_r_data;
  wire                pe_mat_6_23_io_out_r_stop_weight;
  wire                pe_mat_6_23_io_out_r_stall;
  wire       [15:0]   pe_mat_6_23_io_out_c_data;
  wire                pe_mat_6_23_io_out_c_is_weight;
  wire       [15:0]   pe_mat_6_24_io_out_r_data;
  wire                pe_mat_6_24_io_out_r_stop_weight;
  wire                pe_mat_6_24_io_out_r_stall;
  wire       [15:0]   pe_mat_6_24_io_out_c_data;
  wire                pe_mat_6_24_io_out_c_is_weight;
  wire       [15:0]   pe_mat_6_25_io_out_r_data;
  wire                pe_mat_6_25_io_out_r_stop_weight;
  wire                pe_mat_6_25_io_out_r_stall;
  wire       [15:0]   pe_mat_6_25_io_out_c_data;
  wire                pe_mat_6_25_io_out_c_is_weight;
  wire       [15:0]   pe_mat_6_26_io_out_r_data;
  wire                pe_mat_6_26_io_out_r_stop_weight;
  wire                pe_mat_6_26_io_out_r_stall;
  wire       [15:0]   pe_mat_6_26_io_out_c_data;
  wire                pe_mat_6_26_io_out_c_is_weight;
  wire       [15:0]   pe_mat_6_27_io_out_r_data;
  wire                pe_mat_6_27_io_out_r_stop_weight;
  wire                pe_mat_6_27_io_out_r_stall;
  wire       [15:0]   pe_mat_6_27_io_out_c_data;
  wire                pe_mat_6_27_io_out_c_is_weight;
  wire       [15:0]   pe_mat_6_28_io_out_r_data;
  wire                pe_mat_6_28_io_out_r_stop_weight;
  wire                pe_mat_6_28_io_out_r_stall;
  wire       [15:0]   pe_mat_6_28_io_out_c_data;
  wire                pe_mat_6_28_io_out_c_is_weight;
  wire       [15:0]   pe_mat_6_29_io_out_r_data;
  wire                pe_mat_6_29_io_out_r_stop_weight;
  wire                pe_mat_6_29_io_out_r_stall;
  wire       [15:0]   pe_mat_6_29_io_out_c_data;
  wire                pe_mat_6_29_io_out_c_is_weight;
  wire       [15:0]   pe_mat_6_30_io_out_r_data;
  wire                pe_mat_6_30_io_out_r_stop_weight;
  wire                pe_mat_6_30_io_out_r_stall;
  wire       [15:0]   pe_mat_6_30_io_out_c_data;
  wire                pe_mat_6_30_io_out_c_is_weight;
  wire       [15:0]   pe_mat_6_31_io_out_r_data;
  wire                pe_mat_6_31_io_out_r_stop_weight;
  wire                pe_mat_6_31_io_out_r_stall;
  wire       [15:0]   pe_mat_6_31_io_out_c_data;
  wire                pe_mat_6_31_io_out_c_is_weight;
  wire       [15:0]   pe_mat_7_0_io_out_r_data;
  wire                pe_mat_7_0_io_out_r_stop_weight;
  wire                pe_mat_7_0_io_out_r_stall;
  wire       [15:0]   pe_mat_7_0_io_out_c_data;
  wire                pe_mat_7_0_io_out_c_is_weight;
  wire       [15:0]   pe_mat_7_1_io_out_r_data;
  wire                pe_mat_7_1_io_out_r_stop_weight;
  wire                pe_mat_7_1_io_out_r_stall;
  wire       [15:0]   pe_mat_7_1_io_out_c_data;
  wire                pe_mat_7_1_io_out_c_is_weight;
  wire       [15:0]   pe_mat_7_2_io_out_r_data;
  wire                pe_mat_7_2_io_out_r_stop_weight;
  wire                pe_mat_7_2_io_out_r_stall;
  wire       [15:0]   pe_mat_7_2_io_out_c_data;
  wire                pe_mat_7_2_io_out_c_is_weight;
  wire       [15:0]   pe_mat_7_3_io_out_r_data;
  wire                pe_mat_7_3_io_out_r_stop_weight;
  wire                pe_mat_7_3_io_out_r_stall;
  wire       [15:0]   pe_mat_7_3_io_out_c_data;
  wire                pe_mat_7_3_io_out_c_is_weight;
  wire       [15:0]   pe_mat_7_4_io_out_r_data;
  wire                pe_mat_7_4_io_out_r_stop_weight;
  wire                pe_mat_7_4_io_out_r_stall;
  wire       [15:0]   pe_mat_7_4_io_out_c_data;
  wire                pe_mat_7_4_io_out_c_is_weight;
  wire       [15:0]   pe_mat_7_5_io_out_r_data;
  wire                pe_mat_7_5_io_out_r_stop_weight;
  wire                pe_mat_7_5_io_out_r_stall;
  wire       [15:0]   pe_mat_7_5_io_out_c_data;
  wire                pe_mat_7_5_io_out_c_is_weight;
  wire       [15:0]   pe_mat_7_6_io_out_r_data;
  wire                pe_mat_7_6_io_out_r_stop_weight;
  wire                pe_mat_7_6_io_out_r_stall;
  wire       [15:0]   pe_mat_7_6_io_out_c_data;
  wire                pe_mat_7_6_io_out_c_is_weight;
  wire       [15:0]   pe_mat_7_7_io_out_r_data;
  wire                pe_mat_7_7_io_out_r_stop_weight;
  wire                pe_mat_7_7_io_out_r_stall;
  wire       [15:0]   pe_mat_7_7_io_out_c_data;
  wire                pe_mat_7_7_io_out_c_is_weight;
  wire       [15:0]   pe_mat_7_8_io_out_r_data;
  wire                pe_mat_7_8_io_out_r_stop_weight;
  wire                pe_mat_7_8_io_out_r_stall;
  wire       [15:0]   pe_mat_7_8_io_out_c_data;
  wire                pe_mat_7_8_io_out_c_is_weight;
  wire       [15:0]   pe_mat_7_9_io_out_r_data;
  wire                pe_mat_7_9_io_out_r_stop_weight;
  wire                pe_mat_7_9_io_out_r_stall;
  wire       [15:0]   pe_mat_7_9_io_out_c_data;
  wire                pe_mat_7_9_io_out_c_is_weight;
  wire       [15:0]   pe_mat_7_10_io_out_r_data;
  wire                pe_mat_7_10_io_out_r_stop_weight;
  wire                pe_mat_7_10_io_out_r_stall;
  wire       [15:0]   pe_mat_7_10_io_out_c_data;
  wire                pe_mat_7_10_io_out_c_is_weight;
  wire       [15:0]   pe_mat_7_11_io_out_r_data;
  wire                pe_mat_7_11_io_out_r_stop_weight;
  wire                pe_mat_7_11_io_out_r_stall;
  wire       [15:0]   pe_mat_7_11_io_out_c_data;
  wire                pe_mat_7_11_io_out_c_is_weight;
  wire       [15:0]   pe_mat_7_12_io_out_r_data;
  wire                pe_mat_7_12_io_out_r_stop_weight;
  wire                pe_mat_7_12_io_out_r_stall;
  wire       [15:0]   pe_mat_7_12_io_out_c_data;
  wire                pe_mat_7_12_io_out_c_is_weight;
  wire       [15:0]   pe_mat_7_13_io_out_r_data;
  wire                pe_mat_7_13_io_out_r_stop_weight;
  wire                pe_mat_7_13_io_out_r_stall;
  wire       [15:0]   pe_mat_7_13_io_out_c_data;
  wire                pe_mat_7_13_io_out_c_is_weight;
  wire       [15:0]   pe_mat_7_14_io_out_r_data;
  wire                pe_mat_7_14_io_out_r_stop_weight;
  wire                pe_mat_7_14_io_out_r_stall;
  wire       [15:0]   pe_mat_7_14_io_out_c_data;
  wire                pe_mat_7_14_io_out_c_is_weight;
  wire       [15:0]   pe_mat_7_15_io_out_r_data;
  wire                pe_mat_7_15_io_out_r_stop_weight;
  wire                pe_mat_7_15_io_out_r_stall;
  wire       [15:0]   pe_mat_7_15_io_out_c_data;
  wire                pe_mat_7_15_io_out_c_is_weight;
  wire       [15:0]   pe_mat_7_16_io_out_r_data;
  wire                pe_mat_7_16_io_out_r_stop_weight;
  wire                pe_mat_7_16_io_out_r_stall;
  wire       [15:0]   pe_mat_7_16_io_out_c_data;
  wire                pe_mat_7_16_io_out_c_is_weight;
  wire       [15:0]   pe_mat_7_17_io_out_r_data;
  wire                pe_mat_7_17_io_out_r_stop_weight;
  wire                pe_mat_7_17_io_out_r_stall;
  wire       [15:0]   pe_mat_7_17_io_out_c_data;
  wire                pe_mat_7_17_io_out_c_is_weight;
  wire       [15:0]   pe_mat_7_18_io_out_r_data;
  wire                pe_mat_7_18_io_out_r_stop_weight;
  wire                pe_mat_7_18_io_out_r_stall;
  wire       [15:0]   pe_mat_7_18_io_out_c_data;
  wire                pe_mat_7_18_io_out_c_is_weight;
  wire       [15:0]   pe_mat_7_19_io_out_r_data;
  wire                pe_mat_7_19_io_out_r_stop_weight;
  wire                pe_mat_7_19_io_out_r_stall;
  wire       [15:0]   pe_mat_7_19_io_out_c_data;
  wire                pe_mat_7_19_io_out_c_is_weight;
  wire       [15:0]   pe_mat_7_20_io_out_r_data;
  wire                pe_mat_7_20_io_out_r_stop_weight;
  wire                pe_mat_7_20_io_out_r_stall;
  wire       [15:0]   pe_mat_7_20_io_out_c_data;
  wire                pe_mat_7_20_io_out_c_is_weight;
  wire       [15:0]   pe_mat_7_21_io_out_r_data;
  wire                pe_mat_7_21_io_out_r_stop_weight;
  wire                pe_mat_7_21_io_out_r_stall;
  wire       [15:0]   pe_mat_7_21_io_out_c_data;
  wire                pe_mat_7_21_io_out_c_is_weight;
  wire       [15:0]   pe_mat_7_22_io_out_r_data;
  wire                pe_mat_7_22_io_out_r_stop_weight;
  wire                pe_mat_7_22_io_out_r_stall;
  wire       [15:0]   pe_mat_7_22_io_out_c_data;
  wire                pe_mat_7_22_io_out_c_is_weight;
  wire       [15:0]   pe_mat_7_23_io_out_r_data;
  wire                pe_mat_7_23_io_out_r_stop_weight;
  wire                pe_mat_7_23_io_out_r_stall;
  wire       [15:0]   pe_mat_7_23_io_out_c_data;
  wire                pe_mat_7_23_io_out_c_is_weight;
  wire       [15:0]   pe_mat_7_24_io_out_r_data;
  wire                pe_mat_7_24_io_out_r_stop_weight;
  wire                pe_mat_7_24_io_out_r_stall;
  wire       [15:0]   pe_mat_7_24_io_out_c_data;
  wire                pe_mat_7_24_io_out_c_is_weight;
  wire       [15:0]   pe_mat_7_25_io_out_r_data;
  wire                pe_mat_7_25_io_out_r_stop_weight;
  wire                pe_mat_7_25_io_out_r_stall;
  wire       [15:0]   pe_mat_7_25_io_out_c_data;
  wire                pe_mat_7_25_io_out_c_is_weight;
  wire       [15:0]   pe_mat_7_26_io_out_r_data;
  wire                pe_mat_7_26_io_out_r_stop_weight;
  wire                pe_mat_7_26_io_out_r_stall;
  wire       [15:0]   pe_mat_7_26_io_out_c_data;
  wire                pe_mat_7_26_io_out_c_is_weight;
  wire       [15:0]   pe_mat_7_27_io_out_r_data;
  wire                pe_mat_7_27_io_out_r_stop_weight;
  wire                pe_mat_7_27_io_out_r_stall;
  wire       [15:0]   pe_mat_7_27_io_out_c_data;
  wire                pe_mat_7_27_io_out_c_is_weight;
  wire       [15:0]   pe_mat_7_28_io_out_r_data;
  wire                pe_mat_7_28_io_out_r_stop_weight;
  wire                pe_mat_7_28_io_out_r_stall;
  wire       [15:0]   pe_mat_7_28_io_out_c_data;
  wire                pe_mat_7_28_io_out_c_is_weight;
  wire       [15:0]   pe_mat_7_29_io_out_r_data;
  wire                pe_mat_7_29_io_out_r_stop_weight;
  wire                pe_mat_7_29_io_out_r_stall;
  wire       [15:0]   pe_mat_7_29_io_out_c_data;
  wire                pe_mat_7_29_io_out_c_is_weight;
  wire       [15:0]   pe_mat_7_30_io_out_r_data;
  wire                pe_mat_7_30_io_out_r_stop_weight;
  wire                pe_mat_7_30_io_out_r_stall;
  wire       [15:0]   pe_mat_7_30_io_out_c_data;
  wire                pe_mat_7_30_io_out_c_is_weight;
  wire       [15:0]   pe_mat_7_31_io_out_r_data;
  wire                pe_mat_7_31_io_out_r_stop_weight;
  wire                pe_mat_7_31_io_out_r_stall;
  wire       [15:0]   pe_mat_7_31_io_out_c_data;
  wire                pe_mat_7_31_io_out_c_is_weight;
  wire       [15:0]   pe_mat_8_0_io_out_r_data;
  wire                pe_mat_8_0_io_out_r_stop_weight;
  wire                pe_mat_8_0_io_out_r_stall;
  wire       [15:0]   pe_mat_8_0_io_out_c_data;
  wire                pe_mat_8_0_io_out_c_is_weight;
  wire       [15:0]   pe_mat_8_1_io_out_r_data;
  wire                pe_mat_8_1_io_out_r_stop_weight;
  wire                pe_mat_8_1_io_out_r_stall;
  wire       [15:0]   pe_mat_8_1_io_out_c_data;
  wire                pe_mat_8_1_io_out_c_is_weight;
  wire       [15:0]   pe_mat_8_2_io_out_r_data;
  wire                pe_mat_8_2_io_out_r_stop_weight;
  wire                pe_mat_8_2_io_out_r_stall;
  wire       [15:0]   pe_mat_8_2_io_out_c_data;
  wire                pe_mat_8_2_io_out_c_is_weight;
  wire       [15:0]   pe_mat_8_3_io_out_r_data;
  wire                pe_mat_8_3_io_out_r_stop_weight;
  wire                pe_mat_8_3_io_out_r_stall;
  wire       [15:0]   pe_mat_8_3_io_out_c_data;
  wire                pe_mat_8_3_io_out_c_is_weight;
  wire       [15:0]   pe_mat_8_4_io_out_r_data;
  wire                pe_mat_8_4_io_out_r_stop_weight;
  wire                pe_mat_8_4_io_out_r_stall;
  wire       [15:0]   pe_mat_8_4_io_out_c_data;
  wire                pe_mat_8_4_io_out_c_is_weight;
  wire       [15:0]   pe_mat_8_5_io_out_r_data;
  wire                pe_mat_8_5_io_out_r_stop_weight;
  wire                pe_mat_8_5_io_out_r_stall;
  wire       [15:0]   pe_mat_8_5_io_out_c_data;
  wire                pe_mat_8_5_io_out_c_is_weight;
  wire       [15:0]   pe_mat_8_6_io_out_r_data;
  wire                pe_mat_8_6_io_out_r_stop_weight;
  wire                pe_mat_8_6_io_out_r_stall;
  wire       [15:0]   pe_mat_8_6_io_out_c_data;
  wire                pe_mat_8_6_io_out_c_is_weight;
  wire       [15:0]   pe_mat_8_7_io_out_r_data;
  wire                pe_mat_8_7_io_out_r_stop_weight;
  wire                pe_mat_8_7_io_out_r_stall;
  wire       [15:0]   pe_mat_8_7_io_out_c_data;
  wire                pe_mat_8_7_io_out_c_is_weight;
  wire       [15:0]   pe_mat_8_8_io_out_r_data;
  wire                pe_mat_8_8_io_out_r_stop_weight;
  wire                pe_mat_8_8_io_out_r_stall;
  wire       [15:0]   pe_mat_8_8_io_out_c_data;
  wire                pe_mat_8_8_io_out_c_is_weight;
  wire       [15:0]   pe_mat_8_9_io_out_r_data;
  wire                pe_mat_8_9_io_out_r_stop_weight;
  wire                pe_mat_8_9_io_out_r_stall;
  wire       [15:0]   pe_mat_8_9_io_out_c_data;
  wire                pe_mat_8_9_io_out_c_is_weight;
  wire       [15:0]   pe_mat_8_10_io_out_r_data;
  wire                pe_mat_8_10_io_out_r_stop_weight;
  wire                pe_mat_8_10_io_out_r_stall;
  wire       [15:0]   pe_mat_8_10_io_out_c_data;
  wire                pe_mat_8_10_io_out_c_is_weight;
  wire       [15:0]   pe_mat_8_11_io_out_r_data;
  wire                pe_mat_8_11_io_out_r_stop_weight;
  wire                pe_mat_8_11_io_out_r_stall;
  wire       [15:0]   pe_mat_8_11_io_out_c_data;
  wire                pe_mat_8_11_io_out_c_is_weight;
  wire       [15:0]   pe_mat_8_12_io_out_r_data;
  wire                pe_mat_8_12_io_out_r_stop_weight;
  wire                pe_mat_8_12_io_out_r_stall;
  wire       [15:0]   pe_mat_8_12_io_out_c_data;
  wire                pe_mat_8_12_io_out_c_is_weight;
  wire       [15:0]   pe_mat_8_13_io_out_r_data;
  wire                pe_mat_8_13_io_out_r_stop_weight;
  wire                pe_mat_8_13_io_out_r_stall;
  wire       [15:0]   pe_mat_8_13_io_out_c_data;
  wire                pe_mat_8_13_io_out_c_is_weight;
  wire       [15:0]   pe_mat_8_14_io_out_r_data;
  wire                pe_mat_8_14_io_out_r_stop_weight;
  wire                pe_mat_8_14_io_out_r_stall;
  wire       [15:0]   pe_mat_8_14_io_out_c_data;
  wire                pe_mat_8_14_io_out_c_is_weight;
  wire       [15:0]   pe_mat_8_15_io_out_r_data;
  wire                pe_mat_8_15_io_out_r_stop_weight;
  wire                pe_mat_8_15_io_out_r_stall;
  wire       [15:0]   pe_mat_8_15_io_out_c_data;
  wire                pe_mat_8_15_io_out_c_is_weight;
  wire       [15:0]   pe_mat_8_16_io_out_r_data;
  wire                pe_mat_8_16_io_out_r_stop_weight;
  wire                pe_mat_8_16_io_out_r_stall;
  wire       [15:0]   pe_mat_8_16_io_out_c_data;
  wire                pe_mat_8_16_io_out_c_is_weight;
  wire       [15:0]   pe_mat_8_17_io_out_r_data;
  wire                pe_mat_8_17_io_out_r_stop_weight;
  wire                pe_mat_8_17_io_out_r_stall;
  wire       [15:0]   pe_mat_8_17_io_out_c_data;
  wire                pe_mat_8_17_io_out_c_is_weight;
  wire       [15:0]   pe_mat_8_18_io_out_r_data;
  wire                pe_mat_8_18_io_out_r_stop_weight;
  wire                pe_mat_8_18_io_out_r_stall;
  wire       [15:0]   pe_mat_8_18_io_out_c_data;
  wire                pe_mat_8_18_io_out_c_is_weight;
  wire       [15:0]   pe_mat_8_19_io_out_r_data;
  wire                pe_mat_8_19_io_out_r_stop_weight;
  wire                pe_mat_8_19_io_out_r_stall;
  wire       [15:0]   pe_mat_8_19_io_out_c_data;
  wire                pe_mat_8_19_io_out_c_is_weight;
  wire       [15:0]   pe_mat_8_20_io_out_r_data;
  wire                pe_mat_8_20_io_out_r_stop_weight;
  wire                pe_mat_8_20_io_out_r_stall;
  wire       [15:0]   pe_mat_8_20_io_out_c_data;
  wire                pe_mat_8_20_io_out_c_is_weight;
  wire       [15:0]   pe_mat_8_21_io_out_r_data;
  wire                pe_mat_8_21_io_out_r_stop_weight;
  wire                pe_mat_8_21_io_out_r_stall;
  wire       [15:0]   pe_mat_8_21_io_out_c_data;
  wire                pe_mat_8_21_io_out_c_is_weight;
  wire       [15:0]   pe_mat_8_22_io_out_r_data;
  wire                pe_mat_8_22_io_out_r_stop_weight;
  wire                pe_mat_8_22_io_out_r_stall;
  wire       [15:0]   pe_mat_8_22_io_out_c_data;
  wire                pe_mat_8_22_io_out_c_is_weight;
  wire       [15:0]   pe_mat_8_23_io_out_r_data;
  wire                pe_mat_8_23_io_out_r_stop_weight;
  wire                pe_mat_8_23_io_out_r_stall;
  wire       [15:0]   pe_mat_8_23_io_out_c_data;
  wire                pe_mat_8_23_io_out_c_is_weight;
  wire       [15:0]   pe_mat_8_24_io_out_r_data;
  wire                pe_mat_8_24_io_out_r_stop_weight;
  wire                pe_mat_8_24_io_out_r_stall;
  wire       [15:0]   pe_mat_8_24_io_out_c_data;
  wire                pe_mat_8_24_io_out_c_is_weight;
  wire       [15:0]   pe_mat_8_25_io_out_r_data;
  wire                pe_mat_8_25_io_out_r_stop_weight;
  wire                pe_mat_8_25_io_out_r_stall;
  wire       [15:0]   pe_mat_8_25_io_out_c_data;
  wire                pe_mat_8_25_io_out_c_is_weight;
  wire       [15:0]   pe_mat_8_26_io_out_r_data;
  wire                pe_mat_8_26_io_out_r_stop_weight;
  wire                pe_mat_8_26_io_out_r_stall;
  wire       [15:0]   pe_mat_8_26_io_out_c_data;
  wire                pe_mat_8_26_io_out_c_is_weight;
  wire       [15:0]   pe_mat_8_27_io_out_r_data;
  wire                pe_mat_8_27_io_out_r_stop_weight;
  wire                pe_mat_8_27_io_out_r_stall;
  wire       [15:0]   pe_mat_8_27_io_out_c_data;
  wire                pe_mat_8_27_io_out_c_is_weight;
  wire       [15:0]   pe_mat_8_28_io_out_r_data;
  wire                pe_mat_8_28_io_out_r_stop_weight;
  wire                pe_mat_8_28_io_out_r_stall;
  wire       [15:0]   pe_mat_8_28_io_out_c_data;
  wire                pe_mat_8_28_io_out_c_is_weight;
  wire       [15:0]   pe_mat_8_29_io_out_r_data;
  wire                pe_mat_8_29_io_out_r_stop_weight;
  wire                pe_mat_8_29_io_out_r_stall;
  wire       [15:0]   pe_mat_8_29_io_out_c_data;
  wire                pe_mat_8_29_io_out_c_is_weight;
  wire       [15:0]   pe_mat_8_30_io_out_r_data;
  wire                pe_mat_8_30_io_out_r_stop_weight;
  wire                pe_mat_8_30_io_out_r_stall;
  wire       [15:0]   pe_mat_8_30_io_out_c_data;
  wire                pe_mat_8_30_io_out_c_is_weight;
  wire       [15:0]   pe_mat_8_31_io_out_r_data;
  wire                pe_mat_8_31_io_out_r_stop_weight;
  wire                pe_mat_8_31_io_out_r_stall;
  wire       [15:0]   pe_mat_8_31_io_out_c_data;
  wire                pe_mat_8_31_io_out_c_is_weight;
  wire       [15:0]   pe_mat_9_0_io_out_r_data;
  wire                pe_mat_9_0_io_out_r_stop_weight;
  wire                pe_mat_9_0_io_out_r_stall;
  wire       [15:0]   pe_mat_9_0_io_out_c_data;
  wire                pe_mat_9_0_io_out_c_is_weight;
  wire       [15:0]   pe_mat_9_1_io_out_r_data;
  wire                pe_mat_9_1_io_out_r_stop_weight;
  wire                pe_mat_9_1_io_out_r_stall;
  wire       [15:0]   pe_mat_9_1_io_out_c_data;
  wire                pe_mat_9_1_io_out_c_is_weight;
  wire       [15:0]   pe_mat_9_2_io_out_r_data;
  wire                pe_mat_9_2_io_out_r_stop_weight;
  wire                pe_mat_9_2_io_out_r_stall;
  wire       [15:0]   pe_mat_9_2_io_out_c_data;
  wire                pe_mat_9_2_io_out_c_is_weight;
  wire       [15:0]   pe_mat_9_3_io_out_r_data;
  wire                pe_mat_9_3_io_out_r_stop_weight;
  wire                pe_mat_9_3_io_out_r_stall;
  wire       [15:0]   pe_mat_9_3_io_out_c_data;
  wire                pe_mat_9_3_io_out_c_is_weight;
  wire       [15:0]   pe_mat_9_4_io_out_r_data;
  wire                pe_mat_9_4_io_out_r_stop_weight;
  wire                pe_mat_9_4_io_out_r_stall;
  wire       [15:0]   pe_mat_9_4_io_out_c_data;
  wire                pe_mat_9_4_io_out_c_is_weight;
  wire       [15:0]   pe_mat_9_5_io_out_r_data;
  wire                pe_mat_9_5_io_out_r_stop_weight;
  wire                pe_mat_9_5_io_out_r_stall;
  wire       [15:0]   pe_mat_9_5_io_out_c_data;
  wire                pe_mat_9_5_io_out_c_is_weight;
  wire       [15:0]   pe_mat_9_6_io_out_r_data;
  wire                pe_mat_9_6_io_out_r_stop_weight;
  wire                pe_mat_9_6_io_out_r_stall;
  wire       [15:0]   pe_mat_9_6_io_out_c_data;
  wire                pe_mat_9_6_io_out_c_is_weight;
  wire       [15:0]   pe_mat_9_7_io_out_r_data;
  wire                pe_mat_9_7_io_out_r_stop_weight;
  wire                pe_mat_9_7_io_out_r_stall;
  wire       [15:0]   pe_mat_9_7_io_out_c_data;
  wire                pe_mat_9_7_io_out_c_is_weight;
  wire       [15:0]   pe_mat_9_8_io_out_r_data;
  wire                pe_mat_9_8_io_out_r_stop_weight;
  wire                pe_mat_9_8_io_out_r_stall;
  wire       [15:0]   pe_mat_9_8_io_out_c_data;
  wire                pe_mat_9_8_io_out_c_is_weight;
  wire       [15:0]   pe_mat_9_9_io_out_r_data;
  wire                pe_mat_9_9_io_out_r_stop_weight;
  wire                pe_mat_9_9_io_out_r_stall;
  wire       [15:0]   pe_mat_9_9_io_out_c_data;
  wire                pe_mat_9_9_io_out_c_is_weight;
  wire       [15:0]   pe_mat_9_10_io_out_r_data;
  wire                pe_mat_9_10_io_out_r_stop_weight;
  wire                pe_mat_9_10_io_out_r_stall;
  wire       [15:0]   pe_mat_9_10_io_out_c_data;
  wire                pe_mat_9_10_io_out_c_is_weight;
  wire       [15:0]   pe_mat_9_11_io_out_r_data;
  wire                pe_mat_9_11_io_out_r_stop_weight;
  wire                pe_mat_9_11_io_out_r_stall;
  wire       [15:0]   pe_mat_9_11_io_out_c_data;
  wire                pe_mat_9_11_io_out_c_is_weight;
  wire       [15:0]   pe_mat_9_12_io_out_r_data;
  wire                pe_mat_9_12_io_out_r_stop_weight;
  wire                pe_mat_9_12_io_out_r_stall;
  wire       [15:0]   pe_mat_9_12_io_out_c_data;
  wire                pe_mat_9_12_io_out_c_is_weight;
  wire       [15:0]   pe_mat_9_13_io_out_r_data;
  wire                pe_mat_9_13_io_out_r_stop_weight;
  wire                pe_mat_9_13_io_out_r_stall;
  wire       [15:0]   pe_mat_9_13_io_out_c_data;
  wire                pe_mat_9_13_io_out_c_is_weight;
  wire       [15:0]   pe_mat_9_14_io_out_r_data;
  wire                pe_mat_9_14_io_out_r_stop_weight;
  wire                pe_mat_9_14_io_out_r_stall;
  wire       [15:0]   pe_mat_9_14_io_out_c_data;
  wire                pe_mat_9_14_io_out_c_is_weight;
  wire       [15:0]   pe_mat_9_15_io_out_r_data;
  wire                pe_mat_9_15_io_out_r_stop_weight;
  wire                pe_mat_9_15_io_out_r_stall;
  wire       [15:0]   pe_mat_9_15_io_out_c_data;
  wire                pe_mat_9_15_io_out_c_is_weight;
  wire       [15:0]   pe_mat_9_16_io_out_r_data;
  wire                pe_mat_9_16_io_out_r_stop_weight;
  wire                pe_mat_9_16_io_out_r_stall;
  wire       [15:0]   pe_mat_9_16_io_out_c_data;
  wire                pe_mat_9_16_io_out_c_is_weight;
  wire       [15:0]   pe_mat_9_17_io_out_r_data;
  wire                pe_mat_9_17_io_out_r_stop_weight;
  wire                pe_mat_9_17_io_out_r_stall;
  wire       [15:0]   pe_mat_9_17_io_out_c_data;
  wire                pe_mat_9_17_io_out_c_is_weight;
  wire       [15:0]   pe_mat_9_18_io_out_r_data;
  wire                pe_mat_9_18_io_out_r_stop_weight;
  wire                pe_mat_9_18_io_out_r_stall;
  wire       [15:0]   pe_mat_9_18_io_out_c_data;
  wire                pe_mat_9_18_io_out_c_is_weight;
  wire       [15:0]   pe_mat_9_19_io_out_r_data;
  wire                pe_mat_9_19_io_out_r_stop_weight;
  wire                pe_mat_9_19_io_out_r_stall;
  wire       [15:0]   pe_mat_9_19_io_out_c_data;
  wire                pe_mat_9_19_io_out_c_is_weight;
  wire       [15:0]   pe_mat_9_20_io_out_r_data;
  wire                pe_mat_9_20_io_out_r_stop_weight;
  wire                pe_mat_9_20_io_out_r_stall;
  wire       [15:0]   pe_mat_9_20_io_out_c_data;
  wire                pe_mat_9_20_io_out_c_is_weight;
  wire       [15:0]   pe_mat_9_21_io_out_r_data;
  wire                pe_mat_9_21_io_out_r_stop_weight;
  wire                pe_mat_9_21_io_out_r_stall;
  wire       [15:0]   pe_mat_9_21_io_out_c_data;
  wire                pe_mat_9_21_io_out_c_is_weight;
  wire       [15:0]   pe_mat_9_22_io_out_r_data;
  wire                pe_mat_9_22_io_out_r_stop_weight;
  wire                pe_mat_9_22_io_out_r_stall;
  wire       [15:0]   pe_mat_9_22_io_out_c_data;
  wire                pe_mat_9_22_io_out_c_is_weight;
  wire       [15:0]   pe_mat_9_23_io_out_r_data;
  wire                pe_mat_9_23_io_out_r_stop_weight;
  wire                pe_mat_9_23_io_out_r_stall;
  wire       [15:0]   pe_mat_9_23_io_out_c_data;
  wire                pe_mat_9_23_io_out_c_is_weight;
  wire       [15:0]   pe_mat_9_24_io_out_r_data;
  wire                pe_mat_9_24_io_out_r_stop_weight;
  wire                pe_mat_9_24_io_out_r_stall;
  wire       [15:0]   pe_mat_9_24_io_out_c_data;
  wire                pe_mat_9_24_io_out_c_is_weight;
  wire       [15:0]   pe_mat_9_25_io_out_r_data;
  wire                pe_mat_9_25_io_out_r_stop_weight;
  wire                pe_mat_9_25_io_out_r_stall;
  wire       [15:0]   pe_mat_9_25_io_out_c_data;
  wire                pe_mat_9_25_io_out_c_is_weight;
  wire       [15:0]   pe_mat_9_26_io_out_r_data;
  wire                pe_mat_9_26_io_out_r_stop_weight;
  wire                pe_mat_9_26_io_out_r_stall;
  wire       [15:0]   pe_mat_9_26_io_out_c_data;
  wire                pe_mat_9_26_io_out_c_is_weight;
  wire       [15:0]   pe_mat_9_27_io_out_r_data;
  wire                pe_mat_9_27_io_out_r_stop_weight;
  wire                pe_mat_9_27_io_out_r_stall;
  wire       [15:0]   pe_mat_9_27_io_out_c_data;
  wire                pe_mat_9_27_io_out_c_is_weight;
  wire       [15:0]   pe_mat_9_28_io_out_r_data;
  wire                pe_mat_9_28_io_out_r_stop_weight;
  wire                pe_mat_9_28_io_out_r_stall;
  wire       [15:0]   pe_mat_9_28_io_out_c_data;
  wire                pe_mat_9_28_io_out_c_is_weight;
  wire       [15:0]   pe_mat_9_29_io_out_r_data;
  wire                pe_mat_9_29_io_out_r_stop_weight;
  wire                pe_mat_9_29_io_out_r_stall;
  wire       [15:0]   pe_mat_9_29_io_out_c_data;
  wire                pe_mat_9_29_io_out_c_is_weight;
  wire       [15:0]   pe_mat_9_30_io_out_r_data;
  wire                pe_mat_9_30_io_out_r_stop_weight;
  wire                pe_mat_9_30_io_out_r_stall;
  wire       [15:0]   pe_mat_9_30_io_out_c_data;
  wire                pe_mat_9_30_io_out_c_is_weight;
  wire       [15:0]   pe_mat_9_31_io_out_r_data;
  wire                pe_mat_9_31_io_out_r_stop_weight;
  wire                pe_mat_9_31_io_out_r_stall;
  wire       [15:0]   pe_mat_9_31_io_out_c_data;
  wire                pe_mat_9_31_io_out_c_is_weight;
  wire       [15:0]   pe_mat_10_0_io_out_r_data;
  wire                pe_mat_10_0_io_out_r_stop_weight;
  wire                pe_mat_10_0_io_out_r_stall;
  wire       [15:0]   pe_mat_10_0_io_out_c_data;
  wire                pe_mat_10_0_io_out_c_is_weight;
  wire       [15:0]   pe_mat_10_1_io_out_r_data;
  wire                pe_mat_10_1_io_out_r_stop_weight;
  wire                pe_mat_10_1_io_out_r_stall;
  wire       [15:0]   pe_mat_10_1_io_out_c_data;
  wire                pe_mat_10_1_io_out_c_is_weight;
  wire       [15:0]   pe_mat_10_2_io_out_r_data;
  wire                pe_mat_10_2_io_out_r_stop_weight;
  wire                pe_mat_10_2_io_out_r_stall;
  wire       [15:0]   pe_mat_10_2_io_out_c_data;
  wire                pe_mat_10_2_io_out_c_is_weight;
  wire       [15:0]   pe_mat_10_3_io_out_r_data;
  wire                pe_mat_10_3_io_out_r_stop_weight;
  wire                pe_mat_10_3_io_out_r_stall;
  wire       [15:0]   pe_mat_10_3_io_out_c_data;
  wire                pe_mat_10_3_io_out_c_is_weight;
  wire       [15:0]   pe_mat_10_4_io_out_r_data;
  wire                pe_mat_10_4_io_out_r_stop_weight;
  wire                pe_mat_10_4_io_out_r_stall;
  wire       [15:0]   pe_mat_10_4_io_out_c_data;
  wire                pe_mat_10_4_io_out_c_is_weight;
  wire       [15:0]   pe_mat_10_5_io_out_r_data;
  wire                pe_mat_10_5_io_out_r_stop_weight;
  wire                pe_mat_10_5_io_out_r_stall;
  wire       [15:0]   pe_mat_10_5_io_out_c_data;
  wire                pe_mat_10_5_io_out_c_is_weight;
  wire       [15:0]   pe_mat_10_6_io_out_r_data;
  wire                pe_mat_10_6_io_out_r_stop_weight;
  wire                pe_mat_10_6_io_out_r_stall;
  wire       [15:0]   pe_mat_10_6_io_out_c_data;
  wire                pe_mat_10_6_io_out_c_is_weight;
  wire       [15:0]   pe_mat_10_7_io_out_r_data;
  wire                pe_mat_10_7_io_out_r_stop_weight;
  wire                pe_mat_10_7_io_out_r_stall;
  wire       [15:0]   pe_mat_10_7_io_out_c_data;
  wire                pe_mat_10_7_io_out_c_is_weight;
  wire       [15:0]   pe_mat_10_8_io_out_r_data;
  wire                pe_mat_10_8_io_out_r_stop_weight;
  wire                pe_mat_10_8_io_out_r_stall;
  wire       [15:0]   pe_mat_10_8_io_out_c_data;
  wire                pe_mat_10_8_io_out_c_is_weight;
  wire       [15:0]   pe_mat_10_9_io_out_r_data;
  wire                pe_mat_10_9_io_out_r_stop_weight;
  wire                pe_mat_10_9_io_out_r_stall;
  wire       [15:0]   pe_mat_10_9_io_out_c_data;
  wire                pe_mat_10_9_io_out_c_is_weight;
  wire       [15:0]   pe_mat_10_10_io_out_r_data;
  wire                pe_mat_10_10_io_out_r_stop_weight;
  wire                pe_mat_10_10_io_out_r_stall;
  wire       [15:0]   pe_mat_10_10_io_out_c_data;
  wire                pe_mat_10_10_io_out_c_is_weight;
  wire       [15:0]   pe_mat_10_11_io_out_r_data;
  wire                pe_mat_10_11_io_out_r_stop_weight;
  wire                pe_mat_10_11_io_out_r_stall;
  wire       [15:0]   pe_mat_10_11_io_out_c_data;
  wire                pe_mat_10_11_io_out_c_is_weight;
  wire       [15:0]   pe_mat_10_12_io_out_r_data;
  wire                pe_mat_10_12_io_out_r_stop_weight;
  wire                pe_mat_10_12_io_out_r_stall;
  wire       [15:0]   pe_mat_10_12_io_out_c_data;
  wire                pe_mat_10_12_io_out_c_is_weight;
  wire       [15:0]   pe_mat_10_13_io_out_r_data;
  wire                pe_mat_10_13_io_out_r_stop_weight;
  wire                pe_mat_10_13_io_out_r_stall;
  wire       [15:0]   pe_mat_10_13_io_out_c_data;
  wire                pe_mat_10_13_io_out_c_is_weight;
  wire       [15:0]   pe_mat_10_14_io_out_r_data;
  wire                pe_mat_10_14_io_out_r_stop_weight;
  wire                pe_mat_10_14_io_out_r_stall;
  wire       [15:0]   pe_mat_10_14_io_out_c_data;
  wire                pe_mat_10_14_io_out_c_is_weight;
  wire       [15:0]   pe_mat_10_15_io_out_r_data;
  wire                pe_mat_10_15_io_out_r_stop_weight;
  wire                pe_mat_10_15_io_out_r_stall;
  wire       [15:0]   pe_mat_10_15_io_out_c_data;
  wire                pe_mat_10_15_io_out_c_is_weight;
  wire       [15:0]   pe_mat_10_16_io_out_r_data;
  wire                pe_mat_10_16_io_out_r_stop_weight;
  wire                pe_mat_10_16_io_out_r_stall;
  wire       [15:0]   pe_mat_10_16_io_out_c_data;
  wire                pe_mat_10_16_io_out_c_is_weight;
  wire       [15:0]   pe_mat_10_17_io_out_r_data;
  wire                pe_mat_10_17_io_out_r_stop_weight;
  wire                pe_mat_10_17_io_out_r_stall;
  wire       [15:0]   pe_mat_10_17_io_out_c_data;
  wire                pe_mat_10_17_io_out_c_is_weight;
  wire       [15:0]   pe_mat_10_18_io_out_r_data;
  wire                pe_mat_10_18_io_out_r_stop_weight;
  wire                pe_mat_10_18_io_out_r_stall;
  wire       [15:0]   pe_mat_10_18_io_out_c_data;
  wire                pe_mat_10_18_io_out_c_is_weight;
  wire       [15:0]   pe_mat_10_19_io_out_r_data;
  wire                pe_mat_10_19_io_out_r_stop_weight;
  wire                pe_mat_10_19_io_out_r_stall;
  wire       [15:0]   pe_mat_10_19_io_out_c_data;
  wire                pe_mat_10_19_io_out_c_is_weight;
  wire       [15:0]   pe_mat_10_20_io_out_r_data;
  wire                pe_mat_10_20_io_out_r_stop_weight;
  wire                pe_mat_10_20_io_out_r_stall;
  wire       [15:0]   pe_mat_10_20_io_out_c_data;
  wire                pe_mat_10_20_io_out_c_is_weight;
  wire       [15:0]   pe_mat_10_21_io_out_r_data;
  wire                pe_mat_10_21_io_out_r_stop_weight;
  wire                pe_mat_10_21_io_out_r_stall;
  wire       [15:0]   pe_mat_10_21_io_out_c_data;
  wire                pe_mat_10_21_io_out_c_is_weight;
  wire       [15:0]   pe_mat_10_22_io_out_r_data;
  wire                pe_mat_10_22_io_out_r_stop_weight;
  wire                pe_mat_10_22_io_out_r_stall;
  wire       [15:0]   pe_mat_10_22_io_out_c_data;
  wire                pe_mat_10_22_io_out_c_is_weight;
  wire       [15:0]   pe_mat_10_23_io_out_r_data;
  wire                pe_mat_10_23_io_out_r_stop_weight;
  wire                pe_mat_10_23_io_out_r_stall;
  wire       [15:0]   pe_mat_10_23_io_out_c_data;
  wire                pe_mat_10_23_io_out_c_is_weight;
  wire       [15:0]   pe_mat_10_24_io_out_r_data;
  wire                pe_mat_10_24_io_out_r_stop_weight;
  wire                pe_mat_10_24_io_out_r_stall;
  wire       [15:0]   pe_mat_10_24_io_out_c_data;
  wire                pe_mat_10_24_io_out_c_is_weight;
  wire       [15:0]   pe_mat_10_25_io_out_r_data;
  wire                pe_mat_10_25_io_out_r_stop_weight;
  wire                pe_mat_10_25_io_out_r_stall;
  wire       [15:0]   pe_mat_10_25_io_out_c_data;
  wire                pe_mat_10_25_io_out_c_is_weight;
  wire       [15:0]   pe_mat_10_26_io_out_r_data;
  wire                pe_mat_10_26_io_out_r_stop_weight;
  wire                pe_mat_10_26_io_out_r_stall;
  wire       [15:0]   pe_mat_10_26_io_out_c_data;
  wire                pe_mat_10_26_io_out_c_is_weight;
  wire       [15:0]   pe_mat_10_27_io_out_r_data;
  wire                pe_mat_10_27_io_out_r_stop_weight;
  wire                pe_mat_10_27_io_out_r_stall;
  wire       [15:0]   pe_mat_10_27_io_out_c_data;
  wire                pe_mat_10_27_io_out_c_is_weight;
  wire       [15:0]   pe_mat_10_28_io_out_r_data;
  wire                pe_mat_10_28_io_out_r_stop_weight;
  wire                pe_mat_10_28_io_out_r_stall;
  wire       [15:0]   pe_mat_10_28_io_out_c_data;
  wire                pe_mat_10_28_io_out_c_is_weight;
  wire       [15:0]   pe_mat_10_29_io_out_r_data;
  wire                pe_mat_10_29_io_out_r_stop_weight;
  wire                pe_mat_10_29_io_out_r_stall;
  wire       [15:0]   pe_mat_10_29_io_out_c_data;
  wire                pe_mat_10_29_io_out_c_is_weight;
  wire       [15:0]   pe_mat_10_30_io_out_r_data;
  wire                pe_mat_10_30_io_out_r_stop_weight;
  wire                pe_mat_10_30_io_out_r_stall;
  wire       [15:0]   pe_mat_10_30_io_out_c_data;
  wire                pe_mat_10_30_io_out_c_is_weight;
  wire       [15:0]   pe_mat_10_31_io_out_r_data;
  wire                pe_mat_10_31_io_out_r_stop_weight;
  wire                pe_mat_10_31_io_out_r_stall;
  wire       [15:0]   pe_mat_10_31_io_out_c_data;
  wire                pe_mat_10_31_io_out_c_is_weight;
  wire       [15:0]   pe_mat_11_0_io_out_r_data;
  wire                pe_mat_11_0_io_out_r_stop_weight;
  wire                pe_mat_11_0_io_out_r_stall;
  wire       [15:0]   pe_mat_11_0_io_out_c_data;
  wire                pe_mat_11_0_io_out_c_is_weight;
  wire       [15:0]   pe_mat_11_1_io_out_r_data;
  wire                pe_mat_11_1_io_out_r_stop_weight;
  wire                pe_mat_11_1_io_out_r_stall;
  wire       [15:0]   pe_mat_11_1_io_out_c_data;
  wire                pe_mat_11_1_io_out_c_is_weight;
  wire       [15:0]   pe_mat_11_2_io_out_r_data;
  wire                pe_mat_11_2_io_out_r_stop_weight;
  wire                pe_mat_11_2_io_out_r_stall;
  wire       [15:0]   pe_mat_11_2_io_out_c_data;
  wire                pe_mat_11_2_io_out_c_is_weight;
  wire       [15:0]   pe_mat_11_3_io_out_r_data;
  wire                pe_mat_11_3_io_out_r_stop_weight;
  wire                pe_mat_11_3_io_out_r_stall;
  wire       [15:0]   pe_mat_11_3_io_out_c_data;
  wire                pe_mat_11_3_io_out_c_is_weight;
  wire       [15:0]   pe_mat_11_4_io_out_r_data;
  wire                pe_mat_11_4_io_out_r_stop_weight;
  wire                pe_mat_11_4_io_out_r_stall;
  wire       [15:0]   pe_mat_11_4_io_out_c_data;
  wire                pe_mat_11_4_io_out_c_is_weight;
  wire       [15:0]   pe_mat_11_5_io_out_r_data;
  wire                pe_mat_11_5_io_out_r_stop_weight;
  wire                pe_mat_11_5_io_out_r_stall;
  wire       [15:0]   pe_mat_11_5_io_out_c_data;
  wire                pe_mat_11_5_io_out_c_is_weight;
  wire       [15:0]   pe_mat_11_6_io_out_r_data;
  wire                pe_mat_11_6_io_out_r_stop_weight;
  wire                pe_mat_11_6_io_out_r_stall;
  wire       [15:0]   pe_mat_11_6_io_out_c_data;
  wire                pe_mat_11_6_io_out_c_is_weight;
  wire       [15:0]   pe_mat_11_7_io_out_r_data;
  wire                pe_mat_11_7_io_out_r_stop_weight;
  wire                pe_mat_11_7_io_out_r_stall;
  wire       [15:0]   pe_mat_11_7_io_out_c_data;
  wire                pe_mat_11_7_io_out_c_is_weight;
  wire       [15:0]   pe_mat_11_8_io_out_r_data;
  wire                pe_mat_11_8_io_out_r_stop_weight;
  wire                pe_mat_11_8_io_out_r_stall;
  wire       [15:0]   pe_mat_11_8_io_out_c_data;
  wire                pe_mat_11_8_io_out_c_is_weight;
  wire       [15:0]   pe_mat_11_9_io_out_r_data;
  wire                pe_mat_11_9_io_out_r_stop_weight;
  wire                pe_mat_11_9_io_out_r_stall;
  wire       [15:0]   pe_mat_11_9_io_out_c_data;
  wire                pe_mat_11_9_io_out_c_is_weight;
  wire       [15:0]   pe_mat_11_10_io_out_r_data;
  wire                pe_mat_11_10_io_out_r_stop_weight;
  wire                pe_mat_11_10_io_out_r_stall;
  wire       [15:0]   pe_mat_11_10_io_out_c_data;
  wire                pe_mat_11_10_io_out_c_is_weight;
  wire       [15:0]   pe_mat_11_11_io_out_r_data;
  wire                pe_mat_11_11_io_out_r_stop_weight;
  wire                pe_mat_11_11_io_out_r_stall;
  wire       [15:0]   pe_mat_11_11_io_out_c_data;
  wire                pe_mat_11_11_io_out_c_is_weight;
  wire       [15:0]   pe_mat_11_12_io_out_r_data;
  wire                pe_mat_11_12_io_out_r_stop_weight;
  wire                pe_mat_11_12_io_out_r_stall;
  wire       [15:0]   pe_mat_11_12_io_out_c_data;
  wire                pe_mat_11_12_io_out_c_is_weight;
  wire       [15:0]   pe_mat_11_13_io_out_r_data;
  wire                pe_mat_11_13_io_out_r_stop_weight;
  wire                pe_mat_11_13_io_out_r_stall;
  wire       [15:0]   pe_mat_11_13_io_out_c_data;
  wire                pe_mat_11_13_io_out_c_is_weight;
  wire       [15:0]   pe_mat_11_14_io_out_r_data;
  wire                pe_mat_11_14_io_out_r_stop_weight;
  wire                pe_mat_11_14_io_out_r_stall;
  wire       [15:0]   pe_mat_11_14_io_out_c_data;
  wire                pe_mat_11_14_io_out_c_is_weight;
  wire       [15:0]   pe_mat_11_15_io_out_r_data;
  wire                pe_mat_11_15_io_out_r_stop_weight;
  wire                pe_mat_11_15_io_out_r_stall;
  wire       [15:0]   pe_mat_11_15_io_out_c_data;
  wire                pe_mat_11_15_io_out_c_is_weight;
  wire       [15:0]   pe_mat_11_16_io_out_r_data;
  wire                pe_mat_11_16_io_out_r_stop_weight;
  wire                pe_mat_11_16_io_out_r_stall;
  wire       [15:0]   pe_mat_11_16_io_out_c_data;
  wire                pe_mat_11_16_io_out_c_is_weight;
  wire       [15:0]   pe_mat_11_17_io_out_r_data;
  wire                pe_mat_11_17_io_out_r_stop_weight;
  wire                pe_mat_11_17_io_out_r_stall;
  wire       [15:0]   pe_mat_11_17_io_out_c_data;
  wire                pe_mat_11_17_io_out_c_is_weight;
  wire       [15:0]   pe_mat_11_18_io_out_r_data;
  wire                pe_mat_11_18_io_out_r_stop_weight;
  wire                pe_mat_11_18_io_out_r_stall;
  wire       [15:0]   pe_mat_11_18_io_out_c_data;
  wire                pe_mat_11_18_io_out_c_is_weight;
  wire       [15:0]   pe_mat_11_19_io_out_r_data;
  wire                pe_mat_11_19_io_out_r_stop_weight;
  wire                pe_mat_11_19_io_out_r_stall;
  wire       [15:0]   pe_mat_11_19_io_out_c_data;
  wire                pe_mat_11_19_io_out_c_is_weight;
  wire       [15:0]   pe_mat_11_20_io_out_r_data;
  wire                pe_mat_11_20_io_out_r_stop_weight;
  wire                pe_mat_11_20_io_out_r_stall;
  wire       [15:0]   pe_mat_11_20_io_out_c_data;
  wire                pe_mat_11_20_io_out_c_is_weight;
  wire       [15:0]   pe_mat_11_21_io_out_r_data;
  wire                pe_mat_11_21_io_out_r_stop_weight;
  wire                pe_mat_11_21_io_out_r_stall;
  wire       [15:0]   pe_mat_11_21_io_out_c_data;
  wire                pe_mat_11_21_io_out_c_is_weight;
  wire       [15:0]   pe_mat_11_22_io_out_r_data;
  wire                pe_mat_11_22_io_out_r_stop_weight;
  wire                pe_mat_11_22_io_out_r_stall;
  wire       [15:0]   pe_mat_11_22_io_out_c_data;
  wire                pe_mat_11_22_io_out_c_is_weight;
  wire       [15:0]   pe_mat_11_23_io_out_r_data;
  wire                pe_mat_11_23_io_out_r_stop_weight;
  wire                pe_mat_11_23_io_out_r_stall;
  wire       [15:0]   pe_mat_11_23_io_out_c_data;
  wire                pe_mat_11_23_io_out_c_is_weight;
  wire       [15:0]   pe_mat_11_24_io_out_r_data;
  wire                pe_mat_11_24_io_out_r_stop_weight;
  wire                pe_mat_11_24_io_out_r_stall;
  wire       [15:0]   pe_mat_11_24_io_out_c_data;
  wire                pe_mat_11_24_io_out_c_is_weight;
  wire       [15:0]   pe_mat_11_25_io_out_r_data;
  wire                pe_mat_11_25_io_out_r_stop_weight;
  wire                pe_mat_11_25_io_out_r_stall;
  wire       [15:0]   pe_mat_11_25_io_out_c_data;
  wire                pe_mat_11_25_io_out_c_is_weight;
  wire       [15:0]   pe_mat_11_26_io_out_r_data;
  wire                pe_mat_11_26_io_out_r_stop_weight;
  wire                pe_mat_11_26_io_out_r_stall;
  wire       [15:0]   pe_mat_11_26_io_out_c_data;
  wire                pe_mat_11_26_io_out_c_is_weight;
  wire       [15:0]   pe_mat_11_27_io_out_r_data;
  wire                pe_mat_11_27_io_out_r_stop_weight;
  wire                pe_mat_11_27_io_out_r_stall;
  wire       [15:0]   pe_mat_11_27_io_out_c_data;
  wire                pe_mat_11_27_io_out_c_is_weight;
  wire       [15:0]   pe_mat_11_28_io_out_r_data;
  wire                pe_mat_11_28_io_out_r_stop_weight;
  wire                pe_mat_11_28_io_out_r_stall;
  wire       [15:0]   pe_mat_11_28_io_out_c_data;
  wire                pe_mat_11_28_io_out_c_is_weight;
  wire       [15:0]   pe_mat_11_29_io_out_r_data;
  wire                pe_mat_11_29_io_out_r_stop_weight;
  wire                pe_mat_11_29_io_out_r_stall;
  wire       [15:0]   pe_mat_11_29_io_out_c_data;
  wire                pe_mat_11_29_io_out_c_is_weight;
  wire       [15:0]   pe_mat_11_30_io_out_r_data;
  wire                pe_mat_11_30_io_out_r_stop_weight;
  wire                pe_mat_11_30_io_out_r_stall;
  wire       [15:0]   pe_mat_11_30_io_out_c_data;
  wire                pe_mat_11_30_io_out_c_is_weight;
  wire       [15:0]   pe_mat_11_31_io_out_r_data;
  wire                pe_mat_11_31_io_out_r_stop_weight;
  wire                pe_mat_11_31_io_out_r_stall;
  wire       [15:0]   pe_mat_11_31_io_out_c_data;
  wire                pe_mat_11_31_io_out_c_is_weight;
  wire       [15:0]   pe_mat_12_0_io_out_r_data;
  wire                pe_mat_12_0_io_out_r_stop_weight;
  wire                pe_mat_12_0_io_out_r_stall;
  wire       [15:0]   pe_mat_12_0_io_out_c_data;
  wire                pe_mat_12_0_io_out_c_is_weight;
  wire       [15:0]   pe_mat_12_1_io_out_r_data;
  wire                pe_mat_12_1_io_out_r_stop_weight;
  wire                pe_mat_12_1_io_out_r_stall;
  wire       [15:0]   pe_mat_12_1_io_out_c_data;
  wire                pe_mat_12_1_io_out_c_is_weight;
  wire       [15:0]   pe_mat_12_2_io_out_r_data;
  wire                pe_mat_12_2_io_out_r_stop_weight;
  wire                pe_mat_12_2_io_out_r_stall;
  wire       [15:0]   pe_mat_12_2_io_out_c_data;
  wire                pe_mat_12_2_io_out_c_is_weight;
  wire       [15:0]   pe_mat_12_3_io_out_r_data;
  wire                pe_mat_12_3_io_out_r_stop_weight;
  wire                pe_mat_12_3_io_out_r_stall;
  wire       [15:0]   pe_mat_12_3_io_out_c_data;
  wire                pe_mat_12_3_io_out_c_is_weight;
  wire       [15:0]   pe_mat_12_4_io_out_r_data;
  wire                pe_mat_12_4_io_out_r_stop_weight;
  wire                pe_mat_12_4_io_out_r_stall;
  wire       [15:0]   pe_mat_12_4_io_out_c_data;
  wire                pe_mat_12_4_io_out_c_is_weight;
  wire       [15:0]   pe_mat_12_5_io_out_r_data;
  wire                pe_mat_12_5_io_out_r_stop_weight;
  wire                pe_mat_12_5_io_out_r_stall;
  wire       [15:0]   pe_mat_12_5_io_out_c_data;
  wire                pe_mat_12_5_io_out_c_is_weight;
  wire       [15:0]   pe_mat_12_6_io_out_r_data;
  wire                pe_mat_12_6_io_out_r_stop_weight;
  wire                pe_mat_12_6_io_out_r_stall;
  wire       [15:0]   pe_mat_12_6_io_out_c_data;
  wire                pe_mat_12_6_io_out_c_is_weight;
  wire       [15:0]   pe_mat_12_7_io_out_r_data;
  wire                pe_mat_12_7_io_out_r_stop_weight;
  wire                pe_mat_12_7_io_out_r_stall;
  wire       [15:0]   pe_mat_12_7_io_out_c_data;
  wire                pe_mat_12_7_io_out_c_is_weight;
  wire       [15:0]   pe_mat_12_8_io_out_r_data;
  wire                pe_mat_12_8_io_out_r_stop_weight;
  wire                pe_mat_12_8_io_out_r_stall;
  wire       [15:0]   pe_mat_12_8_io_out_c_data;
  wire                pe_mat_12_8_io_out_c_is_weight;
  wire       [15:0]   pe_mat_12_9_io_out_r_data;
  wire                pe_mat_12_9_io_out_r_stop_weight;
  wire                pe_mat_12_9_io_out_r_stall;
  wire       [15:0]   pe_mat_12_9_io_out_c_data;
  wire                pe_mat_12_9_io_out_c_is_weight;
  wire       [15:0]   pe_mat_12_10_io_out_r_data;
  wire                pe_mat_12_10_io_out_r_stop_weight;
  wire                pe_mat_12_10_io_out_r_stall;
  wire       [15:0]   pe_mat_12_10_io_out_c_data;
  wire                pe_mat_12_10_io_out_c_is_weight;
  wire       [15:0]   pe_mat_12_11_io_out_r_data;
  wire                pe_mat_12_11_io_out_r_stop_weight;
  wire                pe_mat_12_11_io_out_r_stall;
  wire       [15:0]   pe_mat_12_11_io_out_c_data;
  wire                pe_mat_12_11_io_out_c_is_weight;
  wire       [15:0]   pe_mat_12_12_io_out_r_data;
  wire                pe_mat_12_12_io_out_r_stop_weight;
  wire                pe_mat_12_12_io_out_r_stall;
  wire       [15:0]   pe_mat_12_12_io_out_c_data;
  wire                pe_mat_12_12_io_out_c_is_weight;
  wire       [15:0]   pe_mat_12_13_io_out_r_data;
  wire                pe_mat_12_13_io_out_r_stop_weight;
  wire                pe_mat_12_13_io_out_r_stall;
  wire       [15:0]   pe_mat_12_13_io_out_c_data;
  wire                pe_mat_12_13_io_out_c_is_weight;
  wire       [15:0]   pe_mat_12_14_io_out_r_data;
  wire                pe_mat_12_14_io_out_r_stop_weight;
  wire                pe_mat_12_14_io_out_r_stall;
  wire       [15:0]   pe_mat_12_14_io_out_c_data;
  wire                pe_mat_12_14_io_out_c_is_weight;
  wire       [15:0]   pe_mat_12_15_io_out_r_data;
  wire                pe_mat_12_15_io_out_r_stop_weight;
  wire                pe_mat_12_15_io_out_r_stall;
  wire       [15:0]   pe_mat_12_15_io_out_c_data;
  wire                pe_mat_12_15_io_out_c_is_weight;
  wire       [15:0]   pe_mat_12_16_io_out_r_data;
  wire                pe_mat_12_16_io_out_r_stop_weight;
  wire                pe_mat_12_16_io_out_r_stall;
  wire       [15:0]   pe_mat_12_16_io_out_c_data;
  wire                pe_mat_12_16_io_out_c_is_weight;
  wire       [15:0]   pe_mat_12_17_io_out_r_data;
  wire                pe_mat_12_17_io_out_r_stop_weight;
  wire                pe_mat_12_17_io_out_r_stall;
  wire       [15:0]   pe_mat_12_17_io_out_c_data;
  wire                pe_mat_12_17_io_out_c_is_weight;
  wire       [15:0]   pe_mat_12_18_io_out_r_data;
  wire                pe_mat_12_18_io_out_r_stop_weight;
  wire                pe_mat_12_18_io_out_r_stall;
  wire       [15:0]   pe_mat_12_18_io_out_c_data;
  wire                pe_mat_12_18_io_out_c_is_weight;
  wire       [15:0]   pe_mat_12_19_io_out_r_data;
  wire                pe_mat_12_19_io_out_r_stop_weight;
  wire                pe_mat_12_19_io_out_r_stall;
  wire       [15:0]   pe_mat_12_19_io_out_c_data;
  wire                pe_mat_12_19_io_out_c_is_weight;
  wire       [15:0]   pe_mat_12_20_io_out_r_data;
  wire                pe_mat_12_20_io_out_r_stop_weight;
  wire                pe_mat_12_20_io_out_r_stall;
  wire       [15:0]   pe_mat_12_20_io_out_c_data;
  wire                pe_mat_12_20_io_out_c_is_weight;
  wire       [15:0]   pe_mat_12_21_io_out_r_data;
  wire                pe_mat_12_21_io_out_r_stop_weight;
  wire                pe_mat_12_21_io_out_r_stall;
  wire       [15:0]   pe_mat_12_21_io_out_c_data;
  wire                pe_mat_12_21_io_out_c_is_weight;
  wire       [15:0]   pe_mat_12_22_io_out_r_data;
  wire                pe_mat_12_22_io_out_r_stop_weight;
  wire                pe_mat_12_22_io_out_r_stall;
  wire       [15:0]   pe_mat_12_22_io_out_c_data;
  wire                pe_mat_12_22_io_out_c_is_weight;
  wire       [15:0]   pe_mat_12_23_io_out_r_data;
  wire                pe_mat_12_23_io_out_r_stop_weight;
  wire                pe_mat_12_23_io_out_r_stall;
  wire       [15:0]   pe_mat_12_23_io_out_c_data;
  wire                pe_mat_12_23_io_out_c_is_weight;
  wire       [15:0]   pe_mat_12_24_io_out_r_data;
  wire                pe_mat_12_24_io_out_r_stop_weight;
  wire                pe_mat_12_24_io_out_r_stall;
  wire       [15:0]   pe_mat_12_24_io_out_c_data;
  wire                pe_mat_12_24_io_out_c_is_weight;
  wire       [15:0]   pe_mat_12_25_io_out_r_data;
  wire                pe_mat_12_25_io_out_r_stop_weight;
  wire                pe_mat_12_25_io_out_r_stall;
  wire       [15:0]   pe_mat_12_25_io_out_c_data;
  wire                pe_mat_12_25_io_out_c_is_weight;
  wire       [15:0]   pe_mat_12_26_io_out_r_data;
  wire                pe_mat_12_26_io_out_r_stop_weight;
  wire                pe_mat_12_26_io_out_r_stall;
  wire       [15:0]   pe_mat_12_26_io_out_c_data;
  wire                pe_mat_12_26_io_out_c_is_weight;
  wire       [15:0]   pe_mat_12_27_io_out_r_data;
  wire                pe_mat_12_27_io_out_r_stop_weight;
  wire                pe_mat_12_27_io_out_r_stall;
  wire       [15:0]   pe_mat_12_27_io_out_c_data;
  wire                pe_mat_12_27_io_out_c_is_weight;
  wire       [15:0]   pe_mat_12_28_io_out_r_data;
  wire                pe_mat_12_28_io_out_r_stop_weight;
  wire                pe_mat_12_28_io_out_r_stall;
  wire       [15:0]   pe_mat_12_28_io_out_c_data;
  wire                pe_mat_12_28_io_out_c_is_weight;
  wire       [15:0]   pe_mat_12_29_io_out_r_data;
  wire                pe_mat_12_29_io_out_r_stop_weight;
  wire                pe_mat_12_29_io_out_r_stall;
  wire       [15:0]   pe_mat_12_29_io_out_c_data;
  wire                pe_mat_12_29_io_out_c_is_weight;
  wire       [15:0]   pe_mat_12_30_io_out_r_data;
  wire                pe_mat_12_30_io_out_r_stop_weight;
  wire                pe_mat_12_30_io_out_r_stall;
  wire       [15:0]   pe_mat_12_30_io_out_c_data;
  wire                pe_mat_12_30_io_out_c_is_weight;
  wire       [15:0]   pe_mat_12_31_io_out_r_data;
  wire                pe_mat_12_31_io_out_r_stop_weight;
  wire                pe_mat_12_31_io_out_r_stall;
  wire       [15:0]   pe_mat_12_31_io_out_c_data;
  wire                pe_mat_12_31_io_out_c_is_weight;
  wire       [15:0]   pe_mat_13_0_io_out_r_data;
  wire                pe_mat_13_0_io_out_r_stop_weight;
  wire                pe_mat_13_0_io_out_r_stall;
  wire       [15:0]   pe_mat_13_0_io_out_c_data;
  wire                pe_mat_13_0_io_out_c_is_weight;
  wire       [15:0]   pe_mat_13_1_io_out_r_data;
  wire                pe_mat_13_1_io_out_r_stop_weight;
  wire                pe_mat_13_1_io_out_r_stall;
  wire       [15:0]   pe_mat_13_1_io_out_c_data;
  wire                pe_mat_13_1_io_out_c_is_weight;
  wire       [15:0]   pe_mat_13_2_io_out_r_data;
  wire                pe_mat_13_2_io_out_r_stop_weight;
  wire                pe_mat_13_2_io_out_r_stall;
  wire       [15:0]   pe_mat_13_2_io_out_c_data;
  wire                pe_mat_13_2_io_out_c_is_weight;
  wire       [15:0]   pe_mat_13_3_io_out_r_data;
  wire                pe_mat_13_3_io_out_r_stop_weight;
  wire                pe_mat_13_3_io_out_r_stall;
  wire       [15:0]   pe_mat_13_3_io_out_c_data;
  wire                pe_mat_13_3_io_out_c_is_weight;
  wire       [15:0]   pe_mat_13_4_io_out_r_data;
  wire                pe_mat_13_4_io_out_r_stop_weight;
  wire                pe_mat_13_4_io_out_r_stall;
  wire       [15:0]   pe_mat_13_4_io_out_c_data;
  wire                pe_mat_13_4_io_out_c_is_weight;
  wire       [15:0]   pe_mat_13_5_io_out_r_data;
  wire                pe_mat_13_5_io_out_r_stop_weight;
  wire                pe_mat_13_5_io_out_r_stall;
  wire       [15:0]   pe_mat_13_5_io_out_c_data;
  wire                pe_mat_13_5_io_out_c_is_weight;
  wire       [15:0]   pe_mat_13_6_io_out_r_data;
  wire                pe_mat_13_6_io_out_r_stop_weight;
  wire                pe_mat_13_6_io_out_r_stall;
  wire       [15:0]   pe_mat_13_6_io_out_c_data;
  wire                pe_mat_13_6_io_out_c_is_weight;
  wire       [15:0]   pe_mat_13_7_io_out_r_data;
  wire                pe_mat_13_7_io_out_r_stop_weight;
  wire                pe_mat_13_7_io_out_r_stall;
  wire       [15:0]   pe_mat_13_7_io_out_c_data;
  wire                pe_mat_13_7_io_out_c_is_weight;
  wire       [15:0]   pe_mat_13_8_io_out_r_data;
  wire                pe_mat_13_8_io_out_r_stop_weight;
  wire                pe_mat_13_8_io_out_r_stall;
  wire       [15:0]   pe_mat_13_8_io_out_c_data;
  wire                pe_mat_13_8_io_out_c_is_weight;
  wire       [15:0]   pe_mat_13_9_io_out_r_data;
  wire                pe_mat_13_9_io_out_r_stop_weight;
  wire                pe_mat_13_9_io_out_r_stall;
  wire       [15:0]   pe_mat_13_9_io_out_c_data;
  wire                pe_mat_13_9_io_out_c_is_weight;
  wire       [15:0]   pe_mat_13_10_io_out_r_data;
  wire                pe_mat_13_10_io_out_r_stop_weight;
  wire                pe_mat_13_10_io_out_r_stall;
  wire       [15:0]   pe_mat_13_10_io_out_c_data;
  wire                pe_mat_13_10_io_out_c_is_weight;
  wire       [15:0]   pe_mat_13_11_io_out_r_data;
  wire                pe_mat_13_11_io_out_r_stop_weight;
  wire                pe_mat_13_11_io_out_r_stall;
  wire       [15:0]   pe_mat_13_11_io_out_c_data;
  wire                pe_mat_13_11_io_out_c_is_weight;
  wire       [15:0]   pe_mat_13_12_io_out_r_data;
  wire                pe_mat_13_12_io_out_r_stop_weight;
  wire                pe_mat_13_12_io_out_r_stall;
  wire       [15:0]   pe_mat_13_12_io_out_c_data;
  wire                pe_mat_13_12_io_out_c_is_weight;
  wire       [15:0]   pe_mat_13_13_io_out_r_data;
  wire                pe_mat_13_13_io_out_r_stop_weight;
  wire                pe_mat_13_13_io_out_r_stall;
  wire       [15:0]   pe_mat_13_13_io_out_c_data;
  wire                pe_mat_13_13_io_out_c_is_weight;
  wire       [15:0]   pe_mat_13_14_io_out_r_data;
  wire                pe_mat_13_14_io_out_r_stop_weight;
  wire                pe_mat_13_14_io_out_r_stall;
  wire       [15:0]   pe_mat_13_14_io_out_c_data;
  wire                pe_mat_13_14_io_out_c_is_weight;
  wire       [15:0]   pe_mat_13_15_io_out_r_data;
  wire                pe_mat_13_15_io_out_r_stop_weight;
  wire                pe_mat_13_15_io_out_r_stall;
  wire       [15:0]   pe_mat_13_15_io_out_c_data;
  wire                pe_mat_13_15_io_out_c_is_weight;
  wire       [15:0]   pe_mat_13_16_io_out_r_data;
  wire                pe_mat_13_16_io_out_r_stop_weight;
  wire                pe_mat_13_16_io_out_r_stall;
  wire       [15:0]   pe_mat_13_16_io_out_c_data;
  wire                pe_mat_13_16_io_out_c_is_weight;
  wire       [15:0]   pe_mat_13_17_io_out_r_data;
  wire                pe_mat_13_17_io_out_r_stop_weight;
  wire                pe_mat_13_17_io_out_r_stall;
  wire       [15:0]   pe_mat_13_17_io_out_c_data;
  wire                pe_mat_13_17_io_out_c_is_weight;
  wire       [15:0]   pe_mat_13_18_io_out_r_data;
  wire                pe_mat_13_18_io_out_r_stop_weight;
  wire                pe_mat_13_18_io_out_r_stall;
  wire       [15:0]   pe_mat_13_18_io_out_c_data;
  wire                pe_mat_13_18_io_out_c_is_weight;
  wire       [15:0]   pe_mat_13_19_io_out_r_data;
  wire                pe_mat_13_19_io_out_r_stop_weight;
  wire                pe_mat_13_19_io_out_r_stall;
  wire       [15:0]   pe_mat_13_19_io_out_c_data;
  wire                pe_mat_13_19_io_out_c_is_weight;
  wire       [15:0]   pe_mat_13_20_io_out_r_data;
  wire                pe_mat_13_20_io_out_r_stop_weight;
  wire                pe_mat_13_20_io_out_r_stall;
  wire       [15:0]   pe_mat_13_20_io_out_c_data;
  wire                pe_mat_13_20_io_out_c_is_weight;
  wire       [15:0]   pe_mat_13_21_io_out_r_data;
  wire                pe_mat_13_21_io_out_r_stop_weight;
  wire                pe_mat_13_21_io_out_r_stall;
  wire       [15:0]   pe_mat_13_21_io_out_c_data;
  wire                pe_mat_13_21_io_out_c_is_weight;
  wire       [15:0]   pe_mat_13_22_io_out_r_data;
  wire                pe_mat_13_22_io_out_r_stop_weight;
  wire                pe_mat_13_22_io_out_r_stall;
  wire       [15:0]   pe_mat_13_22_io_out_c_data;
  wire                pe_mat_13_22_io_out_c_is_weight;
  wire       [15:0]   pe_mat_13_23_io_out_r_data;
  wire                pe_mat_13_23_io_out_r_stop_weight;
  wire                pe_mat_13_23_io_out_r_stall;
  wire       [15:0]   pe_mat_13_23_io_out_c_data;
  wire                pe_mat_13_23_io_out_c_is_weight;
  wire       [15:0]   pe_mat_13_24_io_out_r_data;
  wire                pe_mat_13_24_io_out_r_stop_weight;
  wire                pe_mat_13_24_io_out_r_stall;
  wire       [15:0]   pe_mat_13_24_io_out_c_data;
  wire                pe_mat_13_24_io_out_c_is_weight;
  wire       [15:0]   pe_mat_13_25_io_out_r_data;
  wire                pe_mat_13_25_io_out_r_stop_weight;
  wire                pe_mat_13_25_io_out_r_stall;
  wire       [15:0]   pe_mat_13_25_io_out_c_data;
  wire                pe_mat_13_25_io_out_c_is_weight;
  wire       [15:0]   pe_mat_13_26_io_out_r_data;
  wire                pe_mat_13_26_io_out_r_stop_weight;
  wire                pe_mat_13_26_io_out_r_stall;
  wire       [15:0]   pe_mat_13_26_io_out_c_data;
  wire                pe_mat_13_26_io_out_c_is_weight;
  wire       [15:0]   pe_mat_13_27_io_out_r_data;
  wire                pe_mat_13_27_io_out_r_stop_weight;
  wire                pe_mat_13_27_io_out_r_stall;
  wire       [15:0]   pe_mat_13_27_io_out_c_data;
  wire                pe_mat_13_27_io_out_c_is_weight;
  wire       [15:0]   pe_mat_13_28_io_out_r_data;
  wire                pe_mat_13_28_io_out_r_stop_weight;
  wire                pe_mat_13_28_io_out_r_stall;
  wire       [15:0]   pe_mat_13_28_io_out_c_data;
  wire                pe_mat_13_28_io_out_c_is_weight;
  wire       [15:0]   pe_mat_13_29_io_out_r_data;
  wire                pe_mat_13_29_io_out_r_stop_weight;
  wire                pe_mat_13_29_io_out_r_stall;
  wire       [15:0]   pe_mat_13_29_io_out_c_data;
  wire                pe_mat_13_29_io_out_c_is_weight;
  wire       [15:0]   pe_mat_13_30_io_out_r_data;
  wire                pe_mat_13_30_io_out_r_stop_weight;
  wire                pe_mat_13_30_io_out_r_stall;
  wire       [15:0]   pe_mat_13_30_io_out_c_data;
  wire                pe_mat_13_30_io_out_c_is_weight;
  wire       [15:0]   pe_mat_13_31_io_out_r_data;
  wire                pe_mat_13_31_io_out_r_stop_weight;
  wire                pe_mat_13_31_io_out_r_stall;
  wire       [15:0]   pe_mat_13_31_io_out_c_data;
  wire                pe_mat_13_31_io_out_c_is_weight;
  wire       [15:0]   pe_mat_14_0_io_out_r_data;
  wire                pe_mat_14_0_io_out_r_stop_weight;
  wire                pe_mat_14_0_io_out_r_stall;
  wire       [15:0]   pe_mat_14_0_io_out_c_data;
  wire                pe_mat_14_0_io_out_c_is_weight;
  wire       [15:0]   pe_mat_14_1_io_out_r_data;
  wire                pe_mat_14_1_io_out_r_stop_weight;
  wire                pe_mat_14_1_io_out_r_stall;
  wire       [15:0]   pe_mat_14_1_io_out_c_data;
  wire                pe_mat_14_1_io_out_c_is_weight;
  wire       [15:0]   pe_mat_14_2_io_out_r_data;
  wire                pe_mat_14_2_io_out_r_stop_weight;
  wire                pe_mat_14_2_io_out_r_stall;
  wire       [15:0]   pe_mat_14_2_io_out_c_data;
  wire                pe_mat_14_2_io_out_c_is_weight;
  wire       [15:0]   pe_mat_14_3_io_out_r_data;
  wire                pe_mat_14_3_io_out_r_stop_weight;
  wire                pe_mat_14_3_io_out_r_stall;
  wire       [15:0]   pe_mat_14_3_io_out_c_data;
  wire                pe_mat_14_3_io_out_c_is_weight;
  wire       [15:0]   pe_mat_14_4_io_out_r_data;
  wire                pe_mat_14_4_io_out_r_stop_weight;
  wire                pe_mat_14_4_io_out_r_stall;
  wire       [15:0]   pe_mat_14_4_io_out_c_data;
  wire                pe_mat_14_4_io_out_c_is_weight;
  wire       [15:0]   pe_mat_14_5_io_out_r_data;
  wire                pe_mat_14_5_io_out_r_stop_weight;
  wire                pe_mat_14_5_io_out_r_stall;
  wire       [15:0]   pe_mat_14_5_io_out_c_data;
  wire                pe_mat_14_5_io_out_c_is_weight;
  wire       [15:0]   pe_mat_14_6_io_out_r_data;
  wire                pe_mat_14_6_io_out_r_stop_weight;
  wire                pe_mat_14_6_io_out_r_stall;
  wire       [15:0]   pe_mat_14_6_io_out_c_data;
  wire                pe_mat_14_6_io_out_c_is_weight;
  wire       [15:0]   pe_mat_14_7_io_out_r_data;
  wire                pe_mat_14_7_io_out_r_stop_weight;
  wire                pe_mat_14_7_io_out_r_stall;
  wire       [15:0]   pe_mat_14_7_io_out_c_data;
  wire                pe_mat_14_7_io_out_c_is_weight;
  wire       [15:0]   pe_mat_14_8_io_out_r_data;
  wire                pe_mat_14_8_io_out_r_stop_weight;
  wire                pe_mat_14_8_io_out_r_stall;
  wire       [15:0]   pe_mat_14_8_io_out_c_data;
  wire                pe_mat_14_8_io_out_c_is_weight;
  wire       [15:0]   pe_mat_14_9_io_out_r_data;
  wire                pe_mat_14_9_io_out_r_stop_weight;
  wire                pe_mat_14_9_io_out_r_stall;
  wire       [15:0]   pe_mat_14_9_io_out_c_data;
  wire                pe_mat_14_9_io_out_c_is_weight;
  wire       [15:0]   pe_mat_14_10_io_out_r_data;
  wire                pe_mat_14_10_io_out_r_stop_weight;
  wire                pe_mat_14_10_io_out_r_stall;
  wire       [15:0]   pe_mat_14_10_io_out_c_data;
  wire                pe_mat_14_10_io_out_c_is_weight;
  wire       [15:0]   pe_mat_14_11_io_out_r_data;
  wire                pe_mat_14_11_io_out_r_stop_weight;
  wire                pe_mat_14_11_io_out_r_stall;
  wire       [15:0]   pe_mat_14_11_io_out_c_data;
  wire                pe_mat_14_11_io_out_c_is_weight;
  wire       [15:0]   pe_mat_14_12_io_out_r_data;
  wire                pe_mat_14_12_io_out_r_stop_weight;
  wire                pe_mat_14_12_io_out_r_stall;
  wire       [15:0]   pe_mat_14_12_io_out_c_data;
  wire                pe_mat_14_12_io_out_c_is_weight;
  wire       [15:0]   pe_mat_14_13_io_out_r_data;
  wire                pe_mat_14_13_io_out_r_stop_weight;
  wire                pe_mat_14_13_io_out_r_stall;
  wire       [15:0]   pe_mat_14_13_io_out_c_data;
  wire                pe_mat_14_13_io_out_c_is_weight;
  wire       [15:0]   pe_mat_14_14_io_out_r_data;
  wire                pe_mat_14_14_io_out_r_stop_weight;
  wire                pe_mat_14_14_io_out_r_stall;
  wire       [15:0]   pe_mat_14_14_io_out_c_data;
  wire                pe_mat_14_14_io_out_c_is_weight;
  wire       [15:0]   pe_mat_14_15_io_out_r_data;
  wire                pe_mat_14_15_io_out_r_stop_weight;
  wire                pe_mat_14_15_io_out_r_stall;
  wire       [15:0]   pe_mat_14_15_io_out_c_data;
  wire                pe_mat_14_15_io_out_c_is_weight;
  wire       [15:0]   pe_mat_14_16_io_out_r_data;
  wire                pe_mat_14_16_io_out_r_stop_weight;
  wire                pe_mat_14_16_io_out_r_stall;
  wire       [15:0]   pe_mat_14_16_io_out_c_data;
  wire                pe_mat_14_16_io_out_c_is_weight;
  wire       [15:0]   pe_mat_14_17_io_out_r_data;
  wire                pe_mat_14_17_io_out_r_stop_weight;
  wire                pe_mat_14_17_io_out_r_stall;
  wire       [15:0]   pe_mat_14_17_io_out_c_data;
  wire                pe_mat_14_17_io_out_c_is_weight;
  wire       [15:0]   pe_mat_14_18_io_out_r_data;
  wire                pe_mat_14_18_io_out_r_stop_weight;
  wire                pe_mat_14_18_io_out_r_stall;
  wire       [15:0]   pe_mat_14_18_io_out_c_data;
  wire                pe_mat_14_18_io_out_c_is_weight;
  wire       [15:0]   pe_mat_14_19_io_out_r_data;
  wire                pe_mat_14_19_io_out_r_stop_weight;
  wire                pe_mat_14_19_io_out_r_stall;
  wire       [15:0]   pe_mat_14_19_io_out_c_data;
  wire                pe_mat_14_19_io_out_c_is_weight;
  wire       [15:0]   pe_mat_14_20_io_out_r_data;
  wire                pe_mat_14_20_io_out_r_stop_weight;
  wire                pe_mat_14_20_io_out_r_stall;
  wire       [15:0]   pe_mat_14_20_io_out_c_data;
  wire                pe_mat_14_20_io_out_c_is_weight;
  wire       [15:0]   pe_mat_14_21_io_out_r_data;
  wire                pe_mat_14_21_io_out_r_stop_weight;
  wire                pe_mat_14_21_io_out_r_stall;
  wire       [15:0]   pe_mat_14_21_io_out_c_data;
  wire                pe_mat_14_21_io_out_c_is_weight;
  wire       [15:0]   pe_mat_14_22_io_out_r_data;
  wire                pe_mat_14_22_io_out_r_stop_weight;
  wire                pe_mat_14_22_io_out_r_stall;
  wire       [15:0]   pe_mat_14_22_io_out_c_data;
  wire                pe_mat_14_22_io_out_c_is_weight;
  wire       [15:0]   pe_mat_14_23_io_out_r_data;
  wire                pe_mat_14_23_io_out_r_stop_weight;
  wire                pe_mat_14_23_io_out_r_stall;
  wire       [15:0]   pe_mat_14_23_io_out_c_data;
  wire                pe_mat_14_23_io_out_c_is_weight;
  wire       [15:0]   pe_mat_14_24_io_out_r_data;
  wire                pe_mat_14_24_io_out_r_stop_weight;
  wire                pe_mat_14_24_io_out_r_stall;
  wire       [15:0]   pe_mat_14_24_io_out_c_data;
  wire                pe_mat_14_24_io_out_c_is_weight;
  wire       [15:0]   pe_mat_14_25_io_out_r_data;
  wire                pe_mat_14_25_io_out_r_stop_weight;
  wire                pe_mat_14_25_io_out_r_stall;
  wire       [15:0]   pe_mat_14_25_io_out_c_data;
  wire                pe_mat_14_25_io_out_c_is_weight;
  wire       [15:0]   pe_mat_14_26_io_out_r_data;
  wire                pe_mat_14_26_io_out_r_stop_weight;
  wire                pe_mat_14_26_io_out_r_stall;
  wire       [15:0]   pe_mat_14_26_io_out_c_data;
  wire                pe_mat_14_26_io_out_c_is_weight;
  wire       [15:0]   pe_mat_14_27_io_out_r_data;
  wire                pe_mat_14_27_io_out_r_stop_weight;
  wire                pe_mat_14_27_io_out_r_stall;
  wire       [15:0]   pe_mat_14_27_io_out_c_data;
  wire                pe_mat_14_27_io_out_c_is_weight;
  wire       [15:0]   pe_mat_14_28_io_out_r_data;
  wire                pe_mat_14_28_io_out_r_stop_weight;
  wire                pe_mat_14_28_io_out_r_stall;
  wire       [15:0]   pe_mat_14_28_io_out_c_data;
  wire                pe_mat_14_28_io_out_c_is_weight;
  wire       [15:0]   pe_mat_14_29_io_out_r_data;
  wire                pe_mat_14_29_io_out_r_stop_weight;
  wire                pe_mat_14_29_io_out_r_stall;
  wire       [15:0]   pe_mat_14_29_io_out_c_data;
  wire                pe_mat_14_29_io_out_c_is_weight;
  wire       [15:0]   pe_mat_14_30_io_out_r_data;
  wire                pe_mat_14_30_io_out_r_stop_weight;
  wire                pe_mat_14_30_io_out_r_stall;
  wire       [15:0]   pe_mat_14_30_io_out_c_data;
  wire                pe_mat_14_30_io_out_c_is_weight;
  wire       [15:0]   pe_mat_14_31_io_out_r_data;
  wire                pe_mat_14_31_io_out_r_stop_weight;
  wire                pe_mat_14_31_io_out_r_stall;
  wire       [15:0]   pe_mat_14_31_io_out_c_data;
  wire                pe_mat_14_31_io_out_c_is_weight;
  wire       [15:0]   pe_mat_15_0_io_out_r_data;
  wire                pe_mat_15_0_io_out_r_stop_weight;
  wire                pe_mat_15_0_io_out_r_stall;
  wire       [15:0]   pe_mat_15_0_io_out_c_data;
  wire                pe_mat_15_0_io_out_c_is_weight;
  wire       [15:0]   pe_mat_15_1_io_out_r_data;
  wire                pe_mat_15_1_io_out_r_stop_weight;
  wire                pe_mat_15_1_io_out_r_stall;
  wire       [15:0]   pe_mat_15_1_io_out_c_data;
  wire                pe_mat_15_1_io_out_c_is_weight;
  wire       [15:0]   pe_mat_15_2_io_out_r_data;
  wire                pe_mat_15_2_io_out_r_stop_weight;
  wire                pe_mat_15_2_io_out_r_stall;
  wire       [15:0]   pe_mat_15_2_io_out_c_data;
  wire                pe_mat_15_2_io_out_c_is_weight;
  wire       [15:0]   pe_mat_15_3_io_out_r_data;
  wire                pe_mat_15_3_io_out_r_stop_weight;
  wire                pe_mat_15_3_io_out_r_stall;
  wire       [15:0]   pe_mat_15_3_io_out_c_data;
  wire                pe_mat_15_3_io_out_c_is_weight;
  wire       [15:0]   pe_mat_15_4_io_out_r_data;
  wire                pe_mat_15_4_io_out_r_stop_weight;
  wire                pe_mat_15_4_io_out_r_stall;
  wire       [15:0]   pe_mat_15_4_io_out_c_data;
  wire                pe_mat_15_4_io_out_c_is_weight;
  wire       [15:0]   pe_mat_15_5_io_out_r_data;
  wire                pe_mat_15_5_io_out_r_stop_weight;
  wire                pe_mat_15_5_io_out_r_stall;
  wire       [15:0]   pe_mat_15_5_io_out_c_data;
  wire                pe_mat_15_5_io_out_c_is_weight;
  wire       [15:0]   pe_mat_15_6_io_out_r_data;
  wire                pe_mat_15_6_io_out_r_stop_weight;
  wire                pe_mat_15_6_io_out_r_stall;
  wire       [15:0]   pe_mat_15_6_io_out_c_data;
  wire                pe_mat_15_6_io_out_c_is_weight;
  wire       [15:0]   pe_mat_15_7_io_out_r_data;
  wire                pe_mat_15_7_io_out_r_stop_weight;
  wire                pe_mat_15_7_io_out_r_stall;
  wire       [15:0]   pe_mat_15_7_io_out_c_data;
  wire                pe_mat_15_7_io_out_c_is_weight;
  wire       [15:0]   pe_mat_15_8_io_out_r_data;
  wire                pe_mat_15_8_io_out_r_stop_weight;
  wire                pe_mat_15_8_io_out_r_stall;
  wire       [15:0]   pe_mat_15_8_io_out_c_data;
  wire                pe_mat_15_8_io_out_c_is_weight;
  wire       [15:0]   pe_mat_15_9_io_out_r_data;
  wire                pe_mat_15_9_io_out_r_stop_weight;
  wire                pe_mat_15_9_io_out_r_stall;
  wire       [15:0]   pe_mat_15_9_io_out_c_data;
  wire                pe_mat_15_9_io_out_c_is_weight;
  wire       [15:0]   pe_mat_15_10_io_out_r_data;
  wire                pe_mat_15_10_io_out_r_stop_weight;
  wire                pe_mat_15_10_io_out_r_stall;
  wire       [15:0]   pe_mat_15_10_io_out_c_data;
  wire                pe_mat_15_10_io_out_c_is_weight;
  wire       [15:0]   pe_mat_15_11_io_out_r_data;
  wire                pe_mat_15_11_io_out_r_stop_weight;
  wire                pe_mat_15_11_io_out_r_stall;
  wire       [15:0]   pe_mat_15_11_io_out_c_data;
  wire                pe_mat_15_11_io_out_c_is_weight;
  wire       [15:0]   pe_mat_15_12_io_out_r_data;
  wire                pe_mat_15_12_io_out_r_stop_weight;
  wire                pe_mat_15_12_io_out_r_stall;
  wire       [15:0]   pe_mat_15_12_io_out_c_data;
  wire                pe_mat_15_12_io_out_c_is_weight;
  wire       [15:0]   pe_mat_15_13_io_out_r_data;
  wire                pe_mat_15_13_io_out_r_stop_weight;
  wire                pe_mat_15_13_io_out_r_stall;
  wire       [15:0]   pe_mat_15_13_io_out_c_data;
  wire                pe_mat_15_13_io_out_c_is_weight;
  wire       [15:0]   pe_mat_15_14_io_out_r_data;
  wire                pe_mat_15_14_io_out_r_stop_weight;
  wire                pe_mat_15_14_io_out_r_stall;
  wire       [15:0]   pe_mat_15_14_io_out_c_data;
  wire                pe_mat_15_14_io_out_c_is_weight;
  wire       [15:0]   pe_mat_15_15_io_out_r_data;
  wire                pe_mat_15_15_io_out_r_stop_weight;
  wire                pe_mat_15_15_io_out_r_stall;
  wire       [15:0]   pe_mat_15_15_io_out_c_data;
  wire                pe_mat_15_15_io_out_c_is_weight;
  wire       [15:0]   pe_mat_15_16_io_out_r_data;
  wire                pe_mat_15_16_io_out_r_stop_weight;
  wire                pe_mat_15_16_io_out_r_stall;
  wire       [15:0]   pe_mat_15_16_io_out_c_data;
  wire                pe_mat_15_16_io_out_c_is_weight;
  wire       [15:0]   pe_mat_15_17_io_out_r_data;
  wire                pe_mat_15_17_io_out_r_stop_weight;
  wire                pe_mat_15_17_io_out_r_stall;
  wire       [15:0]   pe_mat_15_17_io_out_c_data;
  wire                pe_mat_15_17_io_out_c_is_weight;
  wire       [15:0]   pe_mat_15_18_io_out_r_data;
  wire                pe_mat_15_18_io_out_r_stop_weight;
  wire                pe_mat_15_18_io_out_r_stall;
  wire       [15:0]   pe_mat_15_18_io_out_c_data;
  wire                pe_mat_15_18_io_out_c_is_weight;
  wire       [15:0]   pe_mat_15_19_io_out_r_data;
  wire                pe_mat_15_19_io_out_r_stop_weight;
  wire                pe_mat_15_19_io_out_r_stall;
  wire       [15:0]   pe_mat_15_19_io_out_c_data;
  wire                pe_mat_15_19_io_out_c_is_weight;
  wire       [15:0]   pe_mat_15_20_io_out_r_data;
  wire                pe_mat_15_20_io_out_r_stop_weight;
  wire                pe_mat_15_20_io_out_r_stall;
  wire       [15:0]   pe_mat_15_20_io_out_c_data;
  wire                pe_mat_15_20_io_out_c_is_weight;
  wire       [15:0]   pe_mat_15_21_io_out_r_data;
  wire                pe_mat_15_21_io_out_r_stop_weight;
  wire                pe_mat_15_21_io_out_r_stall;
  wire       [15:0]   pe_mat_15_21_io_out_c_data;
  wire                pe_mat_15_21_io_out_c_is_weight;
  wire       [15:0]   pe_mat_15_22_io_out_r_data;
  wire                pe_mat_15_22_io_out_r_stop_weight;
  wire                pe_mat_15_22_io_out_r_stall;
  wire       [15:0]   pe_mat_15_22_io_out_c_data;
  wire                pe_mat_15_22_io_out_c_is_weight;
  wire       [15:0]   pe_mat_15_23_io_out_r_data;
  wire                pe_mat_15_23_io_out_r_stop_weight;
  wire                pe_mat_15_23_io_out_r_stall;
  wire       [15:0]   pe_mat_15_23_io_out_c_data;
  wire                pe_mat_15_23_io_out_c_is_weight;
  wire       [15:0]   pe_mat_15_24_io_out_r_data;
  wire                pe_mat_15_24_io_out_r_stop_weight;
  wire                pe_mat_15_24_io_out_r_stall;
  wire       [15:0]   pe_mat_15_24_io_out_c_data;
  wire                pe_mat_15_24_io_out_c_is_weight;
  wire       [15:0]   pe_mat_15_25_io_out_r_data;
  wire                pe_mat_15_25_io_out_r_stop_weight;
  wire                pe_mat_15_25_io_out_r_stall;
  wire       [15:0]   pe_mat_15_25_io_out_c_data;
  wire                pe_mat_15_25_io_out_c_is_weight;
  wire       [15:0]   pe_mat_15_26_io_out_r_data;
  wire                pe_mat_15_26_io_out_r_stop_weight;
  wire                pe_mat_15_26_io_out_r_stall;
  wire       [15:0]   pe_mat_15_26_io_out_c_data;
  wire                pe_mat_15_26_io_out_c_is_weight;
  wire       [15:0]   pe_mat_15_27_io_out_r_data;
  wire                pe_mat_15_27_io_out_r_stop_weight;
  wire                pe_mat_15_27_io_out_r_stall;
  wire       [15:0]   pe_mat_15_27_io_out_c_data;
  wire                pe_mat_15_27_io_out_c_is_weight;
  wire       [15:0]   pe_mat_15_28_io_out_r_data;
  wire                pe_mat_15_28_io_out_r_stop_weight;
  wire                pe_mat_15_28_io_out_r_stall;
  wire       [15:0]   pe_mat_15_28_io_out_c_data;
  wire                pe_mat_15_28_io_out_c_is_weight;
  wire       [15:0]   pe_mat_15_29_io_out_r_data;
  wire                pe_mat_15_29_io_out_r_stop_weight;
  wire                pe_mat_15_29_io_out_r_stall;
  wire       [15:0]   pe_mat_15_29_io_out_c_data;
  wire                pe_mat_15_29_io_out_c_is_weight;
  wire       [15:0]   pe_mat_15_30_io_out_r_data;
  wire                pe_mat_15_30_io_out_r_stop_weight;
  wire                pe_mat_15_30_io_out_r_stall;
  wire       [15:0]   pe_mat_15_30_io_out_c_data;
  wire                pe_mat_15_30_io_out_c_is_weight;
  wire       [15:0]   pe_mat_15_31_io_out_r_data;
  wire                pe_mat_15_31_io_out_r_stop_weight;
  wire                pe_mat_15_31_io_out_r_stall;
  wire       [15:0]   pe_mat_15_31_io_out_c_data;
  wire                pe_mat_15_31_io_out_c_is_weight;
  wire       [15:0]   pe_mat_16_0_io_out_r_data;
  wire                pe_mat_16_0_io_out_r_stop_weight;
  wire                pe_mat_16_0_io_out_r_stall;
  wire       [15:0]   pe_mat_16_0_io_out_c_data;
  wire                pe_mat_16_0_io_out_c_is_weight;
  wire       [15:0]   pe_mat_16_1_io_out_r_data;
  wire                pe_mat_16_1_io_out_r_stop_weight;
  wire                pe_mat_16_1_io_out_r_stall;
  wire       [15:0]   pe_mat_16_1_io_out_c_data;
  wire                pe_mat_16_1_io_out_c_is_weight;
  wire       [15:0]   pe_mat_16_2_io_out_r_data;
  wire                pe_mat_16_2_io_out_r_stop_weight;
  wire                pe_mat_16_2_io_out_r_stall;
  wire       [15:0]   pe_mat_16_2_io_out_c_data;
  wire                pe_mat_16_2_io_out_c_is_weight;
  wire       [15:0]   pe_mat_16_3_io_out_r_data;
  wire                pe_mat_16_3_io_out_r_stop_weight;
  wire                pe_mat_16_3_io_out_r_stall;
  wire       [15:0]   pe_mat_16_3_io_out_c_data;
  wire                pe_mat_16_3_io_out_c_is_weight;
  wire       [15:0]   pe_mat_16_4_io_out_r_data;
  wire                pe_mat_16_4_io_out_r_stop_weight;
  wire                pe_mat_16_4_io_out_r_stall;
  wire       [15:0]   pe_mat_16_4_io_out_c_data;
  wire                pe_mat_16_4_io_out_c_is_weight;
  wire       [15:0]   pe_mat_16_5_io_out_r_data;
  wire                pe_mat_16_5_io_out_r_stop_weight;
  wire                pe_mat_16_5_io_out_r_stall;
  wire       [15:0]   pe_mat_16_5_io_out_c_data;
  wire                pe_mat_16_5_io_out_c_is_weight;
  wire       [15:0]   pe_mat_16_6_io_out_r_data;
  wire                pe_mat_16_6_io_out_r_stop_weight;
  wire                pe_mat_16_6_io_out_r_stall;
  wire       [15:0]   pe_mat_16_6_io_out_c_data;
  wire                pe_mat_16_6_io_out_c_is_weight;
  wire       [15:0]   pe_mat_16_7_io_out_r_data;
  wire                pe_mat_16_7_io_out_r_stop_weight;
  wire                pe_mat_16_7_io_out_r_stall;
  wire       [15:0]   pe_mat_16_7_io_out_c_data;
  wire                pe_mat_16_7_io_out_c_is_weight;
  wire       [15:0]   pe_mat_16_8_io_out_r_data;
  wire                pe_mat_16_8_io_out_r_stop_weight;
  wire                pe_mat_16_8_io_out_r_stall;
  wire       [15:0]   pe_mat_16_8_io_out_c_data;
  wire                pe_mat_16_8_io_out_c_is_weight;
  wire       [15:0]   pe_mat_16_9_io_out_r_data;
  wire                pe_mat_16_9_io_out_r_stop_weight;
  wire                pe_mat_16_9_io_out_r_stall;
  wire       [15:0]   pe_mat_16_9_io_out_c_data;
  wire                pe_mat_16_9_io_out_c_is_weight;
  wire       [15:0]   pe_mat_16_10_io_out_r_data;
  wire                pe_mat_16_10_io_out_r_stop_weight;
  wire                pe_mat_16_10_io_out_r_stall;
  wire       [15:0]   pe_mat_16_10_io_out_c_data;
  wire                pe_mat_16_10_io_out_c_is_weight;
  wire       [15:0]   pe_mat_16_11_io_out_r_data;
  wire                pe_mat_16_11_io_out_r_stop_weight;
  wire                pe_mat_16_11_io_out_r_stall;
  wire       [15:0]   pe_mat_16_11_io_out_c_data;
  wire                pe_mat_16_11_io_out_c_is_weight;
  wire       [15:0]   pe_mat_16_12_io_out_r_data;
  wire                pe_mat_16_12_io_out_r_stop_weight;
  wire                pe_mat_16_12_io_out_r_stall;
  wire       [15:0]   pe_mat_16_12_io_out_c_data;
  wire                pe_mat_16_12_io_out_c_is_weight;
  wire       [15:0]   pe_mat_16_13_io_out_r_data;
  wire                pe_mat_16_13_io_out_r_stop_weight;
  wire                pe_mat_16_13_io_out_r_stall;
  wire       [15:0]   pe_mat_16_13_io_out_c_data;
  wire                pe_mat_16_13_io_out_c_is_weight;
  wire       [15:0]   pe_mat_16_14_io_out_r_data;
  wire                pe_mat_16_14_io_out_r_stop_weight;
  wire                pe_mat_16_14_io_out_r_stall;
  wire       [15:0]   pe_mat_16_14_io_out_c_data;
  wire                pe_mat_16_14_io_out_c_is_weight;
  wire       [15:0]   pe_mat_16_15_io_out_r_data;
  wire                pe_mat_16_15_io_out_r_stop_weight;
  wire                pe_mat_16_15_io_out_r_stall;
  wire       [15:0]   pe_mat_16_15_io_out_c_data;
  wire                pe_mat_16_15_io_out_c_is_weight;
  wire       [15:0]   pe_mat_16_16_io_out_r_data;
  wire                pe_mat_16_16_io_out_r_stop_weight;
  wire                pe_mat_16_16_io_out_r_stall;
  wire       [15:0]   pe_mat_16_16_io_out_c_data;
  wire                pe_mat_16_16_io_out_c_is_weight;
  wire       [15:0]   pe_mat_16_17_io_out_r_data;
  wire                pe_mat_16_17_io_out_r_stop_weight;
  wire                pe_mat_16_17_io_out_r_stall;
  wire       [15:0]   pe_mat_16_17_io_out_c_data;
  wire                pe_mat_16_17_io_out_c_is_weight;
  wire       [15:0]   pe_mat_16_18_io_out_r_data;
  wire                pe_mat_16_18_io_out_r_stop_weight;
  wire                pe_mat_16_18_io_out_r_stall;
  wire       [15:0]   pe_mat_16_18_io_out_c_data;
  wire                pe_mat_16_18_io_out_c_is_weight;
  wire       [15:0]   pe_mat_16_19_io_out_r_data;
  wire                pe_mat_16_19_io_out_r_stop_weight;
  wire                pe_mat_16_19_io_out_r_stall;
  wire       [15:0]   pe_mat_16_19_io_out_c_data;
  wire                pe_mat_16_19_io_out_c_is_weight;
  wire       [15:0]   pe_mat_16_20_io_out_r_data;
  wire                pe_mat_16_20_io_out_r_stop_weight;
  wire                pe_mat_16_20_io_out_r_stall;
  wire       [15:0]   pe_mat_16_20_io_out_c_data;
  wire                pe_mat_16_20_io_out_c_is_weight;
  wire       [15:0]   pe_mat_16_21_io_out_r_data;
  wire                pe_mat_16_21_io_out_r_stop_weight;
  wire                pe_mat_16_21_io_out_r_stall;
  wire       [15:0]   pe_mat_16_21_io_out_c_data;
  wire                pe_mat_16_21_io_out_c_is_weight;
  wire       [15:0]   pe_mat_16_22_io_out_r_data;
  wire                pe_mat_16_22_io_out_r_stop_weight;
  wire                pe_mat_16_22_io_out_r_stall;
  wire       [15:0]   pe_mat_16_22_io_out_c_data;
  wire                pe_mat_16_22_io_out_c_is_weight;
  wire       [15:0]   pe_mat_16_23_io_out_r_data;
  wire                pe_mat_16_23_io_out_r_stop_weight;
  wire                pe_mat_16_23_io_out_r_stall;
  wire       [15:0]   pe_mat_16_23_io_out_c_data;
  wire                pe_mat_16_23_io_out_c_is_weight;
  wire       [15:0]   pe_mat_16_24_io_out_r_data;
  wire                pe_mat_16_24_io_out_r_stop_weight;
  wire                pe_mat_16_24_io_out_r_stall;
  wire       [15:0]   pe_mat_16_24_io_out_c_data;
  wire                pe_mat_16_24_io_out_c_is_weight;
  wire       [15:0]   pe_mat_16_25_io_out_r_data;
  wire                pe_mat_16_25_io_out_r_stop_weight;
  wire                pe_mat_16_25_io_out_r_stall;
  wire       [15:0]   pe_mat_16_25_io_out_c_data;
  wire                pe_mat_16_25_io_out_c_is_weight;
  wire       [15:0]   pe_mat_16_26_io_out_r_data;
  wire                pe_mat_16_26_io_out_r_stop_weight;
  wire                pe_mat_16_26_io_out_r_stall;
  wire       [15:0]   pe_mat_16_26_io_out_c_data;
  wire                pe_mat_16_26_io_out_c_is_weight;
  wire       [15:0]   pe_mat_16_27_io_out_r_data;
  wire                pe_mat_16_27_io_out_r_stop_weight;
  wire                pe_mat_16_27_io_out_r_stall;
  wire       [15:0]   pe_mat_16_27_io_out_c_data;
  wire                pe_mat_16_27_io_out_c_is_weight;
  wire       [15:0]   pe_mat_16_28_io_out_r_data;
  wire                pe_mat_16_28_io_out_r_stop_weight;
  wire                pe_mat_16_28_io_out_r_stall;
  wire       [15:0]   pe_mat_16_28_io_out_c_data;
  wire                pe_mat_16_28_io_out_c_is_weight;
  wire       [15:0]   pe_mat_16_29_io_out_r_data;
  wire                pe_mat_16_29_io_out_r_stop_weight;
  wire                pe_mat_16_29_io_out_r_stall;
  wire       [15:0]   pe_mat_16_29_io_out_c_data;
  wire                pe_mat_16_29_io_out_c_is_weight;
  wire       [15:0]   pe_mat_16_30_io_out_r_data;
  wire                pe_mat_16_30_io_out_r_stop_weight;
  wire                pe_mat_16_30_io_out_r_stall;
  wire       [15:0]   pe_mat_16_30_io_out_c_data;
  wire                pe_mat_16_30_io_out_c_is_weight;
  wire       [15:0]   pe_mat_16_31_io_out_r_data;
  wire                pe_mat_16_31_io_out_r_stop_weight;
  wire                pe_mat_16_31_io_out_r_stall;
  wire       [15:0]   pe_mat_16_31_io_out_c_data;
  wire                pe_mat_16_31_io_out_c_is_weight;
  wire       [15:0]   pe_mat_17_0_io_out_r_data;
  wire                pe_mat_17_0_io_out_r_stop_weight;
  wire                pe_mat_17_0_io_out_r_stall;
  wire       [15:0]   pe_mat_17_0_io_out_c_data;
  wire                pe_mat_17_0_io_out_c_is_weight;
  wire       [15:0]   pe_mat_17_1_io_out_r_data;
  wire                pe_mat_17_1_io_out_r_stop_weight;
  wire                pe_mat_17_1_io_out_r_stall;
  wire       [15:0]   pe_mat_17_1_io_out_c_data;
  wire                pe_mat_17_1_io_out_c_is_weight;
  wire       [15:0]   pe_mat_17_2_io_out_r_data;
  wire                pe_mat_17_2_io_out_r_stop_weight;
  wire                pe_mat_17_2_io_out_r_stall;
  wire       [15:0]   pe_mat_17_2_io_out_c_data;
  wire                pe_mat_17_2_io_out_c_is_weight;
  wire       [15:0]   pe_mat_17_3_io_out_r_data;
  wire                pe_mat_17_3_io_out_r_stop_weight;
  wire                pe_mat_17_3_io_out_r_stall;
  wire       [15:0]   pe_mat_17_3_io_out_c_data;
  wire                pe_mat_17_3_io_out_c_is_weight;
  wire       [15:0]   pe_mat_17_4_io_out_r_data;
  wire                pe_mat_17_4_io_out_r_stop_weight;
  wire                pe_mat_17_4_io_out_r_stall;
  wire       [15:0]   pe_mat_17_4_io_out_c_data;
  wire                pe_mat_17_4_io_out_c_is_weight;
  wire       [15:0]   pe_mat_17_5_io_out_r_data;
  wire                pe_mat_17_5_io_out_r_stop_weight;
  wire                pe_mat_17_5_io_out_r_stall;
  wire       [15:0]   pe_mat_17_5_io_out_c_data;
  wire                pe_mat_17_5_io_out_c_is_weight;
  wire       [15:0]   pe_mat_17_6_io_out_r_data;
  wire                pe_mat_17_6_io_out_r_stop_weight;
  wire                pe_mat_17_6_io_out_r_stall;
  wire       [15:0]   pe_mat_17_6_io_out_c_data;
  wire                pe_mat_17_6_io_out_c_is_weight;
  wire       [15:0]   pe_mat_17_7_io_out_r_data;
  wire                pe_mat_17_7_io_out_r_stop_weight;
  wire                pe_mat_17_7_io_out_r_stall;
  wire       [15:0]   pe_mat_17_7_io_out_c_data;
  wire                pe_mat_17_7_io_out_c_is_weight;
  wire       [15:0]   pe_mat_17_8_io_out_r_data;
  wire                pe_mat_17_8_io_out_r_stop_weight;
  wire                pe_mat_17_8_io_out_r_stall;
  wire       [15:0]   pe_mat_17_8_io_out_c_data;
  wire                pe_mat_17_8_io_out_c_is_weight;
  wire       [15:0]   pe_mat_17_9_io_out_r_data;
  wire                pe_mat_17_9_io_out_r_stop_weight;
  wire                pe_mat_17_9_io_out_r_stall;
  wire       [15:0]   pe_mat_17_9_io_out_c_data;
  wire                pe_mat_17_9_io_out_c_is_weight;
  wire       [15:0]   pe_mat_17_10_io_out_r_data;
  wire                pe_mat_17_10_io_out_r_stop_weight;
  wire                pe_mat_17_10_io_out_r_stall;
  wire       [15:0]   pe_mat_17_10_io_out_c_data;
  wire                pe_mat_17_10_io_out_c_is_weight;
  wire       [15:0]   pe_mat_17_11_io_out_r_data;
  wire                pe_mat_17_11_io_out_r_stop_weight;
  wire                pe_mat_17_11_io_out_r_stall;
  wire       [15:0]   pe_mat_17_11_io_out_c_data;
  wire                pe_mat_17_11_io_out_c_is_weight;
  wire       [15:0]   pe_mat_17_12_io_out_r_data;
  wire                pe_mat_17_12_io_out_r_stop_weight;
  wire                pe_mat_17_12_io_out_r_stall;
  wire       [15:0]   pe_mat_17_12_io_out_c_data;
  wire                pe_mat_17_12_io_out_c_is_weight;
  wire       [15:0]   pe_mat_17_13_io_out_r_data;
  wire                pe_mat_17_13_io_out_r_stop_weight;
  wire                pe_mat_17_13_io_out_r_stall;
  wire       [15:0]   pe_mat_17_13_io_out_c_data;
  wire                pe_mat_17_13_io_out_c_is_weight;
  wire       [15:0]   pe_mat_17_14_io_out_r_data;
  wire                pe_mat_17_14_io_out_r_stop_weight;
  wire                pe_mat_17_14_io_out_r_stall;
  wire       [15:0]   pe_mat_17_14_io_out_c_data;
  wire                pe_mat_17_14_io_out_c_is_weight;
  wire       [15:0]   pe_mat_17_15_io_out_r_data;
  wire                pe_mat_17_15_io_out_r_stop_weight;
  wire                pe_mat_17_15_io_out_r_stall;
  wire       [15:0]   pe_mat_17_15_io_out_c_data;
  wire                pe_mat_17_15_io_out_c_is_weight;
  wire       [15:0]   pe_mat_17_16_io_out_r_data;
  wire                pe_mat_17_16_io_out_r_stop_weight;
  wire                pe_mat_17_16_io_out_r_stall;
  wire       [15:0]   pe_mat_17_16_io_out_c_data;
  wire                pe_mat_17_16_io_out_c_is_weight;
  wire       [15:0]   pe_mat_17_17_io_out_r_data;
  wire                pe_mat_17_17_io_out_r_stop_weight;
  wire                pe_mat_17_17_io_out_r_stall;
  wire       [15:0]   pe_mat_17_17_io_out_c_data;
  wire                pe_mat_17_17_io_out_c_is_weight;
  wire       [15:0]   pe_mat_17_18_io_out_r_data;
  wire                pe_mat_17_18_io_out_r_stop_weight;
  wire                pe_mat_17_18_io_out_r_stall;
  wire       [15:0]   pe_mat_17_18_io_out_c_data;
  wire                pe_mat_17_18_io_out_c_is_weight;
  wire       [15:0]   pe_mat_17_19_io_out_r_data;
  wire                pe_mat_17_19_io_out_r_stop_weight;
  wire                pe_mat_17_19_io_out_r_stall;
  wire       [15:0]   pe_mat_17_19_io_out_c_data;
  wire                pe_mat_17_19_io_out_c_is_weight;
  wire       [15:0]   pe_mat_17_20_io_out_r_data;
  wire                pe_mat_17_20_io_out_r_stop_weight;
  wire                pe_mat_17_20_io_out_r_stall;
  wire       [15:0]   pe_mat_17_20_io_out_c_data;
  wire                pe_mat_17_20_io_out_c_is_weight;
  wire       [15:0]   pe_mat_17_21_io_out_r_data;
  wire                pe_mat_17_21_io_out_r_stop_weight;
  wire                pe_mat_17_21_io_out_r_stall;
  wire       [15:0]   pe_mat_17_21_io_out_c_data;
  wire                pe_mat_17_21_io_out_c_is_weight;
  wire       [15:0]   pe_mat_17_22_io_out_r_data;
  wire                pe_mat_17_22_io_out_r_stop_weight;
  wire                pe_mat_17_22_io_out_r_stall;
  wire       [15:0]   pe_mat_17_22_io_out_c_data;
  wire                pe_mat_17_22_io_out_c_is_weight;
  wire       [15:0]   pe_mat_17_23_io_out_r_data;
  wire                pe_mat_17_23_io_out_r_stop_weight;
  wire                pe_mat_17_23_io_out_r_stall;
  wire       [15:0]   pe_mat_17_23_io_out_c_data;
  wire                pe_mat_17_23_io_out_c_is_weight;
  wire       [15:0]   pe_mat_17_24_io_out_r_data;
  wire                pe_mat_17_24_io_out_r_stop_weight;
  wire                pe_mat_17_24_io_out_r_stall;
  wire       [15:0]   pe_mat_17_24_io_out_c_data;
  wire                pe_mat_17_24_io_out_c_is_weight;
  wire       [15:0]   pe_mat_17_25_io_out_r_data;
  wire                pe_mat_17_25_io_out_r_stop_weight;
  wire                pe_mat_17_25_io_out_r_stall;
  wire       [15:0]   pe_mat_17_25_io_out_c_data;
  wire                pe_mat_17_25_io_out_c_is_weight;
  wire       [15:0]   pe_mat_17_26_io_out_r_data;
  wire                pe_mat_17_26_io_out_r_stop_weight;
  wire                pe_mat_17_26_io_out_r_stall;
  wire       [15:0]   pe_mat_17_26_io_out_c_data;
  wire                pe_mat_17_26_io_out_c_is_weight;
  wire       [15:0]   pe_mat_17_27_io_out_r_data;
  wire                pe_mat_17_27_io_out_r_stop_weight;
  wire                pe_mat_17_27_io_out_r_stall;
  wire       [15:0]   pe_mat_17_27_io_out_c_data;
  wire                pe_mat_17_27_io_out_c_is_weight;
  wire       [15:0]   pe_mat_17_28_io_out_r_data;
  wire                pe_mat_17_28_io_out_r_stop_weight;
  wire                pe_mat_17_28_io_out_r_stall;
  wire       [15:0]   pe_mat_17_28_io_out_c_data;
  wire                pe_mat_17_28_io_out_c_is_weight;
  wire       [15:0]   pe_mat_17_29_io_out_r_data;
  wire                pe_mat_17_29_io_out_r_stop_weight;
  wire                pe_mat_17_29_io_out_r_stall;
  wire       [15:0]   pe_mat_17_29_io_out_c_data;
  wire                pe_mat_17_29_io_out_c_is_weight;
  wire       [15:0]   pe_mat_17_30_io_out_r_data;
  wire                pe_mat_17_30_io_out_r_stop_weight;
  wire                pe_mat_17_30_io_out_r_stall;
  wire       [15:0]   pe_mat_17_30_io_out_c_data;
  wire                pe_mat_17_30_io_out_c_is_weight;
  wire       [15:0]   pe_mat_17_31_io_out_r_data;
  wire                pe_mat_17_31_io_out_r_stop_weight;
  wire                pe_mat_17_31_io_out_r_stall;
  wire       [15:0]   pe_mat_17_31_io_out_c_data;
  wire                pe_mat_17_31_io_out_c_is_weight;
  wire       [15:0]   pe_mat_18_0_io_out_r_data;
  wire                pe_mat_18_0_io_out_r_stop_weight;
  wire                pe_mat_18_0_io_out_r_stall;
  wire       [15:0]   pe_mat_18_0_io_out_c_data;
  wire                pe_mat_18_0_io_out_c_is_weight;
  wire       [15:0]   pe_mat_18_1_io_out_r_data;
  wire                pe_mat_18_1_io_out_r_stop_weight;
  wire                pe_mat_18_1_io_out_r_stall;
  wire       [15:0]   pe_mat_18_1_io_out_c_data;
  wire                pe_mat_18_1_io_out_c_is_weight;
  wire       [15:0]   pe_mat_18_2_io_out_r_data;
  wire                pe_mat_18_2_io_out_r_stop_weight;
  wire                pe_mat_18_2_io_out_r_stall;
  wire       [15:0]   pe_mat_18_2_io_out_c_data;
  wire                pe_mat_18_2_io_out_c_is_weight;
  wire       [15:0]   pe_mat_18_3_io_out_r_data;
  wire                pe_mat_18_3_io_out_r_stop_weight;
  wire                pe_mat_18_3_io_out_r_stall;
  wire       [15:0]   pe_mat_18_3_io_out_c_data;
  wire                pe_mat_18_3_io_out_c_is_weight;
  wire       [15:0]   pe_mat_18_4_io_out_r_data;
  wire                pe_mat_18_4_io_out_r_stop_weight;
  wire                pe_mat_18_4_io_out_r_stall;
  wire       [15:0]   pe_mat_18_4_io_out_c_data;
  wire                pe_mat_18_4_io_out_c_is_weight;
  wire       [15:0]   pe_mat_18_5_io_out_r_data;
  wire                pe_mat_18_5_io_out_r_stop_weight;
  wire                pe_mat_18_5_io_out_r_stall;
  wire       [15:0]   pe_mat_18_5_io_out_c_data;
  wire                pe_mat_18_5_io_out_c_is_weight;
  wire       [15:0]   pe_mat_18_6_io_out_r_data;
  wire                pe_mat_18_6_io_out_r_stop_weight;
  wire                pe_mat_18_6_io_out_r_stall;
  wire       [15:0]   pe_mat_18_6_io_out_c_data;
  wire                pe_mat_18_6_io_out_c_is_weight;
  wire       [15:0]   pe_mat_18_7_io_out_r_data;
  wire                pe_mat_18_7_io_out_r_stop_weight;
  wire                pe_mat_18_7_io_out_r_stall;
  wire       [15:0]   pe_mat_18_7_io_out_c_data;
  wire                pe_mat_18_7_io_out_c_is_weight;
  wire       [15:0]   pe_mat_18_8_io_out_r_data;
  wire                pe_mat_18_8_io_out_r_stop_weight;
  wire                pe_mat_18_8_io_out_r_stall;
  wire       [15:0]   pe_mat_18_8_io_out_c_data;
  wire                pe_mat_18_8_io_out_c_is_weight;
  wire       [15:0]   pe_mat_18_9_io_out_r_data;
  wire                pe_mat_18_9_io_out_r_stop_weight;
  wire                pe_mat_18_9_io_out_r_stall;
  wire       [15:0]   pe_mat_18_9_io_out_c_data;
  wire                pe_mat_18_9_io_out_c_is_weight;
  wire       [15:0]   pe_mat_18_10_io_out_r_data;
  wire                pe_mat_18_10_io_out_r_stop_weight;
  wire                pe_mat_18_10_io_out_r_stall;
  wire       [15:0]   pe_mat_18_10_io_out_c_data;
  wire                pe_mat_18_10_io_out_c_is_weight;
  wire       [15:0]   pe_mat_18_11_io_out_r_data;
  wire                pe_mat_18_11_io_out_r_stop_weight;
  wire                pe_mat_18_11_io_out_r_stall;
  wire       [15:0]   pe_mat_18_11_io_out_c_data;
  wire                pe_mat_18_11_io_out_c_is_weight;
  wire       [15:0]   pe_mat_18_12_io_out_r_data;
  wire                pe_mat_18_12_io_out_r_stop_weight;
  wire                pe_mat_18_12_io_out_r_stall;
  wire       [15:0]   pe_mat_18_12_io_out_c_data;
  wire                pe_mat_18_12_io_out_c_is_weight;
  wire       [15:0]   pe_mat_18_13_io_out_r_data;
  wire                pe_mat_18_13_io_out_r_stop_weight;
  wire                pe_mat_18_13_io_out_r_stall;
  wire       [15:0]   pe_mat_18_13_io_out_c_data;
  wire                pe_mat_18_13_io_out_c_is_weight;
  wire       [15:0]   pe_mat_18_14_io_out_r_data;
  wire                pe_mat_18_14_io_out_r_stop_weight;
  wire                pe_mat_18_14_io_out_r_stall;
  wire       [15:0]   pe_mat_18_14_io_out_c_data;
  wire                pe_mat_18_14_io_out_c_is_weight;
  wire       [15:0]   pe_mat_18_15_io_out_r_data;
  wire                pe_mat_18_15_io_out_r_stop_weight;
  wire                pe_mat_18_15_io_out_r_stall;
  wire       [15:0]   pe_mat_18_15_io_out_c_data;
  wire                pe_mat_18_15_io_out_c_is_weight;
  wire       [15:0]   pe_mat_18_16_io_out_r_data;
  wire                pe_mat_18_16_io_out_r_stop_weight;
  wire                pe_mat_18_16_io_out_r_stall;
  wire       [15:0]   pe_mat_18_16_io_out_c_data;
  wire                pe_mat_18_16_io_out_c_is_weight;
  wire       [15:0]   pe_mat_18_17_io_out_r_data;
  wire                pe_mat_18_17_io_out_r_stop_weight;
  wire                pe_mat_18_17_io_out_r_stall;
  wire       [15:0]   pe_mat_18_17_io_out_c_data;
  wire                pe_mat_18_17_io_out_c_is_weight;
  wire       [15:0]   pe_mat_18_18_io_out_r_data;
  wire                pe_mat_18_18_io_out_r_stop_weight;
  wire                pe_mat_18_18_io_out_r_stall;
  wire       [15:0]   pe_mat_18_18_io_out_c_data;
  wire                pe_mat_18_18_io_out_c_is_weight;
  wire       [15:0]   pe_mat_18_19_io_out_r_data;
  wire                pe_mat_18_19_io_out_r_stop_weight;
  wire                pe_mat_18_19_io_out_r_stall;
  wire       [15:0]   pe_mat_18_19_io_out_c_data;
  wire                pe_mat_18_19_io_out_c_is_weight;
  wire       [15:0]   pe_mat_18_20_io_out_r_data;
  wire                pe_mat_18_20_io_out_r_stop_weight;
  wire                pe_mat_18_20_io_out_r_stall;
  wire       [15:0]   pe_mat_18_20_io_out_c_data;
  wire                pe_mat_18_20_io_out_c_is_weight;
  wire       [15:0]   pe_mat_18_21_io_out_r_data;
  wire                pe_mat_18_21_io_out_r_stop_weight;
  wire                pe_mat_18_21_io_out_r_stall;
  wire       [15:0]   pe_mat_18_21_io_out_c_data;
  wire                pe_mat_18_21_io_out_c_is_weight;
  wire       [15:0]   pe_mat_18_22_io_out_r_data;
  wire                pe_mat_18_22_io_out_r_stop_weight;
  wire                pe_mat_18_22_io_out_r_stall;
  wire       [15:0]   pe_mat_18_22_io_out_c_data;
  wire                pe_mat_18_22_io_out_c_is_weight;
  wire       [15:0]   pe_mat_18_23_io_out_r_data;
  wire                pe_mat_18_23_io_out_r_stop_weight;
  wire                pe_mat_18_23_io_out_r_stall;
  wire       [15:0]   pe_mat_18_23_io_out_c_data;
  wire                pe_mat_18_23_io_out_c_is_weight;
  wire       [15:0]   pe_mat_18_24_io_out_r_data;
  wire                pe_mat_18_24_io_out_r_stop_weight;
  wire                pe_mat_18_24_io_out_r_stall;
  wire       [15:0]   pe_mat_18_24_io_out_c_data;
  wire                pe_mat_18_24_io_out_c_is_weight;
  wire       [15:0]   pe_mat_18_25_io_out_r_data;
  wire                pe_mat_18_25_io_out_r_stop_weight;
  wire                pe_mat_18_25_io_out_r_stall;
  wire       [15:0]   pe_mat_18_25_io_out_c_data;
  wire                pe_mat_18_25_io_out_c_is_weight;
  wire       [15:0]   pe_mat_18_26_io_out_r_data;
  wire                pe_mat_18_26_io_out_r_stop_weight;
  wire                pe_mat_18_26_io_out_r_stall;
  wire       [15:0]   pe_mat_18_26_io_out_c_data;
  wire                pe_mat_18_26_io_out_c_is_weight;
  wire       [15:0]   pe_mat_18_27_io_out_r_data;
  wire                pe_mat_18_27_io_out_r_stop_weight;
  wire                pe_mat_18_27_io_out_r_stall;
  wire       [15:0]   pe_mat_18_27_io_out_c_data;
  wire                pe_mat_18_27_io_out_c_is_weight;
  wire       [15:0]   pe_mat_18_28_io_out_r_data;
  wire                pe_mat_18_28_io_out_r_stop_weight;
  wire                pe_mat_18_28_io_out_r_stall;
  wire       [15:0]   pe_mat_18_28_io_out_c_data;
  wire                pe_mat_18_28_io_out_c_is_weight;
  wire       [15:0]   pe_mat_18_29_io_out_r_data;
  wire                pe_mat_18_29_io_out_r_stop_weight;
  wire                pe_mat_18_29_io_out_r_stall;
  wire       [15:0]   pe_mat_18_29_io_out_c_data;
  wire                pe_mat_18_29_io_out_c_is_weight;
  wire       [15:0]   pe_mat_18_30_io_out_r_data;
  wire                pe_mat_18_30_io_out_r_stop_weight;
  wire                pe_mat_18_30_io_out_r_stall;
  wire       [15:0]   pe_mat_18_30_io_out_c_data;
  wire                pe_mat_18_30_io_out_c_is_weight;
  wire       [15:0]   pe_mat_18_31_io_out_r_data;
  wire                pe_mat_18_31_io_out_r_stop_weight;
  wire                pe_mat_18_31_io_out_r_stall;
  wire       [15:0]   pe_mat_18_31_io_out_c_data;
  wire                pe_mat_18_31_io_out_c_is_weight;
  wire       [15:0]   pe_mat_19_0_io_out_r_data;
  wire                pe_mat_19_0_io_out_r_stop_weight;
  wire                pe_mat_19_0_io_out_r_stall;
  wire       [15:0]   pe_mat_19_0_io_out_c_data;
  wire                pe_mat_19_0_io_out_c_is_weight;
  wire       [15:0]   pe_mat_19_1_io_out_r_data;
  wire                pe_mat_19_1_io_out_r_stop_weight;
  wire                pe_mat_19_1_io_out_r_stall;
  wire       [15:0]   pe_mat_19_1_io_out_c_data;
  wire                pe_mat_19_1_io_out_c_is_weight;
  wire       [15:0]   pe_mat_19_2_io_out_r_data;
  wire                pe_mat_19_2_io_out_r_stop_weight;
  wire                pe_mat_19_2_io_out_r_stall;
  wire       [15:0]   pe_mat_19_2_io_out_c_data;
  wire                pe_mat_19_2_io_out_c_is_weight;
  wire       [15:0]   pe_mat_19_3_io_out_r_data;
  wire                pe_mat_19_3_io_out_r_stop_weight;
  wire                pe_mat_19_3_io_out_r_stall;
  wire       [15:0]   pe_mat_19_3_io_out_c_data;
  wire                pe_mat_19_3_io_out_c_is_weight;
  wire       [15:0]   pe_mat_19_4_io_out_r_data;
  wire                pe_mat_19_4_io_out_r_stop_weight;
  wire                pe_mat_19_4_io_out_r_stall;
  wire       [15:0]   pe_mat_19_4_io_out_c_data;
  wire                pe_mat_19_4_io_out_c_is_weight;
  wire       [15:0]   pe_mat_19_5_io_out_r_data;
  wire                pe_mat_19_5_io_out_r_stop_weight;
  wire                pe_mat_19_5_io_out_r_stall;
  wire       [15:0]   pe_mat_19_5_io_out_c_data;
  wire                pe_mat_19_5_io_out_c_is_weight;
  wire       [15:0]   pe_mat_19_6_io_out_r_data;
  wire                pe_mat_19_6_io_out_r_stop_weight;
  wire                pe_mat_19_6_io_out_r_stall;
  wire       [15:0]   pe_mat_19_6_io_out_c_data;
  wire                pe_mat_19_6_io_out_c_is_weight;
  wire       [15:0]   pe_mat_19_7_io_out_r_data;
  wire                pe_mat_19_7_io_out_r_stop_weight;
  wire                pe_mat_19_7_io_out_r_stall;
  wire       [15:0]   pe_mat_19_7_io_out_c_data;
  wire                pe_mat_19_7_io_out_c_is_weight;
  wire       [15:0]   pe_mat_19_8_io_out_r_data;
  wire                pe_mat_19_8_io_out_r_stop_weight;
  wire                pe_mat_19_8_io_out_r_stall;
  wire       [15:0]   pe_mat_19_8_io_out_c_data;
  wire                pe_mat_19_8_io_out_c_is_weight;
  wire       [15:0]   pe_mat_19_9_io_out_r_data;
  wire                pe_mat_19_9_io_out_r_stop_weight;
  wire                pe_mat_19_9_io_out_r_stall;
  wire       [15:0]   pe_mat_19_9_io_out_c_data;
  wire                pe_mat_19_9_io_out_c_is_weight;
  wire       [15:0]   pe_mat_19_10_io_out_r_data;
  wire                pe_mat_19_10_io_out_r_stop_weight;
  wire                pe_mat_19_10_io_out_r_stall;
  wire       [15:0]   pe_mat_19_10_io_out_c_data;
  wire                pe_mat_19_10_io_out_c_is_weight;
  wire       [15:0]   pe_mat_19_11_io_out_r_data;
  wire                pe_mat_19_11_io_out_r_stop_weight;
  wire                pe_mat_19_11_io_out_r_stall;
  wire       [15:0]   pe_mat_19_11_io_out_c_data;
  wire                pe_mat_19_11_io_out_c_is_weight;
  wire       [15:0]   pe_mat_19_12_io_out_r_data;
  wire                pe_mat_19_12_io_out_r_stop_weight;
  wire                pe_mat_19_12_io_out_r_stall;
  wire       [15:0]   pe_mat_19_12_io_out_c_data;
  wire                pe_mat_19_12_io_out_c_is_weight;
  wire       [15:0]   pe_mat_19_13_io_out_r_data;
  wire                pe_mat_19_13_io_out_r_stop_weight;
  wire                pe_mat_19_13_io_out_r_stall;
  wire       [15:0]   pe_mat_19_13_io_out_c_data;
  wire                pe_mat_19_13_io_out_c_is_weight;
  wire       [15:0]   pe_mat_19_14_io_out_r_data;
  wire                pe_mat_19_14_io_out_r_stop_weight;
  wire                pe_mat_19_14_io_out_r_stall;
  wire       [15:0]   pe_mat_19_14_io_out_c_data;
  wire                pe_mat_19_14_io_out_c_is_weight;
  wire       [15:0]   pe_mat_19_15_io_out_r_data;
  wire                pe_mat_19_15_io_out_r_stop_weight;
  wire                pe_mat_19_15_io_out_r_stall;
  wire       [15:0]   pe_mat_19_15_io_out_c_data;
  wire                pe_mat_19_15_io_out_c_is_weight;
  wire       [15:0]   pe_mat_19_16_io_out_r_data;
  wire                pe_mat_19_16_io_out_r_stop_weight;
  wire                pe_mat_19_16_io_out_r_stall;
  wire       [15:0]   pe_mat_19_16_io_out_c_data;
  wire                pe_mat_19_16_io_out_c_is_weight;
  wire       [15:0]   pe_mat_19_17_io_out_r_data;
  wire                pe_mat_19_17_io_out_r_stop_weight;
  wire                pe_mat_19_17_io_out_r_stall;
  wire       [15:0]   pe_mat_19_17_io_out_c_data;
  wire                pe_mat_19_17_io_out_c_is_weight;
  wire       [15:0]   pe_mat_19_18_io_out_r_data;
  wire                pe_mat_19_18_io_out_r_stop_weight;
  wire                pe_mat_19_18_io_out_r_stall;
  wire       [15:0]   pe_mat_19_18_io_out_c_data;
  wire                pe_mat_19_18_io_out_c_is_weight;
  wire       [15:0]   pe_mat_19_19_io_out_r_data;
  wire                pe_mat_19_19_io_out_r_stop_weight;
  wire                pe_mat_19_19_io_out_r_stall;
  wire       [15:0]   pe_mat_19_19_io_out_c_data;
  wire                pe_mat_19_19_io_out_c_is_weight;
  wire       [15:0]   pe_mat_19_20_io_out_r_data;
  wire                pe_mat_19_20_io_out_r_stop_weight;
  wire                pe_mat_19_20_io_out_r_stall;
  wire       [15:0]   pe_mat_19_20_io_out_c_data;
  wire                pe_mat_19_20_io_out_c_is_weight;
  wire       [15:0]   pe_mat_19_21_io_out_r_data;
  wire                pe_mat_19_21_io_out_r_stop_weight;
  wire                pe_mat_19_21_io_out_r_stall;
  wire       [15:0]   pe_mat_19_21_io_out_c_data;
  wire                pe_mat_19_21_io_out_c_is_weight;
  wire       [15:0]   pe_mat_19_22_io_out_r_data;
  wire                pe_mat_19_22_io_out_r_stop_weight;
  wire                pe_mat_19_22_io_out_r_stall;
  wire       [15:0]   pe_mat_19_22_io_out_c_data;
  wire                pe_mat_19_22_io_out_c_is_weight;
  wire       [15:0]   pe_mat_19_23_io_out_r_data;
  wire                pe_mat_19_23_io_out_r_stop_weight;
  wire                pe_mat_19_23_io_out_r_stall;
  wire       [15:0]   pe_mat_19_23_io_out_c_data;
  wire                pe_mat_19_23_io_out_c_is_weight;
  wire       [15:0]   pe_mat_19_24_io_out_r_data;
  wire                pe_mat_19_24_io_out_r_stop_weight;
  wire                pe_mat_19_24_io_out_r_stall;
  wire       [15:0]   pe_mat_19_24_io_out_c_data;
  wire                pe_mat_19_24_io_out_c_is_weight;
  wire       [15:0]   pe_mat_19_25_io_out_r_data;
  wire                pe_mat_19_25_io_out_r_stop_weight;
  wire                pe_mat_19_25_io_out_r_stall;
  wire       [15:0]   pe_mat_19_25_io_out_c_data;
  wire                pe_mat_19_25_io_out_c_is_weight;
  wire       [15:0]   pe_mat_19_26_io_out_r_data;
  wire                pe_mat_19_26_io_out_r_stop_weight;
  wire                pe_mat_19_26_io_out_r_stall;
  wire       [15:0]   pe_mat_19_26_io_out_c_data;
  wire                pe_mat_19_26_io_out_c_is_weight;
  wire       [15:0]   pe_mat_19_27_io_out_r_data;
  wire                pe_mat_19_27_io_out_r_stop_weight;
  wire                pe_mat_19_27_io_out_r_stall;
  wire       [15:0]   pe_mat_19_27_io_out_c_data;
  wire                pe_mat_19_27_io_out_c_is_weight;
  wire       [15:0]   pe_mat_19_28_io_out_r_data;
  wire                pe_mat_19_28_io_out_r_stop_weight;
  wire                pe_mat_19_28_io_out_r_stall;
  wire       [15:0]   pe_mat_19_28_io_out_c_data;
  wire                pe_mat_19_28_io_out_c_is_weight;
  wire       [15:0]   pe_mat_19_29_io_out_r_data;
  wire                pe_mat_19_29_io_out_r_stop_weight;
  wire                pe_mat_19_29_io_out_r_stall;
  wire       [15:0]   pe_mat_19_29_io_out_c_data;
  wire                pe_mat_19_29_io_out_c_is_weight;
  wire       [15:0]   pe_mat_19_30_io_out_r_data;
  wire                pe_mat_19_30_io_out_r_stop_weight;
  wire                pe_mat_19_30_io_out_r_stall;
  wire       [15:0]   pe_mat_19_30_io_out_c_data;
  wire                pe_mat_19_30_io_out_c_is_weight;
  wire       [15:0]   pe_mat_19_31_io_out_r_data;
  wire                pe_mat_19_31_io_out_r_stop_weight;
  wire                pe_mat_19_31_io_out_r_stall;
  wire       [15:0]   pe_mat_19_31_io_out_c_data;
  wire                pe_mat_19_31_io_out_c_is_weight;
  wire       [15:0]   pe_mat_20_0_io_out_r_data;
  wire                pe_mat_20_0_io_out_r_stop_weight;
  wire                pe_mat_20_0_io_out_r_stall;
  wire       [15:0]   pe_mat_20_0_io_out_c_data;
  wire                pe_mat_20_0_io_out_c_is_weight;
  wire       [15:0]   pe_mat_20_1_io_out_r_data;
  wire                pe_mat_20_1_io_out_r_stop_weight;
  wire                pe_mat_20_1_io_out_r_stall;
  wire       [15:0]   pe_mat_20_1_io_out_c_data;
  wire                pe_mat_20_1_io_out_c_is_weight;
  wire       [15:0]   pe_mat_20_2_io_out_r_data;
  wire                pe_mat_20_2_io_out_r_stop_weight;
  wire                pe_mat_20_2_io_out_r_stall;
  wire       [15:0]   pe_mat_20_2_io_out_c_data;
  wire                pe_mat_20_2_io_out_c_is_weight;
  wire       [15:0]   pe_mat_20_3_io_out_r_data;
  wire                pe_mat_20_3_io_out_r_stop_weight;
  wire                pe_mat_20_3_io_out_r_stall;
  wire       [15:0]   pe_mat_20_3_io_out_c_data;
  wire                pe_mat_20_3_io_out_c_is_weight;
  wire       [15:0]   pe_mat_20_4_io_out_r_data;
  wire                pe_mat_20_4_io_out_r_stop_weight;
  wire                pe_mat_20_4_io_out_r_stall;
  wire       [15:0]   pe_mat_20_4_io_out_c_data;
  wire                pe_mat_20_4_io_out_c_is_weight;
  wire       [15:0]   pe_mat_20_5_io_out_r_data;
  wire                pe_mat_20_5_io_out_r_stop_weight;
  wire                pe_mat_20_5_io_out_r_stall;
  wire       [15:0]   pe_mat_20_5_io_out_c_data;
  wire                pe_mat_20_5_io_out_c_is_weight;
  wire       [15:0]   pe_mat_20_6_io_out_r_data;
  wire                pe_mat_20_6_io_out_r_stop_weight;
  wire                pe_mat_20_6_io_out_r_stall;
  wire       [15:0]   pe_mat_20_6_io_out_c_data;
  wire                pe_mat_20_6_io_out_c_is_weight;
  wire       [15:0]   pe_mat_20_7_io_out_r_data;
  wire                pe_mat_20_7_io_out_r_stop_weight;
  wire                pe_mat_20_7_io_out_r_stall;
  wire       [15:0]   pe_mat_20_7_io_out_c_data;
  wire                pe_mat_20_7_io_out_c_is_weight;
  wire       [15:0]   pe_mat_20_8_io_out_r_data;
  wire                pe_mat_20_8_io_out_r_stop_weight;
  wire                pe_mat_20_8_io_out_r_stall;
  wire       [15:0]   pe_mat_20_8_io_out_c_data;
  wire                pe_mat_20_8_io_out_c_is_weight;
  wire       [15:0]   pe_mat_20_9_io_out_r_data;
  wire                pe_mat_20_9_io_out_r_stop_weight;
  wire                pe_mat_20_9_io_out_r_stall;
  wire       [15:0]   pe_mat_20_9_io_out_c_data;
  wire                pe_mat_20_9_io_out_c_is_weight;
  wire       [15:0]   pe_mat_20_10_io_out_r_data;
  wire                pe_mat_20_10_io_out_r_stop_weight;
  wire                pe_mat_20_10_io_out_r_stall;
  wire       [15:0]   pe_mat_20_10_io_out_c_data;
  wire                pe_mat_20_10_io_out_c_is_weight;
  wire       [15:0]   pe_mat_20_11_io_out_r_data;
  wire                pe_mat_20_11_io_out_r_stop_weight;
  wire                pe_mat_20_11_io_out_r_stall;
  wire       [15:0]   pe_mat_20_11_io_out_c_data;
  wire                pe_mat_20_11_io_out_c_is_weight;
  wire       [15:0]   pe_mat_20_12_io_out_r_data;
  wire                pe_mat_20_12_io_out_r_stop_weight;
  wire                pe_mat_20_12_io_out_r_stall;
  wire       [15:0]   pe_mat_20_12_io_out_c_data;
  wire                pe_mat_20_12_io_out_c_is_weight;
  wire       [15:0]   pe_mat_20_13_io_out_r_data;
  wire                pe_mat_20_13_io_out_r_stop_weight;
  wire                pe_mat_20_13_io_out_r_stall;
  wire       [15:0]   pe_mat_20_13_io_out_c_data;
  wire                pe_mat_20_13_io_out_c_is_weight;
  wire       [15:0]   pe_mat_20_14_io_out_r_data;
  wire                pe_mat_20_14_io_out_r_stop_weight;
  wire                pe_mat_20_14_io_out_r_stall;
  wire       [15:0]   pe_mat_20_14_io_out_c_data;
  wire                pe_mat_20_14_io_out_c_is_weight;
  wire       [15:0]   pe_mat_20_15_io_out_r_data;
  wire                pe_mat_20_15_io_out_r_stop_weight;
  wire                pe_mat_20_15_io_out_r_stall;
  wire       [15:0]   pe_mat_20_15_io_out_c_data;
  wire                pe_mat_20_15_io_out_c_is_weight;
  wire       [15:0]   pe_mat_20_16_io_out_r_data;
  wire                pe_mat_20_16_io_out_r_stop_weight;
  wire                pe_mat_20_16_io_out_r_stall;
  wire       [15:0]   pe_mat_20_16_io_out_c_data;
  wire                pe_mat_20_16_io_out_c_is_weight;
  wire       [15:0]   pe_mat_20_17_io_out_r_data;
  wire                pe_mat_20_17_io_out_r_stop_weight;
  wire                pe_mat_20_17_io_out_r_stall;
  wire       [15:0]   pe_mat_20_17_io_out_c_data;
  wire                pe_mat_20_17_io_out_c_is_weight;
  wire       [15:0]   pe_mat_20_18_io_out_r_data;
  wire                pe_mat_20_18_io_out_r_stop_weight;
  wire                pe_mat_20_18_io_out_r_stall;
  wire       [15:0]   pe_mat_20_18_io_out_c_data;
  wire                pe_mat_20_18_io_out_c_is_weight;
  wire       [15:0]   pe_mat_20_19_io_out_r_data;
  wire                pe_mat_20_19_io_out_r_stop_weight;
  wire                pe_mat_20_19_io_out_r_stall;
  wire       [15:0]   pe_mat_20_19_io_out_c_data;
  wire                pe_mat_20_19_io_out_c_is_weight;
  wire       [15:0]   pe_mat_20_20_io_out_r_data;
  wire                pe_mat_20_20_io_out_r_stop_weight;
  wire                pe_mat_20_20_io_out_r_stall;
  wire       [15:0]   pe_mat_20_20_io_out_c_data;
  wire                pe_mat_20_20_io_out_c_is_weight;
  wire       [15:0]   pe_mat_20_21_io_out_r_data;
  wire                pe_mat_20_21_io_out_r_stop_weight;
  wire                pe_mat_20_21_io_out_r_stall;
  wire       [15:0]   pe_mat_20_21_io_out_c_data;
  wire                pe_mat_20_21_io_out_c_is_weight;
  wire       [15:0]   pe_mat_20_22_io_out_r_data;
  wire                pe_mat_20_22_io_out_r_stop_weight;
  wire                pe_mat_20_22_io_out_r_stall;
  wire       [15:0]   pe_mat_20_22_io_out_c_data;
  wire                pe_mat_20_22_io_out_c_is_weight;
  wire       [15:0]   pe_mat_20_23_io_out_r_data;
  wire                pe_mat_20_23_io_out_r_stop_weight;
  wire                pe_mat_20_23_io_out_r_stall;
  wire       [15:0]   pe_mat_20_23_io_out_c_data;
  wire                pe_mat_20_23_io_out_c_is_weight;
  wire       [15:0]   pe_mat_20_24_io_out_r_data;
  wire                pe_mat_20_24_io_out_r_stop_weight;
  wire                pe_mat_20_24_io_out_r_stall;
  wire       [15:0]   pe_mat_20_24_io_out_c_data;
  wire                pe_mat_20_24_io_out_c_is_weight;
  wire       [15:0]   pe_mat_20_25_io_out_r_data;
  wire                pe_mat_20_25_io_out_r_stop_weight;
  wire                pe_mat_20_25_io_out_r_stall;
  wire       [15:0]   pe_mat_20_25_io_out_c_data;
  wire                pe_mat_20_25_io_out_c_is_weight;
  wire       [15:0]   pe_mat_20_26_io_out_r_data;
  wire                pe_mat_20_26_io_out_r_stop_weight;
  wire                pe_mat_20_26_io_out_r_stall;
  wire       [15:0]   pe_mat_20_26_io_out_c_data;
  wire                pe_mat_20_26_io_out_c_is_weight;
  wire       [15:0]   pe_mat_20_27_io_out_r_data;
  wire                pe_mat_20_27_io_out_r_stop_weight;
  wire                pe_mat_20_27_io_out_r_stall;
  wire       [15:0]   pe_mat_20_27_io_out_c_data;
  wire                pe_mat_20_27_io_out_c_is_weight;
  wire       [15:0]   pe_mat_20_28_io_out_r_data;
  wire                pe_mat_20_28_io_out_r_stop_weight;
  wire                pe_mat_20_28_io_out_r_stall;
  wire       [15:0]   pe_mat_20_28_io_out_c_data;
  wire                pe_mat_20_28_io_out_c_is_weight;
  wire       [15:0]   pe_mat_20_29_io_out_r_data;
  wire                pe_mat_20_29_io_out_r_stop_weight;
  wire                pe_mat_20_29_io_out_r_stall;
  wire       [15:0]   pe_mat_20_29_io_out_c_data;
  wire                pe_mat_20_29_io_out_c_is_weight;
  wire       [15:0]   pe_mat_20_30_io_out_r_data;
  wire                pe_mat_20_30_io_out_r_stop_weight;
  wire                pe_mat_20_30_io_out_r_stall;
  wire       [15:0]   pe_mat_20_30_io_out_c_data;
  wire                pe_mat_20_30_io_out_c_is_weight;
  wire       [15:0]   pe_mat_20_31_io_out_r_data;
  wire                pe_mat_20_31_io_out_r_stop_weight;
  wire                pe_mat_20_31_io_out_r_stall;
  wire       [15:0]   pe_mat_20_31_io_out_c_data;
  wire                pe_mat_20_31_io_out_c_is_weight;
  wire       [15:0]   pe_mat_21_0_io_out_r_data;
  wire                pe_mat_21_0_io_out_r_stop_weight;
  wire                pe_mat_21_0_io_out_r_stall;
  wire       [15:0]   pe_mat_21_0_io_out_c_data;
  wire                pe_mat_21_0_io_out_c_is_weight;
  wire       [15:0]   pe_mat_21_1_io_out_r_data;
  wire                pe_mat_21_1_io_out_r_stop_weight;
  wire                pe_mat_21_1_io_out_r_stall;
  wire       [15:0]   pe_mat_21_1_io_out_c_data;
  wire                pe_mat_21_1_io_out_c_is_weight;
  wire       [15:0]   pe_mat_21_2_io_out_r_data;
  wire                pe_mat_21_2_io_out_r_stop_weight;
  wire                pe_mat_21_2_io_out_r_stall;
  wire       [15:0]   pe_mat_21_2_io_out_c_data;
  wire                pe_mat_21_2_io_out_c_is_weight;
  wire       [15:0]   pe_mat_21_3_io_out_r_data;
  wire                pe_mat_21_3_io_out_r_stop_weight;
  wire                pe_mat_21_3_io_out_r_stall;
  wire       [15:0]   pe_mat_21_3_io_out_c_data;
  wire                pe_mat_21_3_io_out_c_is_weight;
  wire       [15:0]   pe_mat_21_4_io_out_r_data;
  wire                pe_mat_21_4_io_out_r_stop_weight;
  wire                pe_mat_21_4_io_out_r_stall;
  wire       [15:0]   pe_mat_21_4_io_out_c_data;
  wire                pe_mat_21_4_io_out_c_is_weight;
  wire       [15:0]   pe_mat_21_5_io_out_r_data;
  wire                pe_mat_21_5_io_out_r_stop_weight;
  wire                pe_mat_21_5_io_out_r_stall;
  wire       [15:0]   pe_mat_21_5_io_out_c_data;
  wire                pe_mat_21_5_io_out_c_is_weight;
  wire       [15:0]   pe_mat_21_6_io_out_r_data;
  wire                pe_mat_21_6_io_out_r_stop_weight;
  wire                pe_mat_21_6_io_out_r_stall;
  wire       [15:0]   pe_mat_21_6_io_out_c_data;
  wire                pe_mat_21_6_io_out_c_is_weight;
  wire       [15:0]   pe_mat_21_7_io_out_r_data;
  wire                pe_mat_21_7_io_out_r_stop_weight;
  wire                pe_mat_21_7_io_out_r_stall;
  wire       [15:0]   pe_mat_21_7_io_out_c_data;
  wire                pe_mat_21_7_io_out_c_is_weight;
  wire       [15:0]   pe_mat_21_8_io_out_r_data;
  wire                pe_mat_21_8_io_out_r_stop_weight;
  wire                pe_mat_21_8_io_out_r_stall;
  wire       [15:0]   pe_mat_21_8_io_out_c_data;
  wire                pe_mat_21_8_io_out_c_is_weight;
  wire       [15:0]   pe_mat_21_9_io_out_r_data;
  wire                pe_mat_21_9_io_out_r_stop_weight;
  wire                pe_mat_21_9_io_out_r_stall;
  wire       [15:0]   pe_mat_21_9_io_out_c_data;
  wire                pe_mat_21_9_io_out_c_is_weight;
  wire       [15:0]   pe_mat_21_10_io_out_r_data;
  wire                pe_mat_21_10_io_out_r_stop_weight;
  wire                pe_mat_21_10_io_out_r_stall;
  wire       [15:0]   pe_mat_21_10_io_out_c_data;
  wire                pe_mat_21_10_io_out_c_is_weight;
  wire       [15:0]   pe_mat_21_11_io_out_r_data;
  wire                pe_mat_21_11_io_out_r_stop_weight;
  wire                pe_mat_21_11_io_out_r_stall;
  wire       [15:0]   pe_mat_21_11_io_out_c_data;
  wire                pe_mat_21_11_io_out_c_is_weight;
  wire       [15:0]   pe_mat_21_12_io_out_r_data;
  wire                pe_mat_21_12_io_out_r_stop_weight;
  wire                pe_mat_21_12_io_out_r_stall;
  wire       [15:0]   pe_mat_21_12_io_out_c_data;
  wire                pe_mat_21_12_io_out_c_is_weight;
  wire       [15:0]   pe_mat_21_13_io_out_r_data;
  wire                pe_mat_21_13_io_out_r_stop_weight;
  wire                pe_mat_21_13_io_out_r_stall;
  wire       [15:0]   pe_mat_21_13_io_out_c_data;
  wire                pe_mat_21_13_io_out_c_is_weight;
  wire       [15:0]   pe_mat_21_14_io_out_r_data;
  wire                pe_mat_21_14_io_out_r_stop_weight;
  wire                pe_mat_21_14_io_out_r_stall;
  wire       [15:0]   pe_mat_21_14_io_out_c_data;
  wire                pe_mat_21_14_io_out_c_is_weight;
  wire       [15:0]   pe_mat_21_15_io_out_r_data;
  wire                pe_mat_21_15_io_out_r_stop_weight;
  wire                pe_mat_21_15_io_out_r_stall;
  wire       [15:0]   pe_mat_21_15_io_out_c_data;
  wire                pe_mat_21_15_io_out_c_is_weight;
  wire       [15:0]   pe_mat_21_16_io_out_r_data;
  wire                pe_mat_21_16_io_out_r_stop_weight;
  wire                pe_mat_21_16_io_out_r_stall;
  wire       [15:0]   pe_mat_21_16_io_out_c_data;
  wire                pe_mat_21_16_io_out_c_is_weight;
  wire       [15:0]   pe_mat_21_17_io_out_r_data;
  wire                pe_mat_21_17_io_out_r_stop_weight;
  wire                pe_mat_21_17_io_out_r_stall;
  wire       [15:0]   pe_mat_21_17_io_out_c_data;
  wire                pe_mat_21_17_io_out_c_is_weight;
  wire       [15:0]   pe_mat_21_18_io_out_r_data;
  wire                pe_mat_21_18_io_out_r_stop_weight;
  wire                pe_mat_21_18_io_out_r_stall;
  wire       [15:0]   pe_mat_21_18_io_out_c_data;
  wire                pe_mat_21_18_io_out_c_is_weight;
  wire       [15:0]   pe_mat_21_19_io_out_r_data;
  wire                pe_mat_21_19_io_out_r_stop_weight;
  wire                pe_mat_21_19_io_out_r_stall;
  wire       [15:0]   pe_mat_21_19_io_out_c_data;
  wire                pe_mat_21_19_io_out_c_is_weight;
  wire       [15:0]   pe_mat_21_20_io_out_r_data;
  wire                pe_mat_21_20_io_out_r_stop_weight;
  wire                pe_mat_21_20_io_out_r_stall;
  wire       [15:0]   pe_mat_21_20_io_out_c_data;
  wire                pe_mat_21_20_io_out_c_is_weight;
  wire       [15:0]   pe_mat_21_21_io_out_r_data;
  wire                pe_mat_21_21_io_out_r_stop_weight;
  wire                pe_mat_21_21_io_out_r_stall;
  wire       [15:0]   pe_mat_21_21_io_out_c_data;
  wire                pe_mat_21_21_io_out_c_is_weight;
  wire       [15:0]   pe_mat_21_22_io_out_r_data;
  wire                pe_mat_21_22_io_out_r_stop_weight;
  wire                pe_mat_21_22_io_out_r_stall;
  wire       [15:0]   pe_mat_21_22_io_out_c_data;
  wire                pe_mat_21_22_io_out_c_is_weight;
  wire       [15:0]   pe_mat_21_23_io_out_r_data;
  wire                pe_mat_21_23_io_out_r_stop_weight;
  wire                pe_mat_21_23_io_out_r_stall;
  wire       [15:0]   pe_mat_21_23_io_out_c_data;
  wire                pe_mat_21_23_io_out_c_is_weight;
  wire       [15:0]   pe_mat_21_24_io_out_r_data;
  wire                pe_mat_21_24_io_out_r_stop_weight;
  wire                pe_mat_21_24_io_out_r_stall;
  wire       [15:0]   pe_mat_21_24_io_out_c_data;
  wire                pe_mat_21_24_io_out_c_is_weight;
  wire       [15:0]   pe_mat_21_25_io_out_r_data;
  wire                pe_mat_21_25_io_out_r_stop_weight;
  wire                pe_mat_21_25_io_out_r_stall;
  wire       [15:0]   pe_mat_21_25_io_out_c_data;
  wire                pe_mat_21_25_io_out_c_is_weight;
  wire       [15:0]   pe_mat_21_26_io_out_r_data;
  wire                pe_mat_21_26_io_out_r_stop_weight;
  wire                pe_mat_21_26_io_out_r_stall;
  wire       [15:0]   pe_mat_21_26_io_out_c_data;
  wire                pe_mat_21_26_io_out_c_is_weight;
  wire       [15:0]   pe_mat_21_27_io_out_r_data;
  wire                pe_mat_21_27_io_out_r_stop_weight;
  wire                pe_mat_21_27_io_out_r_stall;
  wire       [15:0]   pe_mat_21_27_io_out_c_data;
  wire                pe_mat_21_27_io_out_c_is_weight;
  wire       [15:0]   pe_mat_21_28_io_out_r_data;
  wire                pe_mat_21_28_io_out_r_stop_weight;
  wire                pe_mat_21_28_io_out_r_stall;
  wire       [15:0]   pe_mat_21_28_io_out_c_data;
  wire                pe_mat_21_28_io_out_c_is_weight;
  wire       [15:0]   pe_mat_21_29_io_out_r_data;
  wire                pe_mat_21_29_io_out_r_stop_weight;
  wire                pe_mat_21_29_io_out_r_stall;
  wire       [15:0]   pe_mat_21_29_io_out_c_data;
  wire                pe_mat_21_29_io_out_c_is_weight;
  wire       [15:0]   pe_mat_21_30_io_out_r_data;
  wire                pe_mat_21_30_io_out_r_stop_weight;
  wire                pe_mat_21_30_io_out_r_stall;
  wire       [15:0]   pe_mat_21_30_io_out_c_data;
  wire                pe_mat_21_30_io_out_c_is_weight;
  wire       [15:0]   pe_mat_21_31_io_out_r_data;
  wire                pe_mat_21_31_io_out_r_stop_weight;
  wire                pe_mat_21_31_io_out_r_stall;
  wire       [15:0]   pe_mat_21_31_io_out_c_data;
  wire                pe_mat_21_31_io_out_c_is_weight;
  wire       [15:0]   pe_mat_22_0_io_out_r_data;
  wire                pe_mat_22_0_io_out_r_stop_weight;
  wire                pe_mat_22_0_io_out_r_stall;
  wire       [15:0]   pe_mat_22_0_io_out_c_data;
  wire                pe_mat_22_0_io_out_c_is_weight;
  wire       [15:0]   pe_mat_22_1_io_out_r_data;
  wire                pe_mat_22_1_io_out_r_stop_weight;
  wire                pe_mat_22_1_io_out_r_stall;
  wire       [15:0]   pe_mat_22_1_io_out_c_data;
  wire                pe_mat_22_1_io_out_c_is_weight;
  wire       [15:0]   pe_mat_22_2_io_out_r_data;
  wire                pe_mat_22_2_io_out_r_stop_weight;
  wire                pe_mat_22_2_io_out_r_stall;
  wire       [15:0]   pe_mat_22_2_io_out_c_data;
  wire                pe_mat_22_2_io_out_c_is_weight;
  wire       [15:0]   pe_mat_22_3_io_out_r_data;
  wire                pe_mat_22_3_io_out_r_stop_weight;
  wire                pe_mat_22_3_io_out_r_stall;
  wire       [15:0]   pe_mat_22_3_io_out_c_data;
  wire                pe_mat_22_3_io_out_c_is_weight;
  wire       [15:0]   pe_mat_22_4_io_out_r_data;
  wire                pe_mat_22_4_io_out_r_stop_weight;
  wire                pe_mat_22_4_io_out_r_stall;
  wire       [15:0]   pe_mat_22_4_io_out_c_data;
  wire                pe_mat_22_4_io_out_c_is_weight;
  wire       [15:0]   pe_mat_22_5_io_out_r_data;
  wire                pe_mat_22_5_io_out_r_stop_weight;
  wire                pe_mat_22_5_io_out_r_stall;
  wire       [15:0]   pe_mat_22_5_io_out_c_data;
  wire                pe_mat_22_5_io_out_c_is_weight;
  wire       [15:0]   pe_mat_22_6_io_out_r_data;
  wire                pe_mat_22_6_io_out_r_stop_weight;
  wire                pe_mat_22_6_io_out_r_stall;
  wire       [15:0]   pe_mat_22_6_io_out_c_data;
  wire                pe_mat_22_6_io_out_c_is_weight;
  wire       [15:0]   pe_mat_22_7_io_out_r_data;
  wire                pe_mat_22_7_io_out_r_stop_weight;
  wire                pe_mat_22_7_io_out_r_stall;
  wire       [15:0]   pe_mat_22_7_io_out_c_data;
  wire                pe_mat_22_7_io_out_c_is_weight;
  wire       [15:0]   pe_mat_22_8_io_out_r_data;
  wire                pe_mat_22_8_io_out_r_stop_weight;
  wire                pe_mat_22_8_io_out_r_stall;
  wire       [15:0]   pe_mat_22_8_io_out_c_data;
  wire                pe_mat_22_8_io_out_c_is_weight;
  wire       [15:0]   pe_mat_22_9_io_out_r_data;
  wire                pe_mat_22_9_io_out_r_stop_weight;
  wire                pe_mat_22_9_io_out_r_stall;
  wire       [15:0]   pe_mat_22_9_io_out_c_data;
  wire                pe_mat_22_9_io_out_c_is_weight;
  wire       [15:0]   pe_mat_22_10_io_out_r_data;
  wire                pe_mat_22_10_io_out_r_stop_weight;
  wire                pe_mat_22_10_io_out_r_stall;
  wire       [15:0]   pe_mat_22_10_io_out_c_data;
  wire                pe_mat_22_10_io_out_c_is_weight;
  wire       [15:0]   pe_mat_22_11_io_out_r_data;
  wire                pe_mat_22_11_io_out_r_stop_weight;
  wire                pe_mat_22_11_io_out_r_stall;
  wire       [15:0]   pe_mat_22_11_io_out_c_data;
  wire                pe_mat_22_11_io_out_c_is_weight;
  wire       [15:0]   pe_mat_22_12_io_out_r_data;
  wire                pe_mat_22_12_io_out_r_stop_weight;
  wire                pe_mat_22_12_io_out_r_stall;
  wire       [15:0]   pe_mat_22_12_io_out_c_data;
  wire                pe_mat_22_12_io_out_c_is_weight;
  wire       [15:0]   pe_mat_22_13_io_out_r_data;
  wire                pe_mat_22_13_io_out_r_stop_weight;
  wire                pe_mat_22_13_io_out_r_stall;
  wire       [15:0]   pe_mat_22_13_io_out_c_data;
  wire                pe_mat_22_13_io_out_c_is_weight;
  wire       [15:0]   pe_mat_22_14_io_out_r_data;
  wire                pe_mat_22_14_io_out_r_stop_weight;
  wire                pe_mat_22_14_io_out_r_stall;
  wire       [15:0]   pe_mat_22_14_io_out_c_data;
  wire                pe_mat_22_14_io_out_c_is_weight;
  wire       [15:0]   pe_mat_22_15_io_out_r_data;
  wire                pe_mat_22_15_io_out_r_stop_weight;
  wire                pe_mat_22_15_io_out_r_stall;
  wire       [15:0]   pe_mat_22_15_io_out_c_data;
  wire                pe_mat_22_15_io_out_c_is_weight;
  wire       [15:0]   pe_mat_22_16_io_out_r_data;
  wire                pe_mat_22_16_io_out_r_stop_weight;
  wire                pe_mat_22_16_io_out_r_stall;
  wire       [15:0]   pe_mat_22_16_io_out_c_data;
  wire                pe_mat_22_16_io_out_c_is_weight;
  wire       [15:0]   pe_mat_22_17_io_out_r_data;
  wire                pe_mat_22_17_io_out_r_stop_weight;
  wire                pe_mat_22_17_io_out_r_stall;
  wire       [15:0]   pe_mat_22_17_io_out_c_data;
  wire                pe_mat_22_17_io_out_c_is_weight;
  wire       [15:0]   pe_mat_22_18_io_out_r_data;
  wire                pe_mat_22_18_io_out_r_stop_weight;
  wire                pe_mat_22_18_io_out_r_stall;
  wire       [15:0]   pe_mat_22_18_io_out_c_data;
  wire                pe_mat_22_18_io_out_c_is_weight;
  wire       [15:0]   pe_mat_22_19_io_out_r_data;
  wire                pe_mat_22_19_io_out_r_stop_weight;
  wire                pe_mat_22_19_io_out_r_stall;
  wire       [15:0]   pe_mat_22_19_io_out_c_data;
  wire                pe_mat_22_19_io_out_c_is_weight;
  wire       [15:0]   pe_mat_22_20_io_out_r_data;
  wire                pe_mat_22_20_io_out_r_stop_weight;
  wire                pe_mat_22_20_io_out_r_stall;
  wire       [15:0]   pe_mat_22_20_io_out_c_data;
  wire                pe_mat_22_20_io_out_c_is_weight;
  wire       [15:0]   pe_mat_22_21_io_out_r_data;
  wire                pe_mat_22_21_io_out_r_stop_weight;
  wire                pe_mat_22_21_io_out_r_stall;
  wire       [15:0]   pe_mat_22_21_io_out_c_data;
  wire                pe_mat_22_21_io_out_c_is_weight;
  wire       [15:0]   pe_mat_22_22_io_out_r_data;
  wire                pe_mat_22_22_io_out_r_stop_weight;
  wire                pe_mat_22_22_io_out_r_stall;
  wire       [15:0]   pe_mat_22_22_io_out_c_data;
  wire                pe_mat_22_22_io_out_c_is_weight;
  wire       [15:0]   pe_mat_22_23_io_out_r_data;
  wire                pe_mat_22_23_io_out_r_stop_weight;
  wire                pe_mat_22_23_io_out_r_stall;
  wire       [15:0]   pe_mat_22_23_io_out_c_data;
  wire                pe_mat_22_23_io_out_c_is_weight;
  wire       [15:0]   pe_mat_22_24_io_out_r_data;
  wire                pe_mat_22_24_io_out_r_stop_weight;
  wire                pe_mat_22_24_io_out_r_stall;
  wire       [15:0]   pe_mat_22_24_io_out_c_data;
  wire                pe_mat_22_24_io_out_c_is_weight;
  wire       [15:0]   pe_mat_22_25_io_out_r_data;
  wire                pe_mat_22_25_io_out_r_stop_weight;
  wire                pe_mat_22_25_io_out_r_stall;
  wire       [15:0]   pe_mat_22_25_io_out_c_data;
  wire                pe_mat_22_25_io_out_c_is_weight;
  wire       [15:0]   pe_mat_22_26_io_out_r_data;
  wire                pe_mat_22_26_io_out_r_stop_weight;
  wire                pe_mat_22_26_io_out_r_stall;
  wire       [15:0]   pe_mat_22_26_io_out_c_data;
  wire                pe_mat_22_26_io_out_c_is_weight;
  wire       [15:0]   pe_mat_22_27_io_out_r_data;
  wire                pe_mat_22_27_io_out_r_stop_weight;
  wire                pe_mat_22_27_io_out_r_stall;
  wire       [15:0]   pe_mat_22_27_io_out_c_data;
  wire                pe_mat_22_27_io_out_c_is_weight;
  wire       [15:0]   pe_mat_22_28_io_out_r_data;
  wire                pe_mat_22_28_io_out_r_stop_weight;
  wire                pe_mat_22_28_io_out_r_stall;
  wire       [15:0]   pe_mat_22_28_io_out_c_data;
  wire                pe_mat_22_28_io_out_c_is_weight;
  wire       [15:0]   pe_mat_22_29_io_out_r_data;
  wire                pe_mat_22_29_io_out_r_stop_weight;
  wire                pe_mat_22_29_io_out_r_stall;
  wire       [15:0]   pe_mat_22_29_io_out_c_data;
  wire                pe_mat_22_29_io_out_c_is_weight;
  wire       [15:0]   pe_mat_22_30_io_out_r_data;
  wire                pe_mat_22_30_io_out_r_stop_weight;
  wire                pe_mat_22_30_io_out_r_stall;
  wire       [15:0]   pe_mat_22_30_io_out_c_data;
  wire                pe_mat_22_30_io_out_c_is_weight;
  wire       [15:0]   pe_mat_22_31_io_out_r_data;
  wire                pe_mat_22_31_io_out_r_stop_weight;
  wire                pe_mat_22_31_io_out_r_stall;
  wire       [15:0]   pe_mat_22_31_io_out_c_data;
  wire                pe_mat_22_31_io_out_c_is_weight;
  wire       [15:0]   pe_mat_23_0_io_out_r_data;
  wire                pe_mat_23_0_io_out_r_stop_weight;
  wire                pe_mat_23_0_io_out_r_stall;
  wire       [15:0]   pe_mat_23_0_io_out_c_data;
  wire                pe_mat_23_0_io_out_c_is_weight;
  wire       [15:0]   pe_mat_23_1_io_out_r_data;
  wire                pe_mat_23_1_io_out_r_stop_weight;
  wire                pe_mat_23_1_io_out_r_stall;
  wire       [15:0]   pe_mat_23_1_io_out_c_data;
  wire                pe_mat_23_1_io_out_c_is_weight;
  wire       [15:0]   pe_mat_23_2_io_out_r_data;
  wire                pe_mat_23_2_io_out_r_stop_weight;
  wire                pe_mat_23_2_io_out_r_stall;
  wire       [15:0]   pe_mat_23_2_io_out_c_data;
  wire                pe_mat_23_2_io_out_c_is_weight;
  wire       [15:0]   pe_mat_23_3_io_out_r_data;
  wire                pe_mat_23_3_io_out_r_stop_weight;
  wire                pe_mat_23_3_io_out_r_stall;
  wire       [15:0]   pe_mat_23_3_io_out_c_data;
  wire                pe_mat_23_3_io_out_c_is_weight;
  wire       [15:0]   pe_mat_23_4_io_out_r_data;
  wire                pe_mat_23_4_io_out_r_stop_weight;
  wire                pe_mat_23_4_io_out_r_stall;
  wire       [15:0]   pe_mat_23_4_io_out_c_data;
  wire                pe_mat_23_4_io_out_c_is_weight;
  wire       [15:0]   pe_mat_23_5_io_out_r_data;
  wire                pe_mat_23_5_io_out_r_stop_weight;
  wire                pe_mat_23_5_io_out_r_stall;
  wire       [15:0]   pe_mat_23_5_io_out_c_data;
  wire                pe_mat_23_5_io_out_c_is_weight;
  wire       [15:0]   pe_mat_23_6_io_out_r_data;
  wire                pe_mat_23_6_io_out_r_stop_weight;
  wire                pe_mat_23_6_io_out_r_stall;
  wire       [15:0]   pe_mat_23_6_io_out_c_data;
  wire                pe_mat_23_6_io_out_c_is_weight;
  wire       [15:0]   pe_mat_23_7_io_out_r_data;
  wire                pe_mat_23_7_io_out_r_stop_weight;
  wire                pe_mat_23_7_io_out_r_stall;
  wire       [15:0]   pe_mat_23_7_io_out_c_data;
  wire                pe_mat_23_7_io_out_c_is_weight;
  wire       [15:0]   pe_mat_23_8_io_out_r_data;
  wire                pe_mat_23_8_io_out_r_stop_weight;
  wire                pe_mat_23_8_io_out_r_stall;
  wire       [15:0]   pe_mat_23_8_io_out_c_data;
  wire                pe_mat_23_8_io_out_c_is_weight;
  wire       [15:0]   pe_mat_23_9_io_out_r_data;
  wire                pe_mat_23_9_io_out_r_stop_weight;
  wire                pe_mat_23_9_io_out_r_stall;
  wire       [15:0]   pe_mat_23_9_io_out_c_data;
  wire                pe_mat_23_9_io_out_c_is_weight;
  wire       [15:0]   pe_mat_23_10_io_out_r_data;
  wire                pe_mat_23_10_io_out_r_stop_weight;
  wire                pe_mat_23_10_io_out_r_stall;
  wire       [15:0]   pe_mat_23_10_io_out_c_data;
  wire                pe_mat_23_10_io_out_c_is_weight;
  wire       [15:0]   pe_mat_23_11_io_out_r_data;
  wire                pe_mat_23_11_io_out_r_stop_weight;
  wire                pe_mat_23_11_io_out_r_stall;
  wire       [15:0]   pe_mat_23_11_io_out_c_data;
  wire                pe_mat_23_11_io_out_c_is_weight;
  wire       [15:0]   pe_mat_23_12_io_out_r_data;
  wire                pe_mat_23_12_io_out_r_stop_weight;
  wire                pe_mat_23_12_io_out_r_stall;
  wire       [15:0]   pe_mat_23_12_io_out_c_data;
  wire                pe_mat_23_12_io_out_c_is_weight;
  wire       [15:0]   pe_mat_23_13_io_out_r_data;
  wire                pe_mat_23_13_io_out_r_stop_weight;
  wire                pe_mat_23_13_io_out_r_stall;
  wire       [15:0]   pe_mat_23_13_io_out_c_data;
  wire                pe_mat_23_13_io_out_c_is_weight;
  wire       [15:0]   pe_mat_23_14_io_out_r_data;
  wire                pe_mat_23_14_io_out_r_stop_weight;
  wire                pe_mat_23_14_io_out_r_stall;
  wire       [15:0]   pe_mat_23_14_io_out_c_data;
  wire                pe_mat_23_14_io_out_c_is_weight;
  wire       [15:0]   pe_mat_23_15_io_out_r_data;
  wire                pe_mat_23_15_io_out_r_stop_weight;
  wire                pe_mat_23_15_io_out_r_stall;
  wire       [15:0]   pe_mat_23_15_io_out_c_data;
  wire                pe_mat_23_15_io_out_c_is_weight;
  wire       [15:0]   pe_mat_23_16_io_out_r_data;
  wire                pe_mat_23_16_io_out_r_stop_weight;
  wire                pe_mat_23_16_io_out_r_stall;
  wire       [15:0]   pe_mat_23_16_io_out_c_data;
  wire                pe_mat_23_16_io_out_c_is_weight;
  wire       [15:0]   pe_mat_23_17_io_out_r_data;
  wire                pe_mat_23_17_io_out_r_stop_weight;
  wire                pe_mat_23_17_io_out_r_stall;
  wire       [15:0]   pe_mat_23_17_io_out_c_data;
  wire                pe_mat_23_17_io_out_c_is_weight;
  wire       [15:0]   pe_mat_23_18_io_out_r_data;
  wire                pe_mat_23_18_io_out_r_stop_weight;
  wire                pe_mat_23_18_io_out_r_stall;
  wire       [15:0]   pe_mat_23_18_io_out_c_data;
  wire                pe_mat_23_18_io_out_c_is_weight;
  wire       [15:0]   pe_mat_23_19_io_out_r_data;
  wire                pe_mat_23_19_io_out_r_stop_weight;
  wire                pe_mat_23_19_io_out_r_stall;
  wire       [15:0]   pe_mat_23_19_io_out_c_data;
  wire                pe_mat_23_19_io_out_c_is_weight;
  wire       [15:0]   pe_mat_23_20_io_out_r_data;
  wire                pe_mat_23_20_io_out_r_stop_weight;
  wire                pe_mat_23_20_io_out_r_stall;
  wire       [15:0]   pe_mat_23_20_io_out_c_data;
  wire                pe_mat_23_20_io_out_c_is_weight;
  wire       [15:0]   pe_mat_23_21_io_out_r_data;
  wire                pe_mat_23_21_io_out_r_stop_weight;
  wire                pe_mat_23_21_io_out_r_stall;
  wire       [15:0]   pe_mat_23_21_io_out_c_data;
  wire                pe_mat_23_21_io_out_c_is_weight;
  wire       [15:0]   pe_mat_23_22_io_out_r_data;
  wire                pe_mat_23_22_io_out_r_stop_weight;
  wire                pe_mat_23_22_io_out_r_stall;
  wire       [15:0]   pe_mat_23_22_io_out_c_data;
  wire                pe_mat_23_22_io_out_c_is_weight;
  wire       [15:0]   pe_mat_23_23_io_out_r_data;
  wire                pe_mat_23_23_io_out_r_stop_weight;
  wire                pe_mat_23_23_io_out_r_stall;
  wire       [15:0]   pe_mat_23_23_io_out_c_data;
  wire                pe_mat_23_23_io_out_c_is_weight;
  wire       [15:0]   pe_mat_23_24_io_out_r_data;
  wire                pe_mat_23_24_io_out_r_stop_weight;
  wire                pe_mat_23_24_io_out_r_stall;
  wire       [15:0]   pe_mat_23_24_io_out_c_data;
  wire                pe_mat_23_24_io_out_c_is_weight;
  wire       [15:0]   pe_mat_23_25_io_out_r_data;
  wire                pe_mat_23_25_io_out_r_stop_weight;
  wire                pe_mat_23_25_io_out_r_stall;
  wire       [15:0]   pe_mat_23_25_io_out_c_data;
  wire                pe_mat_23_25_io_out_c_is_weight;
  wire       [15:0]   pe_mat_23_26_io_out_r_data;
  wire                pe_mat_23_26_io_out_r_stop_weight;
  wire                pe_mat_23_26_io_out_r_stall;
  wire       [15:0]   pe_mat_23_26_io_out_c_data;
  wire                pe_mat_23_26_io_out_c_is_weight;
  wire       [15:0]   pe_mat_23_27_io_out_r_data;
  wire                pe_mat_23_27_io_out_r_stop_weight;
  wire                pe_mat_23_27_io_out_r_stall;
  wire       [15:0]   pe_mat_23_27_io_out_c_data;
  wire                pe_mat_23_27_io_out_c_is_weight;
  wire       [15:0]   pe_mat_23_28_io_out_r_data;
  wire                pe_mat_23_28_io_out_r_stop_weight;
  wire                pe_mat_23_28_io_out_r_stall;
  wire       [15:0]   pe_mat_23_28_io_out_c_data;
  wire                pe_mat_23_28_io_out_c_is_weight;
  wire       [15:0]   pe_mat_23_29_io_out_r_data;
  wire                pe_mat_23_29_io_out_r_stop_weight;
  wire                pe_mat_23_29_io_out_r_stall;
  wire       [15:0]   pe_mat_23_29_io_out_c_data;
  wire                pe_mat_23_29_io_out_c_is_weight;
  wire       [15:0]   pe_mat_23_30_io_out_r_data;
  wire                pe_mat_23_30_io_out_r_stop_weight;
  wire                pe_mat_23_30_io_out_r_stall;
  wire       [15:0]   pe_mat_23_30_io_out_c_data;
  wire                pe_mat_23_30_io_out_c_is_weight;
  wire       [15:0]   pe_mat_23_31_io_out_r_data;
  wire                pe_mat_23_31_io_out_r_stop_weight;
  wire                pe_mat_23_31_io_out_r_stall;
  wire       [15:0]   pe_mat_23_31_io_out_c_data;
  wire                pe_mat_23_31_io_out_c_is_weight;
  wire       [15:0]   pe_mat_24_0_io_out_r_data;
  wire                pe_mat_24_0_io_out_r_stop_weight;
  wire                pe_mat_24_0_io_out_r_stall;
  wire       [15:0]   pe_mat_24_0_io_out_c_data;
  wire                pe_mat_24_0_io_out_c_is_weight;
  wire       [15:0]   pe_mat_24_1_io_out_r_data;
  wire                pe_mat_24_1_io_out_r_stop_weight;
  wire                pe_mat_24_1_io_out_r_stall;
  wire       [15:0]   pe_mat_24_1_io_out_c_data;
  wire                pe_mat_24_1_io_out_c_is_weight;
  wire       [15:0]   pe_mat_24_2_io_out_r_data;
  wire                pe_mat_24_2_io_out_r_stop_weight;
  wire                pe_mat_24_2_io_out_r_stall;
  wire       [15:0]   pe_mat_24_2_io_out_c_data;
  wire                pe_mat_24_2_io_out_c_is_weight;
  wire       [15:0]   pe_mat_24_3_io_out_r_data;
  wire                pe_mat_24_3_io_out_r_stop_weight;
  wire                pe_mat_24_3_io_out_r_stall;
  wire       [15:0]   pe_mat_24_3_io_out_c_data;
  wire                pe_mat_24_3_io_out_c_is_weight;
  wire       [15:0]   pe_mat_24_4_io_out_r_data;
  wire                pe_mat_24_4_io_out_r_stop_weight;
  wire                pe_mat_24_4_io_out_r_stall;
  wire       [15:0]   pe_mat_24_4_io_out_c_data;
  wire                pe_mat_24_4_io_out_c_is_weight;
  wire       [15:0]   pe_mat_24_5_io_out_r_data;
  wire                pe_mat_24_5_io_out_r_stop_weight;
  wire                pe_mat_24_5_io_out_r_stall;
  wire       [15:0]   pe_mat_24_5_io_out_c_data;
  wire                pe_mat_24_5_io_out_c_is_weight;
  wire       [15:0]   pe_mat_24_6_io_out_r_data;
  wire                pe_mat_24_6_io_out_r_stop_weight;
  wire                pe_mat_24_6_io_out_r_stall;
  wire       [15:0]   pe_mat_24_6_io_out_c_data;
  wire                pe_mat_24_6_io_out_c_is_weight;
  wire       [15:0]   pe_mat_24_7_io_out_r_data;
  wire                pe_mat_24_7_io_out_r_stop_weight;
  wire                pe_mat_24_7_io_out_r_stall;
  wire       [15:0]   pe_mat_24_7_io_out_c_data;
  wire                pe_mat_24_7_io_out_c_is_weight;
  wire       [15:0]   pe_mat_24_8_io_out_r_data;
  wire                pe_mat_24_8_io_out_r_stop_weight;
  wire                pe_mat_24_8_io_out_r_stall;
  wire       [15:0]   pe_mat_24_8_io_out_c_data;
  wire                pe_mat_24_8_io_out_c_is_weight;
  wire       [15:0]   pe_mat_24_9_io_out_r_data;
  wire                pe_mat_24_9_io_out_r_stop_weight;
  wire                pe_mat_24_9_io_out_r_stall;
  wire       [15:0]   pe_mat_24_9_io_out_c_data;
  wire                pe_mat_24_9_io_out_c_is_weight;
  wire       [15:0]   pe_mat_24_10_io_out_r_data;
  wire                pe_mat_24_10_io_out_r_stop_weight;
  wire                pe_mat_24_10_io_out_r_stall;
  wire       [15:0]   pe_mat_24_10_io_out_c_data;
  wire                pe_mat_24_10_io_out_c_is_weight;
  wire       [15:0]   pe_mat_24_11_io_out_r_data;
  wire                pe_mat_24_11_io_out_r_stop_weight;
  wire                pe_mat_24_11_io_out_r_stall;
  wire       [15:0]   pe_mat_24_11_io_out_c_data;
  wire                pe_mat_24_11_io_out_c_is_weight;
  wire       [15:0]   pe_mat_24_12_io_out_r_data;
  wire                pe_mat_24_12_io_out_r_stop_weight;
  wire                pe_mat_24_12_io_out_r_stall;
  wire       [15:0]   pe_mat_24_12_io_out_c_data;
  wire                pe_mat_24_12_io_out_c_is_weight;
  wire       [15:0]   pe_mat_24_13_io_out_r_data;
  wire                pe_mat_24_13_io_out_r_stop_weight;
  wire                pe_mat_24_13_io_out_r_stall;
  wire       [15:0]   pe_mat_24_13_io_out_c_data;
  wire                pe_mat_24_13_io_out_c_is_weight;
  wire       [15:0]   pe_mat_24_14_io_out_r_data;
  wire                pe_mat_24_14_io_out_r_stop_weight;
  wire                pe_mat_24_14_io_out_r_stall;
  wire       [15:0]   pe_mat_24_14_io_out_c_data;
  wire                pe_mat_24_14_io_out_c_is_weight;
  wire       [15:0]   pe_mat_24_15_io_out_r_data;
  wire                pe_mat_24_15_io_out_r_stop_weight;
  wire                pe_mat_24_15_io_out_r_stall;
  wire       [15:0]   pe_mat_24_15_io_out_c_data;
  wire                pe_mat_24_15_io_out_c_is_weight;
  wire       [15:0]   pe_mat_24_16_io_out_r_data;
  wire                pe_mat_24_16_io_out_r_stop_weight;
  wire                pe_mat_24_16_io_out_r_stall;
  wire       [15:0]   pe_mat_24_16_io_out_c_data;
  wire                pe_mat_24_16_io_out_c_is_weight;
  wire       [15:0]   pe_mat_24_17_io_out_r_data;
  wire                pe_mat_24_17_io_out_r_stop_weight;
  wire                pe_mat_24_17_io_out_r_stall;
  wire       [15:0]   pe_mat_24_17_io_out_c_data;
  wire                pe_mat_24_17_io_out_c_is_weight;
  wire       [15:0]   pe_mat_24_18_io_out_r_data;
  wire                pe_mat_24_18_io_out_r_stop_weight;
  wire                pe_mat_24_18_io_out_r_stall;
  wire       [15:0]   pe_mat_24_18_io_out_c_data;
  wire                pe_mat_24_18_io_out_c_is_weight;
  wire       [15:0]   pe_mat_24_19_io_out_r_data;
  wire                pe_mat_24_19_io_out_r_stop_weight;
  wire                pe_mat_24_19_io_out_r_stall;
  wire       [15:0]   pe_mat_24_19_io_out_c_data;
  wire                pe_mat_24_19_io_out_c_is_weight;
  wire       [15:0]   pe_mat_24_20_io_out_r_data;
  wire                pe_mat_24_20_io_out_r_stop_weight;
  wire                pe_mat_24_20_io_out_r_stall;
  wire       [15:0]   pe_mat_24_20_io_out_c_data;
  wire                pe_mat_24_20_io_out_c_is_weight;
  wire       [15:0]   pe_mat_24_21_io_out_r_data;
  wire                pe_mat_24_21_io_out_r_stop_weight;
  wire                pe_mat_24_21_io_out_r_stall;
  wire       [15:0]   pe_mat_24_21_io_out_c_data;
  wire                pe_mat_24_21_io_out_c_is_weight;
  wire       [15:0]   pe_mat_24_22_io_out_r_data;
  wire                pe_mat_24_22_io_out_r_stop_weight;
  wire                pe_mat_24_22_io_out_r_stall;
  wire       [15:0]   pe_mat_24_22_io_out_c_data;
  wire                pe_mat_24_22_io_out_c_is_weight;
  wire       [15:0]   pe_mat_24_23_io_out_r_data;
  wire                pe_mat_24_23_io_out_r_stop_weight;
  wire                pe_mat_24_23_io_out_r_stall;
  wire       [15:0]   pe_mat_24_23_io_out_c_data;
  wire                pe_mat_24_23_io_out_c_is_weight;
  wire       [15:0]   pe_mat_24_24_io_out_r_data;
  wire                pe_mat_24_24_io_out_r_stop_weight;
  wire                pe_mat_24_24_io_out_r_stall;
  wire       [15:0]   pe_mat_24_24_io_out_c_data;
  wire                pe_mat_24_24_io_out_c_is_weight;
  wire       [15:0]   pe_mat_24_25_io_out_r_data;
  wire                pe_mat_24_25_io_out_r_stop_weight;
  wire                pe_mat_24_25_io_out_r_stall;
  wire       [15:0]   pe_mat_24_25_io_out_c_data;
  wire                pe_mat_24_25_io_out_c_is_weight;
  wire       [15:0]   pe_mat_24_26_io_out_r_data;
  wire                pe_mat_24_26_io_out_r_stop_weight;
  wire                pe_mat_24_26_io_out_r_stall;
  wire       [15:0]   pe_mat_24_26_io_out_c_data;
  wire                pe_mat_24_26_io_out_c_is_weight;
  wire       [15:0]   pe_mat_24_27_io_out_r_data;
  wire                pe_mat_24_27_io_out_r_stop_weight;
  wire                pe_mat_24_27_io_out_r_stall;
  wire       [15:0]   pe_mat_24_27_io_out_c_data;
  wire                pe_mat_24_27_io_out_c_is_weight;
  wire       [15:0]   pe_mat_24_28_io_out_r_data;
  wire                pe_mat_24_28_io_out_r_stop_weight;
  wire                pe_mat_24_28_io_out_r_stall;
  wire       [15:0]   pe_mat_24_28_io_out_c_data;
  wire                pe_mat_24_28_io_out_c_is_weight;
  wire       [15:0]   pe_mat_24_29_io_out_r_data;
  wire                pe_mat_24_29_io_out_r_stop_weight;
  wire                pe_mat_24_29_io_out_r_stall;
  wire       [15:0]   pe_mat_24_29_io_out_c_data;
  wire                pe_mat_24_29_io_out_c_is_weight;
  wire       [15:0]   pe_mat_24_30_io_out_r_data;
  wire                pe_mat_24_30_io_out_r_stop_weight;
  wire                pe_mat_24_30_io_out_r_stall;
  wire       [15:0]   pe_mat_24_30_io_out_c_data;
  wire                pe_mat_24_30_io_out_c_is_weight;
  wire       [15:0]   pe_mat_24_31_io_out_r_data;
  wire                pe_mat_24_31_io_out_r_stop_weight;
  wire                pe_mat_24_31_io_out_r_stall;
  wire       [15:0]   pe_mat_24_31_io_out_c_data;
  wire                pe_mat_24_31_io_out_c_is_weight;
  wire       [15:0]   pe_mat_25_0_io_out_r_data;
  wire                pe_mat_25_0_io_out_r_stop_weight;
  wire                pe_mat_25_0_io_out_r_stall;
  wire       [15:0]   pe_mat_25_0_io_out_c_data;
  wire                pe_mat_25_0_io_out_c_is_weight;
  wire       [15:0]   pe_mat_25_1_io_out_r_data;
  wire                pe_mat_25_1_io_out_r_stop_weight;
  wire                pe_mat_25_1_io_out_r_stall;
  wire       [15:0]   pe_mat_25_1_io_out_c_data;
  wire                pe_mat_25_1_io_out_c_is_weight;
  wire       [15:0]   pe_mat_25_2_io_out_r_data;
  wire                pe_mat_25_2_io_out_r_stop_weight;
  wire                pe_mat_25_2_io_out_r_stall;
  wire       [15:0]   pe_mat_25_2_io_out_c_data;
  wire                pe_mat_25_2_io_out_c_is_weight;
  wire       [15:0]   pe_mat_25_3_io_out_r_data;
  wire                pe_mat_25_3_io_out_r_stop_weight;
  wire                pe_mat_25_3_io_out_r_stall;
  wire       [15:0]   pe_mat_25_3_io_out_c_data;
  wire                pe_mat_25_3_io_out_c_is_weight;
  wire       [15:0]   pe_mat_25_4_io_out_r_data;
  wire                pe_mat_25_4_io_out_r_stop_weight;
  wire                pe_mat_25_4_io_out_r_stall;
  wire       [15:0]   pe_mat_25_4_io_out_c_data;
  wire                pe_mat_25_4_io_out_c_is_weight;
  wire       [15:0]   pe_mat_25_5_io_out_r_data;
  wire                pe_mat_25_5_io_out_r_stop_weight;
  wire                pe_mat_25_5_io_out_r_stall;
  wire       [15:0]   pe_mat_25_5_io_out_c_data;
  wire                pe_mat_25_5_io_out_c_is_weight;
  wire       [15:0]   pe_mat_25_6_io_out_r_data;
  wire                pe_mat_25_6_io_out_r_stop_weight;
  wire                pe_mat_25_6_io_out_r_stall;
  wire       [15:0]   pe_mat_25_6_io_out_c_data;
  wire                pe_mat_25_6_io_out_c_is_weight;
  wire       [15:0]   pe_mat_25_7_io_out_r_data;
  wire                pe_mat_25_7_io_out_r_stop_weight;
  wire                pe_mat_25_7_io_out_r_stall;
  wire       [15:0]   pe_mat_25_7_io_out_c_data;
  wire                pe_mat_25_7_io_out_c_is_weight;
  wire       [15:0]   pe_mat_25_8_io_out_r_data;
  wire                pe_mat_25_8_io_out_r_stop_weight;
  wire                pe_mat_25_8_io_out_r_stall;
  wire       [15:0]   pe_mat_25_8_io_out_c_data;
  wire                pe_mat_25_8_io_out_c_is_weight;
  wire       [15:0]   pe_mat_25_9_io_out_r_data;
  wire                pe_mat_25_9_io_out_r_stop_weight;
  wire                pe_mat_25_9_io_out_r_stall;
  wire       [15:0]   pe_mat_25_9_io_out_c_data;
  wire                pe_mat_25_9_io_out_c_is_weight;
  wire       [15:0]   pe_mat_25_10_io_out_r_data;
  wire                pe_mat_25_10_io_out_r_stop_weight;
  wire                pe_mat_25_10_io_out_r_stall;
  wire       [15:0]   pe_mat_25_10_io_out_c_data;
  wire                pe_mat_25_10_io_out_c_is_weight;
  wire       [15:0]   pe_mat_25_11_io_out_r_data;
  wire                pe_mat_25_11_io_out_r_stop_weight;
  wire                pe_mat_25_11_io_out_r_stall;
  wire       [15:0]   pe_mat_25_11_io_out_c_data;
  wire                pe_mat_25_11_io_out_c_is_weight;
  wire       [15:0]   pe_mat_25_12_io_out_r_data;
  wire                pe_mat_25_12_io_out_r_stop_weight;
  wire                pe_mat_25_12_io_out_r_stall;
  wire       [15:0]   pe_mat_25_12_io_out_c_data;
  wire                pe_mat_25_12_io_out_c_is_weight;
  wire       [15:0]   pe_mat_25_13_io_out_r_data;
  wire                pe_mat_25_13_io_out_r_stop_weight;
  wire                pe_mat_25_13_io_out_r_stall;
  wire       [15:0]   pe_mat_25_13_io_out_c_data;
  wire                pe_mat_25_13_io_out_c_is_weight;
  wire       [15:0]   pe_mat_25_14_io_out_r_data;
  wire                pe_mat_25_14_io_out_r_stop_weight;
  wire                pe_mat_25_14_io_out_r_stall;
  wire       [15:0]   pe_mat_25_14_io_out_c_data;
  wire                pe_mat_25_14_io_out_c_is_weight;
  wire       [15:0]   pe_mat_25_15_io_out_r_data;
  wire                pe_mat_25_15_io_out_r_stop_weight;
  wire                pe_mat_25_15_io_out_r_stall;
  wire       [15:0]   pe_mat_25_15_io_out_c_data;
  wire                pe_mat_25_15_io_out_c_is_weight;
  wire       [15:0]   pe_mat_25_16_io_out_r_data;
  wire                pe_mat_25_16_io_out_r_stop_weight;
  wire                pe_mat_25_16_io_out_r_stall;
  wire       [15:0]   pe_mat_25_16_io_out_c_data;
  wire                pe_mat_25_16_io_out_c_is_weight;
  wire       [15:0]   pe_mat_25_17_io_out_r_data;
  wire                pe_mat_25_17_io_out_r_stop_weight;
  wire                pe_mat_25_17_io_out_r_stall;
  wire       [15:0]   pe_mat_25_17_io_out_c_data;
  wire                pe_mat_25_17_io_out_c_is_weight;
  wire       [15:0]   pe_mat_25_18_io_out_r_data;
  wire                pe_mat_25_18_io_out_r_stop_weight;
  wire                pe_mat_25_18_io_out_r_stall;
  wire       [15:0]   pe_mat_25_18_io_out_c_data;
  wire                pe_mat_25_18_io_out_c_is_weight;
  wire       [15:0]   pe_mat_25_19_io_out_r_data;
  wire                pe_mat_25_19_io_out_r_stop_weight;
  wire                pe_mat_25_19_io_out_r_stall;
  wire       [15:0]   pe_mat_25_19_io_out_c_data;
  wire                pe_mat_25_19_io_out_c_is_weight;
  wire       [15:0]   pe_mat_25_20_io_out_r_data;
  wire                pe_mat_25_20_io_out_r_stop_weight;
  wire                pe_mat_25_20_io_out_r_stall;
  wire       [15:0]   pe_mat_25_20_io_out_c_data;
  wire                pe_mat_25_20_io_out_c_is_weight;
  wire       [15:0]   pe_mat_25_21_io_out_r_data;
  wire                pe_mat_25_21_io_out_r_stop_weight;
  wire                pe_mat_25_21_io_out_r_stall;
  wire       [15:0]   pe_mat_25_21_io_out_c_data;
  wire                pe_mat_25_21_io_out_c_is_weight;
  wire       [15:0]   pe_mat_25_22_io_out_r_data;
  wire                pe_mat_25_22_io_out_r_stop_weight;
  wire                pe_mat_25_22_io_out_r_stall;
  wire       [15:0]   pe_mat_25_22_io_out_c_data;
  wire                pe_mat_25_22_io_out_c_is_weight;
  wire       [15:0]   pe_mat_25_23_io_out_r_data;
  wire                pe_mat_25_23_io_out_r_stop_weight;
  wire                pe_mat_25_23_io_out_r_stall;
  wire       [15:0]   pe_mat_25_23_io_out_c_data;
  wire                pe_mat_25_23_io_out_c_is_weight;
  wire       [15:0]   pe_mat_25_24_io_out_r_data;
  wire                pe_mat_25_24_io_out_r_stop_weight;
  wire                pe_mat_25_24_io_out_r_stall;
  wire       [15:0]   pe_mat_25_24_io_out_c_data;
  wire                pe_mat_25_24_io_out_c_is_weight;
  wire       [15:0]   pe_mat_25_25_io_out_r_data;
  wire                pe_mat_25_25_io_out_r_stop_weight;
  wire                pe_mat_25_25_io_out_r_stall;
  wire       [15:0]   pe_mat_25_25_io_out_c_data;
  wire                pe_mat_25_25_io_out_c_is_weight;
  wire       [15:0]   pe_mat_25_26_io_out_r_data;
  wire                pe_mat_25_26_io_out_r_stop_weight;
  wire                pe_mat_25_26_io_out_r_stall;
  wire       [15:0]   pe_mat_25_26_io_out_c_data;
  wire                pe_mat_25_26_io_out_c_is_weight;
  wire       [15:0]   pe_mat_25_27_io_out_r_data;
  wire                pe_mat_25_27_io_out_r_stop_weight;
  wire                pe_mat_25_27_io_out_r_stall;
  wire       [15:0]   pe_mat_25_27_io_out_c_data;
  wire                pe_mat_25_27_io_out_c_is_weight;
  wire       [15:0]   pe_mat_25_28_io_out_r_data;
  wire                pe_mat_25_28_io_out_r_stop_weight;
  wire                pe_mat_25_28_io_out_r_stall;
  wire       [15:0]   pe_mat_25_28_io_out_c_data;
  wire                pe_mat_25_28_io_out_c_is_weight;
  wire       [15:0]   pe_mat_25_29_io_out_r_data;
  wire                pe_mat_25_29_io_out_r_stop_weight;
  wire                pe_mat_25_29_io_out_r_stall;
  wire       [15:0]   pe_mat_25_29_io_out_c_data;
  wire                pe_mat_25_29_io_out_c_is_weight;
  wire       [15:0]   pe_mat_25_30_io_out_r_data;
  wire                pe_mat_25_30_io_out_r_stop_weight;
  wire                pe_mat_25_30_io_out_r_stall;
  wire       [15:0]   pe_mat_25_30_io_out_c_data;
  wire                pe_mat_25_30_io_out_c_is_weight;
  wire       [15:0]   pe_mat_25_31_io_out_r_data;
  wire                pe_mat_25_31_io_out_r_stop_weight;
  wire                pe_mat_25_31_io_out_r_stall;
  wire       [15:0]   pe_mat_25_31_io_out_c_data;
  wire                pe_mat_25_31_io_out_c_is_weight;
  wire       [15:0]   pe_mat_26_0_io_out_r_data;
  wire                pe_mat_26_0_io_out_r_stop_weight;
  wire                pe_mat_26_0_io_out_r_stall;
  wire       [15:0]   pe_mat_26_0_io_out_c_data;
  wire                pe_mat_26_0_io_out_c_is_weight;
  wire       [15:0]   pe_mat_26_1_io_out_r_data;
  wire                pe_mat_26_1_io_out_r_stop_weight;
  wire                pe_mat_26_1_io_out_r_stall;
  wire       [15:0]   pe_mat_26_1_io_out_c_data;
  wire                pe_mat_26_1_io_out_c_is_weight;
  wire       [15:0]   pe_mat_26_2_io_out_r_data;
  wire                pe_mat_26_2_io_out_r_stop_weight;
  wire                pe_mat_26_2_io_out_r_stall;
  wire       [15:0]   pe_mat_26_2_io_out_c_data;
  wire                pe_mat_26_2_io_out_c_is_weight;
  wire       [15:0]   pe_mat_26_3_io_out_r_data;
  wire                pe_mat_26_3_io_out_r_stop_weight;
  wire                pe_mat_26_3_io_out_r_stall;
  wire       [15:0]   pe_mat_26_3_io_out_c_data;
  wire                pe_mat_26_3_io_out_c_is_weight;
  wire       [15:0]   pe_mat_26_4_io_out_r_data;
  wire                pe_mat_26_4_io_out_r_stop_weight;
  wire                pe_mat_26_4_io_out_r_stall;
  wire       [15:0]   pe_mat_26_4_io_out_c_data;
  wire                pe_mat_26_4_io_out_c_is_weight;
  wire       [15:0]   pe_mat_26_5_io_out_r_data;
  wire                pe_mat_26_5_io_out_r_stop_weight;
  wire                pe_mat_26_5_io_out_r_stall;
  wire       [15:0]   pe_mat_26_5_io_out_c_data;
  wire                pe_mat_26_5_io_out_c_is_weight;
  wire       [15:0]   pe_mat_26_6_io_out_r_data;
  wire                pe_mat_26_6_io_out_r_stop_weight;
  wire                pe_mat_26_6_io_out_r_stall;
  wire       [15:0]   pe_mat_26_6_io_out_c_data;
  wire                pe_mat_26_6_io_out_c_is_weight;
  wire       [15:0]   pe_mat_26_7_io_out_r_data;
  wire                pe_mat_26_7_io_out_r_stop_weight;
  wire                pe_mat_26_7_io_out_r_stall;
  wire       [15:0]   pe_mat_26_7_io_out_c_data;
  wire                pe_mat_26_7_io_out_c_is_weight;
  wire       [15:0]   pe_mat_26_8_io_out_r_data;
  wire                pe_mat_26_8_io_out_r_stop_weight;
  wire                pe_mat_26_8_io_out_r_stall;
  wire       [15:0]   pe_mat_26_8_io_out_c_data;
  wire                pe_mat_26_8_io_out_c_is_weight;
  wire       [15:0]   pe_mat_26_9_io_out_r_data;
  wire                pe_mat_26_9_io_out_r_stop_weight;
  wire                pe_mat_26_9_io_out_r_stall;
  wire       [15:0]   pe_mat_26_9_io_out_c_data;
  wire                pe_mat_26_9_io_out_c_is_weight;
  wire       [15:0]   pe_mat_26_10_io_out_r_data;
  wire                pe_mat_26_10_io_out_r_stop_weight;
  wire                pe_mat_26_10_io_out_r_stall;
  wire       [15:0]   pe_mat_26_10_io_out_c_data;
  wire                pe_mat_26_10_io_out_c_is_weight;
  wire       [15:0]   pe_mat_26_11_io_out_r_data;
  wire                pe_mat_26_11_io_out_r_stop_weight;
  wire                pe_mat_26_11_io_out_r_stall;
  wire       [15:0]   pe_mat_26_11_io_out_c_data;
  wire                pe_mat_26_11_io_out_c_is_weight;
  wire       [15:0]   pe_mat_26_12_io_out_r_data;
  wire                pe_mat_26_12_io_out_r_stop_weight;
  wire                pe_mat_26_12_io_out_r_stall;
  wire       [15:0]   pe_mat_26_12_io_out_c_data;
  wire                pe_mat_26_12_io_out_c_is_weight;
  wire       [15:0]   pe_mat_26_13_io_out_r_data;
  wire                pe_mat_26_13_io_out_r_stop_weight;
  wire                pe_mat_26_13_io_out_r_stall;
  wire       [15:0]   pe_mat_26_13_io_out_c_data;
  wire                pe_mat_26_13_io_out_c_is_weight;
  wire       [15:0]   pe_mat_26_14_io_out_r_data;
  wire                pe_mat_26_14_io_out_r_stop_weight;
  wire                pe_mat_26_14_io_out_r_stall;
  wire       [15:0]   pe_mat_26_14_io_out_c_data;
  wire                pe_mat_26_14_io_out_c_is_weight;
  wire       [15:0]   pe_mat_26_15_io_out_r_data;
  wire                pe_mat_26_15_io_out_r_stop_weight;
  wire                pe_mat_26_15_io_out_r_stall;
  wire       [15:0]   pe_mat_26_15_io_out_c_data;
  wire                pe_mat_26_15_io_out_c_is_weight;
  wire       [15:0]   pe_mat_26_16_io_out_r_data;
  wire                pe_mat_26_16_io_out_r_stop_weight;
  wire                pe_mat_26_16_io_out_r_stall;
  wire       [15:0]   pe_mat_26_16_io_out_c_data;
  wire                pe_mat_26_16_io_out_c_is_weight;
  wire       [15:0]   pe_mat_26_17_io_out_r_data;
  wire                pe_mat_26_17_io_out_r_stop_weight;
  wire                pe_mat_26_17_io_out_r_stall;
  wire       [15:0]   pe_mat_26_17_io_out_c_data;
  wire                pe_mat_26_17_io_out_c_is_weight;
  wire       [15:0]   pe_mat_26_18_io_out_r_data;
  wire                pe_mat_26_18_io_out_r_stop_weight;
  wire                pe_mat_26_18_io_out_r_stall;
  wire       [15:0]   pe_mat_26_18_io_out_c_data;
  wire                pe_mat_26_18_io_out_c_is_weight;
  wire       [15:0]   pe_mat_26_19_io_out_r_data;
  wire                pe_mat_26_19_io_out_r_stop_weight;
  wire                pe_mat_26_19_io_out_r_stall;
  wire       [15:0]   pe_mat_26_19_io_out_c_data;
  wire                pe_mat_26_19_io_out_c_is_weight;
  wire       [15:0]   pe_mat_26_20_io_out_r_data;
  wire                pe_mat_26_20_io_out_r_stop_weight;
  wire                pe_mat_26_20_io_out_r_stall;
  wire       [15:0]   pe_mat_26_20_io_out_c_data;
  wire                pe_mat_26_20_io_out_c_is_weight;
  wire       [15:0]   pe_mat_26_21_io_out_r_data;
  wire                pe_mat_26_21_io_out_r_stop_weight;
  wire                pe_mat_26_21_io_out_r_stall;
  wire       [15:0]   pe_mat_26_21_io_out_c_data;
  wire                pe_mat_26_21_io_out_c_is_weight;
  wire       [15:0]   pe_mat_26_22_io_out_r_data;
  wire                pe_mat_26_22_io_out_r_stop_weight;
  wire                pe_mat_26_22_io_out_r_stall;
  wire       [15:0]   pe_mat_26_22_io_out_c_data;
  wire                pe_mat_26_22_io_out_c_is_weight;
  wire       [15:0]   pe_mat_26_23_io_out_r_data;
  wire                pe_mat_26_23_io_out_r_stop_weight;
  wire                pe_mat_26_23_io_out_r_stall;
  wire       [15:0]   pe_mat_26_23_io_out_c_data;
  wire                pe_mat_26_23_io_out_c_is_weight;
  wire       [15:0]   pe_mat_26_24_io_out_r_data;
  wire                pe_mat_26_24_io_out_r_stop_weight;
  wire                pe_mat_26_24_io_out_r_stall;
  wire       [15:0]   pe_mat_26_24_io_out_c_data;
  wire                pe_mat_26_24_io_out_c_is_weight;
  wire       [15:0]   pe_mat_26_25_io_out_r_data;
  wire                pe_mat_26_25_io_out_r_stop_weight;
  wire                pe_mat_26_25_io_out_r_stall;
  wire       [15:0]   pe_mat_26_25_io_out_c_data;
  wire                pe_mat_26_25_io_out_c_is_weight;
  wire       [15:0]   pe_mat_26_26_io_out_r_data;
  wire                pe_mat_26_26_io_out_r_stop_weight;
  wire                pe_mat_26_26_io_out_r_stall;
  wire       [15:0]   pe_mat_26_26_io_out_c_data;
  wire                pe_mat_26_26_io_out_c_is_weight;
  wire       [15:0]   pe_mat_26_27_io_out_r_data;
  wire                pe_mat_26_27_io_out_r_stop_weight;
  wire                pe_mat_26_27_io_out_r_stall;
  wire       [15:0]   pe_mat_26_27_io_out_c_data;
  wire                pe_mat_26_27_io_out_c_is_weight;
  wire       [15:0]   pe_mat_26_28_io_out_r_data;
  wire                pe_mat_26_28_io_out_r_stop_weight;
  wire                pe_mat_26_28_io_out_r_stall;
  wire       [15:0]   pe_mat_26_28_io_out_c_data;
  wire                pe_mat_26_28_io_out_c_is_weight;
  wire       [15:0]   pe_mat_26_29_io_out_r_data;
  wire                pe_mat_26_29_io_out_r_stop_weight;
  wire                pe_mat_26_29_io_out_r_stall;
  wire       [15:0]   pe_mat_26_29_io_out_c_data;
  wire                pe_mat_26_29_io_out_c_is_weight;
  wire       [15:0]   pe_mat_26_30_io_out_r_data;
  wire                pe_mat_26_30_io_out_r_stop_weight;
  wire                pe_mat_26_30_io_out_r_stall;
  wire       [15:0]   pe_mat_26_30_io_out_c_data;
  wire                pe_mat_26_30_io_out_c_is_weight;
  wire       [15:0]   pe_mat_26_31_io_out_r_data;
  wire                pe_mat_26_31_io_out_r_stop_weight;
  wire                pe_mat_26_31_io_out_r_stall;
  wire       [15:0]   pe_mat_26_31_io_out_c_data;
  wire                pe_mat_26_31_io_out_c_is_weight;
  wire       [15:0]   pe_mat_27_0_io_out_r_data;
  wire                pe_mat_27_0_io_out_r_stop_weight;
  wire                pe_mat_27_0_io_out_r_stall;
  wire       [15:0]   pe_mat_27_0_io_out_c_data;
  wire                pe_mat_27_0_io_out_c_is_weight;
  wire       [15:0]   pe_mat_27_1_io_out_r_data;
  wire                pe_mat_27_1_io_out_r_stop_weight;
  wire                pe_mat_27_1_io_out_r_stall;
  wire       [15:0]   pe_mat_27_1_io_out_c_data;
  wire                pe_mat_27_1_io_out_c_is_weight;
  wire       [15:0]   pe_mat_27_2_io_out_r_data;
  wire                pe_mat_27_2_io_out_r_stop_weight;
  wire                pe_mat_27_2_io_out_r_stall;
  wire       [15:0]   pe_mat_27_2_io_out_c_data;
  wire                pe_mat_27_2_io_out_c_is_weight;
  wire       [15:0]   pe_mat_27_3_io_out_r_data;
  wire                pe_mat_27_3_io_out_r_stop_weight;
  wire                pe_mat_27_3_io_out_r_stall;
  wire       [15:0]   pe_mat_27_3_io_out_c_data;
  wire                pe_mat_27_3_io_out_c_is_weight;
  wire       [15:0]   pe_mat_27_4_io_out_r_data;
  wire                pe_mat_27_4_io_out_r_stop_weight;
  wire                pe_mat_27_4_io_out_r_stall;
  wire       [15:0]   pe_mat_27_4_io_out_c_data;
  wire                pe_mat_27_4_io_out_c_is_weight;
  wire       [15:0]   pe_mat_27_5_io_out_r_data;
  wire                pe_mat_27_5_io_out_r_stop_weight;
  wire                pe_mat_27_5_io_out_r_stall;
  wire       [15:0]   pe_mat_27_5_io_out_c_data;
  wire                pe_mat_27_5_io_out_c_is_weight;
  wire       [15:0]   pe_mat_27_6_io_out_r_data;
  wire                pe_mat_27_6_io_out_r_stop_weight;
  wire                pe_mat_27_6_io_out_r_stall;
  wire       [15:0]   pe_mat_27_6_io_out_c_data;
  wire                pe_mat_27_6_io_out_c_is_weight;
  wire       [15:0]   pe_mat_27_7_io_out_r_data;
  wire                pe_mat_27_7_io_out_r_stop_weight;
  wire                pe_mat_27_7_io_out_r_stall;
  wire       [15:0]   pe_mat_27_7_io_out_c_data;
  wire                pe_mat_27_7_io_out_c_is_weight;
  wire       [15:0]   pe_mat_27_8_io_out_r_data;
  wire                pe_mat_27_8_io_out_r_stop_weight;
  wire                pe_mat_27_8_io_out_r_stall;
  wire       [15:0]   pe_mat_27_8_io_out_c_data;
  wire                pe_mat_27_8_io_out_c_is_weight;
  wire       [15:0]   pe_mat_27_9_io_out_r_data;
  wire                pe_mat_27_9_io_out_r_stop_weight;
  wire                pe_mat_27_9_io_out_r_stall;
  wire       [15:0]   pe_mat_27_9_io_out_c_data;
  wire                pe_mat_27_9_io_out_c_is_weight;
  wire       [15:0]   pe_mat_27_10_io_out_r_data;
  wire                pe_mat_27_10_io_out_r_stop_weight;
  wire                pe_mat_27_10_io_out_r_stall;
  wire       [15:0]   pe_mat_27_10_io_out_c_data;
  wire                pe_mat_27_10_io_out_c_is_weight;
  wire       [15:0]   pe_mat_27_11_io_out_r_data;
  wire                pe_mat_27_11_io_out_r_stop_weight;
  wire                pe_mat_27_11_io_out_r_stall;
  wire       [15:0]   pe_mat_27_11_io_out_c_data;
  wire                pe_mat_27_11_io_out_c_is_weight;
  wire       [15:0]   pe_mat_27_12_io_out_r_data;
  wire                pe_mat_27_12_io_out_r_stop_weight;
  wire                pe_mat_27_12_io_out_r_stall;
  wire       [15:0]   pe_mat_27_12_io_out_c_data;
  wire                pe_mat_27_12_io_out_c_is_weight;
  wire       [15:0]   pe_mat_27_13_io_out_r_data;
  wire                pe_mat_27_13_io_out_r_stop_weight;
  wire                pe_mat_27_13_io_out_r_stall;
  wire       [15:0]   pe_mat_27_13_io_out_c_data;
  wire                pe_mat_27_13_io_out_c_is_weight;
  wire       [15:0]   pe_mat_27_14_io_out_r_data;
  wire                pe_mat_27_14_io_out_r_stop_weight;
  wire                pe_mat_27_14_io_out_r_stall;
  wire       [15:0]   pe_mat_27_14_io_out_c_data;
  wire                pe_mat_27_14_io_out_c_is_weight;
  wire       [15:0]   pe_mat_27_15_io_out_r_data;
  wire                pe_mat_27_15_io_out_r_stop_weight;
  wire                pe_mat_27_15_io_out_r_stall;
  wire       [15:0]   pe_mat_27_15_io_out_c_data;
  wire                pe_mat_27_15_io_out_c_is_weight;
  wire       [15:0]   pe_mat_27_16_io_out_r_data;
  wire                pe_mat_27_16_io_out_r_stop_weight;
  wire                pe_mat_27_16_io_out_r_stall;
  wire       [15:0]   pe_mat_27_16_io_out_c_data;
  wire                pe_mat_27_16_io_out_c_is_weight;
  wire       [15:0]   pe_mat_27_17_io_out_r_data;
  wire                pe_mat_27_17_io_out_r_stop_weight;
  wire                pe_mat_27_17_io_out_r_stall;
  wire       [15:0]   pe_mat_27_17_io_out_c_data;
  wire                pe_mat_27_17_io_out_c_is_weight;
  wire       [15:0]   pe_mat_27_18_io_out_r_data;
  wire                pe_mat_27_18_io_out_r_stop_weight;
  wire                pe_mat_27_18_io_out_r_stall;
  wire       [15:0]   pe_mat_27_18_io_out_c_data;
  wire                pe_mat_27_18_io_out_c_is_weight;
  wire       [15:0]   pe_mat_27_19_io_out_r_data;
  wire                pe_mat_27_19_io_out_r_stop_weight;
  wire                pe_mat_27_19_io_out_r_stall;
  wire       [15:0]   pe_mat_27_19_io_out_c_data;
  wire                pe_mat_27_19_io_out_c_is_weight;
  wire       [15:0]   pe_mat_27_20_io_out_r_data;
  wire                pe_mat_27_20_io_out_r_stop_weight;
  wire                pe_mat_27_20_io_out_r_stall;
  wire       [15:0]   pe_mat_27_20_io_out_c_data;
  wire                pe_mat_27_20_io_out_c_is_weight;
  wire       [15:0]   pe_mat_27_21_io_out_r_data;
  wire                pe_mat_27_21_io_out_r_stop_weight;
  wire                pe_mat_27_21_io_out_r_stall;
  wire       [15:0]   pe_mat_27_21_io_out_c_data;
  wire                pe_mat_27_21_io_out_c_is_weight;
  wire       [15:0]   pe_mat_27_22_io_out_r_data;
  wire                pe_mat_27_22_io_out_r_stop_weight;
  wire                pe_mat_27_22_io_out_r_stall;
  wire       [15:0]   pe_mat_27_22_io_out_c_data;
  wire                pe_mat_27_22_io_out_c_is_weight;
  wire       [15:0]   pe_mat_27_23_io_out_r_data;
  wire                pe_mat_27_23_io_out_r_stop_weight;
  wire                pe_mat_27_23_io_out_r_stall;
  wire       [15:0]   pe_mat_27_23_io_out_c_data;
  wire                pe_mat_27_23_io_out_c_is_weight;
  wire       [15:0]   pe_mat_27_24_io_out_r_data;
  wire                pe_mat_27_24_io_out_r_stop_weight;
  wire                pe_mat_27_24_io_out_r_stall;
  wire       [15:0]   pe_mat_27_24_io_out_c_data;
  wire                pe_mat_27_24_io_out_c_is_weight;
  wire       [15:0]   pe_mat_27_25_io_out_r_data;
  wire                pe_mat_27_25_io_out_r_stop_weight;
  wire                pe_mat_27_25_io_out_r_stall;
  wire       [15:0]   pe_mat_27_25_io_out_c_data;
  wire                pe_mat_27_25_io_out_c_is_weight;
  wire       [15:0]   pe_mat_27_26_io_out_r_data;
  wire                pe_mat_27_26_io_out_r_stop_weight;
  wire                pe_mat_27_26_io_out_r_stall;
  wire       [15:0]   pe_mat_27_26_io_out_c_data;
  wire                pe_mat_27_26_io_out_c_is_weight;
  wire       [15:0]   pe_mat_27_27_io_out_r_data;
  wire                pe_mat_27_27_io_out_r_stop_weight;
  wire                pe_mat_27_27_io_out_r_stall;
  wire       [15:0]   pe_mat_27_27_io_out_c_data;
  wire                pe_mat_27_27_io_out_c_is_weight;
  wire       [15:0]   pe_mat_27_28_io_out_r_data;
  wire                pe_mat_27_28_io_out_r_stop_weight;
  wire                pe_mat_27_28_io_out_r_stall;
  wire       [15:0]   pe_mat_27_28_io_out_c_data;
  wire                pe_mat_27_28_io_out_c_is_weight;
  wire       [15:0]   pe_mat_27_29_io_out_r_data;
  wire                pe_mat_27_29_io_out_r_stop_weight;
  wire                pe_mat_27_29_io_out_r_stall;
  wire       [15:0]   pe_mat_27_29_io_out_c_data;
  wire                pe_mat_27_29_io_out_c_is_weight;
  wire       [15:0]   pe_mat_27_30_io_out_r_data;
  wire                pe_mat_27_30_io_out_r_stop_weight;
  wire                pe_mat_27_30_io_out_r_stall;
  wire       [15:0]   pe_mat_27_30_io_out_c_data;
  wire                pe_mat_27_30_io_out_c_is_weight;
  wire       [15:0]   pe_mat_27_31_io_out_r_data;
  wire                pe_mat_27_31_io_out_r_stop_weight;
  wire                pe_mat_27_31_io_out_r_stall;
  wire       [15:0]   pe_mat_27_31_io_out_c_data;
  wire                pe_mat_27_31_io_out_c_is_weight;
  wire       [15:0]   pe_mat_28_0_io_out_r_data;
  wire                pe_mat_28_0_io_out_r_stop_weight;
  wire                pe_mat_28_0_io_out_r_stall;
  wire       [15:0]   pe_mat_28_0_io_out_c_data;
  wire                pe_mat_28_0_io_out_c_is_weight;
  wire       [15:0]   pe_mat_28_1_io_out_r_data;
  wire                pe_mat_28_1_io_out_r_stop_weight;
  wire                pe_mat_28_1_io_out_r_stall;
  wire       [15:0]   pe_mat_28_1_io_out_c_data;
  wire                pe_mat_28_1_io_out_c_is_weight;
  wire       [15:0]   pe_mat_28_2_io_out_r_data;
  wire                pe_mat_28_2_io_out_r_stop_weight;
  wire                pe_mat_28_2_io_out_r_stall;
  wire       [15:0]   pe_mat_28_2_io_out_c_data;
  wire                pe_mat_28_2_io_out_c_is_weight;
  wire       [15:0]   pe_mat_28_3_io_out_r_data;
  wire                pe_mat_28_3_io_out_r_stop_weight;
  wire                pe_mat_28_3_io_out_r_stall;
  wire       [15:0]   pe_mat_28_3_io_out_c_data;
  wire                pe_mat_28_3_io_out_c_is_weight;
  wire       [15:0]   pe_mat_28_4_io_out_r_data;
  wire                pe_mat_28_4_io_out_r_stop_weight;
  wire                pe_mat_28_4_io_out_r_stall;
  wire       [15:0]   pe_mat_28_4_io_out_c_data;
  wire                pe_mat_28_4_io_out_c_is_weight;
  wire       [15:0]   pe_mat_28_5_io_out_r_data;
  wire                pe_mat_28_5_io_out_r_stop_weight;
  wire                pe_mat_28_5_io_out_r_stall;
  wire       [15:0]   pe_mat_28_5_io_out_c_data;
  wire                pe_mat_28_5_io_out_c_is_weight;
  wire       [15:0]   pe_mat_28_6_io_out_r_data;
  wire                pe_mat_28_6_io_out_r_stop_weight;
  wire                pe_mat_28_6_io_out_r_stall;
  wire       [15:0]   pe_mat_28_6_io_out_c_data;
  wire                pe_mat_28_6_io_out_c_is_weight;
  wire       [15:0]   pe_mat_28_7_io_out_r_data;
  wire                pe_mat_28_7_io_out_r_stop_weight;
  wire                pe_mat_28_7_io_out_r_stall;
  wire       [15:0]   pe_mat_28_7_io_out_c_data;
  wire                pe_mat_28_7_io_out_c_is_weight;
  wire       [15:0]   pe_mat_28_8_io_out_r_data;
  wire                pe_mat_28_8_io_out_r_stop_weight;
  wire                pe_mat_28_8_io_out_r_stall;
  wire       [15:0]   pe_mat_28_8_io_out_c_data;
  wire                pe_mat_28_8_io_out_c_is_weight;
  wire       [15:0]   pe_mat_28_9_io_out_r_data;
  wire                pe_mat_28_9_io_out_r_stop_weight;
  wire                pe_mat_28_9_io_out_r_stall;
  wire       [15:0]   pe_mat_28_9_io_out_c_data;
  wire                pe_mat_28_9_io_out_c_is_weight;
  wire       [15:0]   pe_mat_28_10_io_out_r_data;
  wire                pe_mat_28_10_io_out_r_stop_weight;
  wire                pe_mat_28_10_io_out_r_stall;
  wire       [15:0]   pe_mat_28_10_io_out_c_data;
  wire                pe_mat_28_10_io_out_c_is_weight;
  wire       [15:0]   pe_mat_28_11_io_out_r_data;
  wire                pe_mat_28_11_io_out_r_stop_weight;
  wire                pe_mat_28_11_io_out_r_stall;
  wire       [15:0]   pe_mat_28_11_io_out_c_data;
  wire                pe_mat_28_11_io_out_c_is_weight;
  wire       [15:0]   pe_mat_28_12_io_out_r_data;
  wire                pe_mat_28_12_io_out_r_stop_weight;
  wire                pe_mat_28_12_io_out_r_stall;
  wire       [15:0]   pe_mat_28_12_io_out_c_data;
  wire                pe_mat_28_12_io_out_c_is_weight;
  wire       [15:0]   pe_mat_28_13_io_out_r_data;
  wire                pe_mat_28_13_io_out_r_stop_weight;
  wire                pe_mat_28_13_io_out_r_stall;
  wire       [15:0]   pe_mat_28_13_io_out_c_data;
  wire                pe_mat_28_13_io_out_c_is_weight;
  wire       [15:0]   pe_mat_28_14_io_out_r_data;
  wire                pe_mat_28_14_io_out_r_stop_weight;
  wire                pe_mat_28_14_io_out_r_stall;
  wire       [15:0]   pe_mat_28_14_io_out_c_data;
  wire                pe_mat_28_14_io_out_c_is_weight;
  wire       [15:0]   pe_mat_28_15_io_out_r_data;
  wire                pe_mat_28_15_io_out_r_stop_weight;
  wire                pe_mat_28_15_io_out_r_stall;
  wire       [15:0]   pe_mat_28_15_io_out_c_data;
  wire                pe_mat_28_15_io_out_c_is_weight;
  wire       [15:0]   pe_mat_28_16_io_out_r_data;
  wire                pe_mat_28_16_io_out_r_stop_weight;
  wire                pe_mat_28_16_io_out_r_stall;
  wire       [15:0]   pe_mat_28_16_io_out_c_data;
  wire                pe_mat_28_16_io_out_c_is_weight;
  wire       [15:0]   pe_mat_28_17_io_out_r_data;
  wire                pe_mat_28_17_io_out_r_stop_weight;
  wire                pe_mat_28_17_io_out_r_stall;
  wire       [15:0]   pe_mat_28_17_io_out_c_data;
  wire                pe_mat_28_17_io_out_c_is_weight;
  wire       [15:0]   pe_mat_28_18_io_out_r_data;
  wire                pe_mat_28_18_io_out_r_stop_weight;
  wire                pe_mat_28_18_io_out_r_stall;
  wire       [15:0]   pe_mat_28_18_io_out_c_data;
  wire                pe_mat_28_18_io_out_c_is_weight;
  wire       [15:0]   pe_mat_28_19_io_out_r_data;
  wire                pe_mat_28_19_io_out_r_stop_weight;
  wire                pe_mat_28_19_io_out_r_stall;
  wire       [15:0]   pe_mat_28_19_io_out_c_data;
  wire                pe_mat_28_19_io_out_c_is_weight;
  wire       [15:0]   pe_mat_28_20_io_out_r_data;
  wire                pe_mat_28_20_io_out_r_stop_weight;
  wire                pe_mat_28_20_io_out_r_stall;
  wire       [15:0]   pe_mat_28_20_io_out_c_data;
  wire                pe_mat_28_20_io_out_c_is_weight;
  wire       [15:0]   pe_mat_28_21_io_out_r_data;
  wire                pe_mat_28_21_io_out_r_stop_weight;
  wire                pe_mat_28_21_io_out_r_stall;
  wire       [15:0]   pe_mat_28_21_io_out_c_data;
  wire                pe_mat_28_21_io_out_c_is_weight;
  wire       [15:0]   pe_mat_28_22_io_out_r_data;
  wire                pe_mat_28_22_io_out_r_stop_weight;
  wire                pe_mat_28_22_io_out_r_stall;
  wire       [15:0]   pe_mat_28_22_io_out_c_data;
  wire                pe_mat_28_22_io_out_c_is_weight;
  wire       [15:0]   pe_mat_28_23_io_out_r_data;
  wire                pe_mat_28_23_io_out_r_stop_weight;
  wire                pe_mat_28_23_io_out_r_stall;
  wire       [15:0]   pe_mat_28_23_io_out_c_data;
  wire                pe_mat_28_23_io_out_c_is_weight;
  wire       [15:0]   pe_mat_28_24_io_out_r_data;
  wire                pe_mat_28_24_io_out_r_stop_weight;
  wire                pe_mat_28_24_io_out_r_stall;
  wire       [15:0]   pe_mat_28_24_io_out_c_data;
  wire                pe_mat_28_24_io_out_c_is_weight;
  wire       [15:0]   pe_mat_28_25_io_out_r_data;
  wire                pe_mat_28_25_io_out_r_stop_weight;
  wire                pe_mat_28_25_io_out_r_stall;
  wire       [15:0]   pe_mat_28_25_io_out_c_data;
  wire                pe_mat_28_25_io_out_c_is_weight;
  wire       [15:0]   pe_mat_28_26_io_out_r_data;
  wire                pe_mat_28_26_io_out_r_stop_weight;
  wire                pe_mat_28_26_io_out_r_stall;
  wire       [15:0]   pe_mat_28_26_io_out_c_data;
  wire                pe_mat_28_26_io_out_c_is_weight;
  wire       [15:0]   pe_mat_28_27_io_out_r_data;
  wire                pe_mat_28_27_io_out_r_stop_weight;
  wire                pe_mat_28_27_io_out_r_stall;
  wire       [15:0]   pe_mat_28_27_io_out_c_data;
  wire                pe_mat_28_27_io_out_c_is_weight;
  wire       [15:0]   pe_mat_28_28_io_out_r_data;
  wire                pe_mat_28_28_io_out_r_stop_weight;
  wire                pe_mat_28_28_io_out_r_stall;
  wire       [15:0]   pe_mat_28_28_io_out_c_data;
  wire                pe_mat_28_28_io_out_c_is_weight;
  wire       [15:0]   pe_mat_28_29_io_out_r_data;
  wire                pe_mat_28_29_io_out_r_stop_weight;
  wire                pe_mat_28_29_io_out_r_stall;
  wire       [15:0]   pe_mat_28_29_io_out_c_data;
  wire                pe_mat_28_29_io_out_c_is_weight;
  wire       [15:0]   pe_mat_28_30_io_out_r_data;
  wire                pe_mat_28_30_io_out_r_stop_weight;
  wire                pe_mat_28_30_io_out_r_stall;
  wire       [15:0]   pe_mat_28_30_io_out_c_data;
  wire                pe_mat_28_30_io_out_c_is_weight;
  wire       [15:0]   pe_mat_28_31_io_out_r_data;
  wire                pe_mat_28_31_io_out_r_stop_weight;
  wire                pe_mat_28_31_io_out_r_stall;
  wire       [15:0]   pe_mat_28_31_io_out_c_data;
  wire                pe_mat_28_31_io_out_c_is_weight;
  wire       [15:0]   pe_mat_29_0_io_out_r_data;
  wire                pe_mat_29_0_io_out_r_stop_weight;
  wire                pe_mat_29_0_io_out_r_stall;
  wire       [15:0]   pe_mat_29_0_io_out_c_data;
  wire                pe_mat_29_0_io_out_c_is_weight;
  wire       [15:0]   pe_mat_29_1_io_out_r_data;
  wire                pe_mat_29_1_io_out_r_stop_weight;
  wire                pe_mat_29_1_io_out_r_stall;
  wire       [15:0]   pe_mat_29_1_io_out_c_data;
  wire                pe_mat_29_1_io_out_c_is_weight;
  wire       [15:0]   pe_mat_29_2_io_out_r_data;
  wire                pe_mat_29_2_io_out_r_stop_weight;
  wire                pe_mat_29_2_io_out_r_stall;
  wire       [15:0]   pe_mat_29_2_io_out_c_data;
  wire                pe_mat_29_2_io_out_c_is_weight;
  wire       [15:0]   pe_mat_29_3_io_out_r_data;
  wire                pe_mat_29_3_io_out_r_stop_weight;
  wire                pe_mat_29_3_io_out_r_stall;
  wire       [15:0]   pe_mat_29_3_io_out_c_data;
  wire                pe_mat_29_3_io_out_c_is_weight;
  wire       [15:0]   pe_mat_29_4_io_out_r_data;
  wire                pe_mat_29_4_io_out_r_stop_weight;
  wire                pe_mat_29_4_io_out_r_stall;
  wire       [15:0]   pe_mat_29_4_io_out_c_data;
  wire                pe_mat_29_4_io_out_c_is_weight;
  wire       [15:0]   pe_mat_29_5_io_out_r_data;
  wire                pe_mat_29_5_io_out_r_stop_weight;
  wire                pe_mat_29_5_io_out_r_stall;
  wire       [15:0]   pe_mat_29_5_io_out_c_data;
  wire                pe_mat_29_5_io_out_c_is_weight;
  wire       [15:0]   pe_mat_29_6_io_out_r_data;
  wire                pe_mat_29_6_io_out_r_stop_weight;
  wire                pe_mat_29_6_io_out_r_stall;
  wire       [15:0]   pe_mat_29_6_io_out_c_data;
  wire                pe_mat_29_6_io_out_c_is_weight;
  wire       [15:0]   pe_mat_29_7_io_out_r_data;
  wire                pe_mat_29_7_io_out_r_stop_weight;
  wire                pe_mat_29_7_io_out_r_stall;
  wire       [15:0]   pe_mat_29_7_io_out_c_data;
  wire                pe_mat_29_7_io_out_c_is_weight;
  wire       [15:0]   pe_mat_29_8_io_out_r_data;
  wire                pe_mat_29_8_io_out_r_stop_weight;
  wire                pe_mat_29_8_io_out_r_stall;
  wire       [15:0]   pe_mat_29_8_io_out_c_data;
  wire                pe_mat_29_8_io_out_c_is_weight;
  wire       [15:0]   pe_mat_29_9_io_out_r_data;
  wire                pe_mat_29_9_io_out_r_stop_weight;
  wire                pe_mat_29_9_io_out_r_stall;
  wire       [15:0]   pe_mat_29_9_io_out_c_data;
  wire                pe_mat_29_9_io_out_c_is_weight;
  wire       [15:0]   pe_mat_29_10_io_out_r_data;
  wire                pe_mat_29_10_io_out_r_stop_weight;
  wire                pe_mat_29_10_io_out_r_stall;
  wire       [15:0]   pe_mat_29_10_io_out_c_data;
  wire                pe_mat_29_10_io_out_c_is_weight;
  wire       [15:0]   pe_mat_29_11_io_out_r_data;
  wire                pe_mat_29_11_io_out_r_stop_weight;
  wire                pe_mat_29_11_io_out_r_stall;
  wire       [15:0]   pe_mat_29_11_io_out_c_data;
  wire                pe_mat_29_11_io_out_c_is_weight;
  wire       [15:0]   pe_mat_29_12_io_out_r_data;
  wire                pe_mat_29_12_io_out_r_stop_weight;
  wire                pe_mat_29_12_io_out_r_stall;
  wire       [15:0]   pe_mat_29_12_io_out_c_data;
  wire                pe_mat_29_12_io_out_c_is_weight;
  wire       [15:0]   pe_mat_29_13_io_out_r_data;
  wire                pe_mat_29_13_io_out_r_stop_weight;
  wire                pe_mat_29_13_io_out_r_stall;
  wire       [15:0]   pe_mat_29_13_io_out_c_data;
  wire                pe_mat_29_13_io_out_c_is_weight;
  wire       [15:0]   pe_mat_29_14_io_out_r_data;
  wire                pe_mat_29_14_io_out_r_stop_weight;
  wire                pe_mat_29_14_io_out_r_stall;
  wire       [15:0]   pe_mat_29_14_io_out_c_data;
  wire                pe_mat_29_14_io_out_c_is_weight;
  wire       [15:0]   pe_mat_29_15_io_out_r_data;
  wire                pe_mat_29_15_io_out_r_stop_weight;
  wire                pe_mat_29_15_io_out_r_stall;
  wire       [15:0]   pe_mat_29_15_io_out_c_data;
  wire                pe_mat_29_15_io_out_c_is_weight;
  wire       [15:0]   pe_mat_29_16_io_out_r_data;
  wire                pe_mat_29_16_io_out_r_stop_weight;
  wire                pe_mat_29_16_io_out_r_stall;
  wire       [15:0]   pe_mat_29_16_io_out_c_data;
  wire                pe_mat_29_16_io_out_c_is_weight;
  wire       [15:0]   pe_mat_29_17_io_out_r_data;
  wire                pe_mat_29_17_io_out_r_stop_weight;
  wire                pe_mat_29_17_io_out_r_stall;
  wire       [15:0]   pe_mat_29_17_io_out_c_data;
  wire                pe_mat_29_17_io_out_c_is_weight;
  wire       [15:0]   pe_mat_29_18_io_out_r_data;
  wire                pe_mat_29_18_io_out_r_stop_weight;
  wire                pe_mat_29_18_io_out_r_stall;
  wire       [15:0]   pe_mat_29_18_io_out_c_data;
  wire                pe_mat_29_18_io_out_c_is_weight;
  wire       [15:0]   pe_mat_29_19_io_out_r_data;
  wire                pe_mat_29_19_io_out_r_stop_weight;
  wire                pe_mat_29_19_io_out_r_stall;
  wire       [15:0]   pe_mat_29_19_io_out_c_data;
  wire                pe_mat_29_19_io_out_c_is_weight;
  wire       [15:0]   pe_mat_29_20_io_out_r_data;
  wire                pe_mat_29_20_io_out_r_stop_weight;
  wire                pe_mat_29_20_io_out_r_stall;
  wire       [15:0]   pe_mat_29_20_io_out_c_data;
  wire                pe_mat_29_20_io_out_c_is_weight;
  wire       [15:0]   pe_mat_29_21_io_out_r_data;
  wire                pe_mat_29_21_io_out_r_stop_weight;
  wire                pe_mat_29_21_io_out_r_stall;
  wire       [15:0]   pe_mat_29_21_io_out_c_data;
  wire                pe_mat_29_21_io_out_c_is_weight;
  wire       [15:0]   pe_mat_29_22_io_out_r_data;
  wire                pe_mat_29_22_io_out_r_stop_weight;
  wire                pe_mat_29_22_io_out_r_stall;
  wire       [15:0]   pe_mat_29_22_io_out_c_data;
  wire                pe_mat_29_22_io_out_c_is_weight;
  wire       [15:0]   pe_mat_29_23_io_out_r_data;
  wire                pe_mat_29_23_io_out_r_stop_weight;
  wire                pe_mat_29_23_io_out_r_stall;
  wire       [15:0]   pe_mat_29_23_io_out_c_data;
  wire                pe_mat_29_23_io_out_c_is_weight;
  wire       [15:0]   pe_mat_29_24_io_out_r_data;
  wire                pe_mat_29_24_io_out_r_stop_weight;
  wire                pe_mat_29_24_io_out_r_stall;
  wire       [15:0]   pe_mat_29_24_io_out_c_data;
  wire                pe_mat_29_24_io_out_c_is_weight;
  wire       [15:0]   pe_mat_29_25_io_out_r_data;
  wire                pe_mat_29_25_io_out_r_stop_weight;
  wire                pe_mat_29_25_io_out_r_stall;
  wire       [15:0]   pe_mat_29_25_io_out_c_data;
  wire                pe_mat_29_25_io_out_c_is_weight;
  wire       [15:0]   pe_mat_29_26_io_out_r_data;
  wire                pe_mat_29_26_io_out_r_stop_weight;
  wire                pe_mat_29_26_io_out_r_stall;
  wire       [15:0]   pe_mat_29_26_io_out_c_data;
  wire                pe_mat_29_26_io_out_c_is_weight;
  wire       [15:0]   pe_mat_29_27_io_out_r_data;
  wire                pe_mat_29_27_io_out_r_stop_weight;
  wire                pe_mat_29_27_io_out_r_stall;
  wire       [15:0]   pe_mat_29_27_io_out_c_data;
  wire                pe_mat_29_27_io_out_c_is_weight;
  wire       [15:0]   pe_mat_29_28_io_out_r_data;
  wire                pe_mat_29_28_io_out_r_stop_weight;
  wire                pe_mat_29_28_io_out_r_stall;
  wire       [15:0]   pe_mat_29_28_io_out_c_data;
  wire                pe_mat_29_28_io_out_c_is_weight;
  wire       [15:0]   pe_mat_29_29_io_out_r_data;
  wire                pe_mat_29_29_io_out_r_stop_weight;
  wire                pe_mat_29_29_io_out_r_stall;
  wire       [15:0]   pe_mat_29_29_io_out_c_data;
  wire                pe_mat_29_29_io_out_c_is_weight;
  wire       [15:0]   pe_mat_29_30_io_out_r_data;
  wire                pe_mat_29_30_io_out_r_stop_weight;
  wire                pe_mat_29_30_io_out_r_stall;
  wire       [15:0]   pe_mat_29_30_io_out_c_data;
  wire                pe_mat_29_30_io_out_c_is_weight;
  wire       [15:0]   pe_mat_29_31_io_out_r_data;
  wire                pe_mat_29_31_io_out_r_stop_weight;
  wire                pe_mat_29_31_io_out_r_stall;
  wire       [15:0]   pe_mat_29_31_io_out_c_data;
  wire                pe_mat_29_31_io_out_c_is_weight;
  wire       [15:0]   pe_mat_30_0_io_out_r_data;
  wire                pe_mat_30_0_io_out_r_stop_weight;
  wire                pe_mat_30_0_io_out_r_stall;
  wire       [15:0]   pe_mat_30_0_io_out_c_data;
  wire                pe_mat_30_0_io_out_c_is_weight;
  wire       [15:0]   pe_mat_30_1_io_out_r_data;
  wire                pe_mat_30_1_io_out_r_stop_weight;
  wire                pe_mat_30_1_io_out_r_stall;
  wire       [15:0]   pe_mat_30_1_io_out_c_data;
  wire                pe_mat_30_1_io_out_c_is_weight;
  wire       [15:0]   pe_mat_30_2_io_out_r_data;
  wire                pe_mat_30_2_io_out_r_stop_weight;
  wire                pe_mat_30_2_io_out_r_stall;
  wire       [15:0]   pe_mat_30_2_io_out_c_data;
  wire                pe_mat_30_2_io_out_c_is_weight;
  wire       [15:0]   pe_mat_30_3_io_out_r_data;
  wire                pe_mat_30_3_io_out_r_stop_weight;
  wire                pe_mat_30_3_io_out_r_stall;
  wire       [15:0]   pe_mat_30_3_io_out_c_data;
  wire                pe_mat_30_3_io_out_c_is_weight;
  wire       [15:0]   pe_mat_30_4_io_out_r_data;
  wire                pe_mat_30_4_io_out_r_stop_weight;
  wire                pe_mat_30_4_io_out_r_stall;
  wire       [15:0]   pe_mat_30_4_io_out_c_data;
  wire                pe_mat_30_4_io_out_c_is_weight;
  wire       [15:0]   pe_mat_30_5_io_out_r_data;
  wire                pe_mat_30_5_io_out_r_stop_weight;
  wire                pe_mat_30_5_io_out_r_stall;
  wire       [15:0]   pe_mat_30_5_io_out_c_data;
  wire                pe_mat_30_5_io_out_c_is_weight;
  wire       [15:0]   pe_mat_30_6_io_out_r_data;
  wire                pe_mat_30_6_io_out_r_stop_weight;
  wire                pe_mat_30_6_io_out_r_stall;
  wire       [15:0]   pe_mat_30_6_io_out_c_data;
  wire                pe_mat_30_6_io_out_c_is_weight;
  wire       [15:0]   pe_mat_30_7_io_out_r_data;
  wire                pe_mat_30_7_io_out_r_stop_weight;
  wire                pe_mat_30_7_io_out_r_stall;
  wire       [15:0]   pe_mat_30_7_io_out_c_data;
  wire                pe_mat_30_7_io_out_c_is_weight;
  wire       [15:0]   pe_mat_30_8_io_out_r_data;
  wire                pe_mat_30_8_io_out_r_stop_weight;
  wire                pe_mat_30_8_io_out_r_stall;
  wire       [15:0]   pe_mat_30_8_io_out_c_data;
  wire                pe_mat_30_8_io_out_c_is_weight;
  wire       [15:0]   pe_mat_30_9_io_out_r_data;
  wire                pe_mat_30_9_io_out_r_stop_weight;
  wire                pe_mat_30_9_io_out_r_stall;
  wire       [15:0]   pe_mat_30_9_io_out_c_data;
  wire                pe_mat_30_9_io_out_c_is_weight;
  wire       [15:0]   pe_mat_30_10_io_out_r_data;
  wire                pe_mat_30_10_io_out_r_stop_weight;
  wire                pe_mat_30_10_io_out_r_stall;
  wire       [15:0]   pe_mat_30_10_io_out_c_data;
  wire                pe_mat_30_10_io_out_c_is_weight;
  wire       [15:0]   pe_mat_30_11_io_out_r_data;
  wire                pe_mat_30_11_io_out_r_stop_weight;
  wire                pe_mat_30_11_io_out_r_stall;
  wire       [15:0]   pe_mat_30_11_io_out_c_data;
  wire                pe_mat_30_11_io_out_c_is_weight;
  wire       [15:0]   pe_mat_30_12_io_out_r_data;
  wire                pe_mat_30_12_io_out_r_stop_weight;
  wire                pe_mat_30_12_io_out_r_stall;
  wire       [15:0]   pe_mat_30_12_io_out_c_data;
  wire                pe_mat_30_12_io_out_c_is_weight;
  wire       [15:0]   pe_mat_30_13_io_out_r_data;
  wire                pe_mat_30_13_io_out_r_stop_weight;
  wire                pe_mat_30_13_io_out_r_stall;
  wire       [15:0]   pe_mat_30_13_io_out_c_data;
  wire                pe_mat_30_13_io_out_c_is_weight;
  wire       [15:0]   pe_mat_30_14_io_out_r_data;
  wire                pe_mat_30_14_io_out_r_stop_weight;
  wire                pe_mat_30_14_io_out_r_stall;
  wire       [15:0]   pe_mat_30_14_io_out_c_data;
  wire                pe_mat_30_14_io_out_c_is_weight;
  wire       [15:0]   pe_mat_30_15_io_out_r_data;
  wire                pe_mat_30_15_io_out_r_stop_weight;
  wire                pe_mat_30_15_io_out_r_stall;
  wire       [15:0]   pe_mat_30_15_io_out_c_data;
  wire                pe_mat_30_15_io_out_c_is_weight;
  wire       [15:0]   pe_mat_30_16_io_out_r_data;
  wire                pe_mat_30_16_io_out_r_stop_weight;
  wire                pe_mat_30_16_io_out_r_stall;
  wire       [15:0]   pe_mat_30_16_io_out_c_data;
  wire                pe_mat_30_16_io_out_c_is_weight;
  wire       [15:0]   pe_mat_30_17_io_out_r_data;
  wire                pe_mat_30_17_io_out_r_stop_weight;
  wire                pe_mat_30_17_io_out_r_stall;
  wire       [15:0]   pe_mat_30_17_io_out_c_data;
  wire                pe_mat_30_17_io_out_c_is_weight;
  wire       [15:0]   pe_mat_30_18_io_out_r_data;
  wire                pe_mat_30_18_io_out_r_stop_weight;
  wire                pe_mat_30_18_io_out_r_stall;
  wire       [15:0]   pe_mat_30_18_io_out_c_data;
  wire                pe_mat_30_18_io_out_c_is_weight;
  wire       [15:0]   pe_mat_30_19_io_out_r_data;
  wire                pe_mat_30_19_io_out_r_stop_weight;
  wire                pe_mat_30_19_io_out_r_stall;
  wire       [15:0]   pe_mat_30_19_io_out_c_data;
  wire                pe_mat_30_19_io_out_c_is_weight;
  wire       [15:0]   pe_mat_30_20_io_out_r_data;
  wire                pe_mat_30_20_io_out_r_stop_weight;
  wire                pe_mat_30_20_io_out_r_stall;
  wire       [15:0]   pe_mat_30_20_io_out_c_data;
  wire                pe_mat_30_20_io_out_c_is_weight;
  wire       [15:0]   pe_mat_30_21_io_out_r_data;
  wire                pe_mat_30_21_io_out_r_stop_weight;
  wire                pe_mat_30_21_io_out_r_stall;
  wire       [15:0]   pe_mat_30_21_io_out_c_data;
  wire                pe_mat_30_21_io_out_c_is_weight;
  wire       [15:0]   pe_mat_30_22_io_out_r_data;
  wire                pe_mat_30_22_io_out_r_stop_weight;
  wire                pe_mat_30_22_io_out_r_stall;
  wire       [15:0]   pe_mat_30_22_io_out_c_data;
  wire                pe_mat_30_22_io_out_c_is_weight;
  wire       [15:0]   pe_mat_30_23_io_out_r_data;
  wire                pe_mat_30_23_io_out_r_stop_weight;
  wire                pe_mat_30_23_io_out_r_stall;
  wire       [15:0]   pe_mat_30_23_io_out_c_data;
  wire                pe_mat_30_23_io_out_c_is_weight;
  wire       [15:0]   pe_mat_30_24_io_out_r_data;
  wire                pe_mat_30_24_io_out_r_stop_weight;
  wire                pe_mat_30_24_io_out_r_stall;
  wire       [15:0]   pe_mat_30_24_io_out_c_data;
  wire                pe_mat_30_24_io_out_c_is_weight;
  wire       [15:0]   pe_mat_30_25_io_out_r_data;
  wire                pe_mat_30_25_io_out_r_stop_weight;
  wire                pe_mat_30_25_io_out_r_stall;
  wire       [15:0]   pe_mat_30_25_io_out_c_data;
  wire                pe_mat_30_25_io_out_c_is_weight;
  wire       [15:0]   pe_mat_30_26_io_out_r_data;
  wire                pe_mat_30_26_io_out_r_stop_weight;
  wire                pe_mat_30_26_io_out_r_stall;
  wire       [15:0]   pe_mat_30_26_io_out_c_data;
  wire                pe_mat_30_26_io_out_c_is_weight;
  wire       [15:0]   pe_mat_30_27_io_out_r_data;
  wire                pe_mat_30_27_io_out_r_stop_weight;
  wire                pe_mat_30_27_io_out_r_stall;
  wire       [15:0]   pe_mat_30_27_io_out_c_data;
  wire                pe_mat_30_27_io_out_c_is_weight;
  wire       [15:0]   pe_mat_30_28_io_out_r_data;
  wire                pe_mat_30_28_io_out_r_stop_weight;
  wire                pe_mat_30_28_io_out_r_stall;
  wire       [15:0]   pe_mat_30_28_io_out_c_data;
  wire                pe_mat_30_28_io_out_c_is_weight;
  wire       [15:0]   pe_mat_30_29_io_out_r_data;
  wire                pe_mat_30_29_io_out_r_stop_weight;
  wire                pe_mat_30_29_io_out_r_stall;
  wire       [15:0]   pe_mat_30_29_io_out_c_data;
  wire                pe_mat_30_29_io_out_c_is_weight;
  wire       [15:0]   pe_mat_30_30_io_out_r_data;
  wire                pe_mat_30_30_io_out_r_stop_weight;
  wire                pe_mat_30_30_io_out_r_stall;
  wire       [15:0]   pe_mat_30_30_io_out_c_data;
  wire                pe_mat_30_30_io_out_c_is_weight;
  wire       [15:0]   pe_mat_30_31_io_out_r_data;
  wire                pe_mat_30_31_io_out_r_stop_weight;
  wire                pe_mat_30_31_io_out_r_stall;
  wire       [15:0]   pe_mat_30_31_io_out_c_data;
  wire                pe_mat_30_31_io_out_c_is_weight;
  wire       [15:0]   pe_mat_31_0_io_out_r_data;
  wire                pe_mat_31_0_io_out_r_stop_weight;
  wire                pe_mat_31_0_io_out_r_stall;
  wire       [15:0]   pe_mat_31_0_io_out_c_data;
  wire                pe_mat_31_0_io_out_c_is_weight;
  wire       [15:0]   pe_mat_31_1_io_out_r_data;
  wire                pe_mat_31_1_io_out_r_stop_weight;
  wire                pe_mat_31_1_io_out_r_stall;
  wire       [15:0]   pe_mat_31_1_io_out_c_data;
  wire                pe_mat_31_1_io_out_c_is_weight;
  wire       [15:0]   pe_mat_31_2_io_out_r_data;
  wire                pe_mat_31_2_io_out_r_stop_weight;
  wire                pe_mat_31_2_io_out_r_stall;
  wire       [15:0]   pe_mat_31_2_io_out_c_data;
  wire                pe_mat_31_2_io_out_c_is_weight;
  wire       [15:0]   pe_mat_31_3_io_out_r_data;
  wire                pe_mat_31_3_io_out_r_stop_weight;
  wire                pe_mat_31_3_io_out_r_stall;
  wire       [15:0]   pe_mat_31_3_io_out_c_data;
  wire                pe_mat_31_3_io_out_c_is_weight;
  wire       [15:0]   pe_mat_31_4_io_out_r_data;
  wire                pe_mat_31_4_io_out_r_stop_weight;
  wire                pe_mat_31_4_io_out_r_stall;
  wire       [15:0]   pe_mat_31_4_io_out_c_data;
  wire                pe_mat_31_4_io_out_c_is_weight;
  wire       [15:0]   pe_mat_31_5_io_out_r_data;
  wire                pe_mat_31_5_io_out_r_stop_weight;
  wire                pe_mat_31_5_io_out_r_stall;
  wire       [15:0]   pe_mat_31_5_io_out_c_data;
  wire                pe_mat_31_5_io_out_c_is_weight;
  wire       [15:0]   pe_mat_31_6_io_out_r_data;
  wire                pe_mat_31_6_io_out_r_stop_weight;
  wire                pe_mat_31_6_io_out_r_stall;
  wire       [15:0]   pe_mat_31_6_io_out_c_data;
  wire                pe_mat_31_6_io_out_c_is_weight;
  wire       [15:0]   pe_mat_31_7_io_out_r_data;
  wire                pe_mat_31_7_io_out_r_stop_weight;
  wire                pe_mat_31_7_io_out_r_stall;
  wire       [15:0]   pe_mat_31_7_io_out_c_data;
  wire                pe_mat_31_7_io_out_c_is_weight;
  wire       [15:0]   pe_mat_31_8_io_out_r_data;
  wire                pe_mat_31_8_io_out_r_stop_weight;
  wire                pe_mat_31_8_io_out_r_stall;
  wire       [15:0]   pe_mat_31_8_io_out_c_data;
  wire                pe_mat_31_8_io_out_c_is_weight;
  wire       [15:0]   pe_mat_31_9_io_out_r_data;
  wire                pe_mat_31_9_io_out_r_stop_weight;
  wire                pe_mat_31_9_io_out_r_stall;
  wire       [15:0]   pe_mat_31_9_io_out_c_data;
  wire                pe_mat_31_9_io_out_c_is_weight;
  wire       [15:0]   pe_mat_31_10_io_out_r_data;
  wire                pe_mat_31_10_io_out_r_stop_weight;
  wire                pe_mat_31_10_io_out_r_stall;
  wire       [15:0]   pe_mat_31_10_io_out_c_data;
  wire                pe_mat_31_10_io_out_c_is_weight;
  wire       [15:0]   pe_mat_31_11_io_out_r_data;
  wire                pe_mat_31_11_io_out_r_stop_weight;
  wire                pe_mat_31_11_io_out_r_stall;
  wire       [15:0]   pe_mat_31_11_io_out_c_data;
  wire                pe_mat_31_11_io_out_c_is_weight;
  wire       [15:0]   pe_mat_31_12_io_out_r_data;
  wire                pe_mat_31_12_io_out_r_stop_weight;
  wire                pe_mat_31_12_io_out_r_stall;
  wire       [15:0]   pe_mat_31_12_io_out_c_data;
  wire                pe_mat_31_12_io_out_c_is_weight;
  wire       [15:0]   pe_mat_31_13_io_out_r_data;
  wire                pe_mat_31_13_io_out_r_stop_weight;
  wire                pe_mat_31_13_io_out_r_stall;
  wire       [15:0]   pe_mat_31_13_io_out_c_data;
  wire                pe_mat_31_13_io_out_c_is_weight;
  wire       [15:0]   pe_mat_31_14_io_out_r_data;
  wire                pe_mat_31_14_io_out_r_stop_weight;
  wire                pe_mat_31_14_io_out_r_stall;
  wire       [15:0]   pe_mat_31_14_io_out_c_data;
  wire                pe_mat_31_14_io_out_c_is_weight;
  wire       [15:0]   pe_mat_31_15_io_out_r_data;
  wire                pe_mat_31_15_io_out_r_stop_weight;
  wire                pe_mat_31_15_io_out_r_stall;
  wire       [15:0]   pe_mat_31_15_io_out_c_data;
  wire                pe_mat_31_15_io_out_c_is_weight;
  wire       [15:0]   pe_mat_31_16_io_out_r_data;
  wire                pe_mat_31_16_io_out_r_stop_weight;
  wire                pe_mat_31_16_io_out_r_stall;
  wire       [15:0]   pe_mat_31_16_io_out_c_data;
  wire                pe_mat_31_16_io_out_c_is_weight;
  wire       [15:0]   pe_mat_31_17_io_out_r_data;
  wire                pe_mat_31_17_io_out_r_stop_weight;
  wire                pe_mat_31_17_io_out_r_stall;
  wire       [15:0]   pe_mat_31_17_io_out_c_data;
  wire                pe_mat_31_17_io_out_c_is_weight;
  wire       [15:0]   pe_mat_31_18_io_out_r_data;
  wire                pe_mat_31_18_io_out_r_stop_weight;
  wire                pe_mat_31_18_io_out_r_stall;
  wire       [15:0]   pe_mat_31_18_io_out_c_data;
  wire                pe_mat_31_18_io_out_c_is_weight;
  wire       [15:0]   pe_mat_31_19_io_out_r_data;
  wire                pe_mat_31_19_io_out_r_stop_weight;
  wire                pe_mat_31_19_io_out_r_stall;
  wire       [15:0]   pe_mat_31_19_io_out_c_data;
  wire                pe_mat_31_19_io_out_c_is_weight;
  wire       [15:0]   pe_mat_31_20_io_out_r_data;
  wire                pe_mat_31_20_io_out_r_stop_weight;
  wire                pe_mat_31_20_io_out_r_stall;
  wire       [15:0]   pe_mat_31_20_io_out_c_data;
  wire                pe_mat_31_20_io_out_c_is_weight;
  wire       [15:0]   pe_mat_31_21_io_out_r_data;
  wire                pe_mat_31_21_io_out_r_stop_weight;
  wire                pe_mat_31_21_io_out_r_stall;
  wire       [15:0]   pe_mat_31_21_io_out_c_data;
  wire                pe_mat_31_21_io_out_c_is_weight;
  wire       [15:0]   pe_mat_31_22_io_out_r_data;
  wire                pe_mat_31_22_io_out_r_stop_weight;
  wire                pe_mat_31_22_io_out_r_stall;
  wire       [15:0]   pe_mat_31_22_io_out_c_data;
  wire                pe_mat_31_22_io_out_c_is_weight;
  wire       [15:0]   pe_mat_31_23_io_out_r_data;
  wire                pe_mat_31_23_io_out_r_stop_weight;
  wire                pe_mat_31_23_io_out_r_stall;
  wire       [15:0]   pe_mat_31_23_io_out_c_data;
  wire                pe_mat_31_23_io_out_c_is_weight;
  wire       [15:0]   pe_mat_31_24_io_out_r_data;
  wire                pe_mat_31_24_io_out_r_stop_weight;
  wire                pe_mat_31_24_io_out_r_stall;
  wire       [15:0]   pe_mat_31_24_io_out_c_data;
  wire                pe_mat_31_24_io_out_c_is_weight;
  wire       [15:0]   pe_mat_31_25_io_out_r_data;
  wire                pe_mat_31_25_io_out_r_stop_weight;
  wire                pe_mat_31_25_io_out_r_stall;
  wire       [15:0]   pe_mat_31_25_io_out_c_data;
  wire                pe_mat_31_25_io_out_c_is_weight;
  wire       [15:0]   pe_mat_31_26_io_out_r_data;
  wire                pe_mat_31_26_io_out_r_stop_weight;
  wire                pe_mat_31_26_io_out_r_stall;
  wire       [15:0]   pe_mat_31_26_io_out_c_data;
  wire                pe_mat_31_26_io_out_c_is_weight;
  wire       [15:0]   pe_mat_31_27_io_out_r_data;
  wire                pe_mat_31_27_io_out_r_stop_weight;
  wire                pe_mat_31_27_io_out_r_stall;
  wire       [15:0]   pe_mat_31_27_io_out_c_data;
  wire                pe_mat_31_27_io_out_c_is_weight;
  wire       [15:0]   pe_mat_31_28_io_out_r_data;
  wire                pe_mat_31_28_io_out_r_stop_weight;
  wire                pe_mat_31_28_io_out_r_stall;
  wire       [15:0]   pe_mat_31_28_io_out_c_data;
  wire                pe_mat_31_28_io_out_c_is_weight;
  wire       [15:0]   pe_mat_31_29_io_out_r_data;
  wire                pe_mat_31_29_io_out_r_stop_weight;
  wire                pe_mat_31_29_io_out_r_stall;
  wire       [15:0]   pe_mat_31_29_io_out_c_data;
  wire                pe_mat_31_29_io_out_c_is_weight;
  wire       [15:0]   pe_mat_31_30_io_out_r_data;
  wire                pe_mat_31_30_io_out_r_stop_weight;
  wire                pe_mat_31_30_io_out_r_stall;
  wire       [15:0]   pe_mat_31_30_io_out_c_data;
  wire                pe_mat_31_30_io_out_c_is_weight;
  wire       [15:0]   pe_mat_31_31_io_out_r_data;
  wire                pe_mat_31_31_io_out_r_stop_weight;
  wire                pe_mat_31_31_io_out_r_stall;
  wire       [15:0]   pe_mat_31_31_io_out_c_data;
  wire                pe_mat_31_31_io_out_c_is_weight;

  PEWS_1023 pe_mat_0_0 (
    .io_in_r_data         (io_in_r_0_data[15:0]           ), //i
    .io_in_r_stop_weight  (io_in_r_0_stop_weight          ), //i
    .io_in_r_stall        (io_in_r_0_stall                ), //i
    .io_out_r_data        (pe_mat_0_0_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_0_0_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_0_0_io_out_r_stall      ), //o
    .io_in_c_data         (io_in_c_0_data[15:0]           ), //i
    .io_in_c_is_weight    (io_in_c_0_is_weight            ), //i
    .io_out_c_data        (pe_mat_0_0_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_0_0_io_out_c_is_weight  ), //o
    .clk                  (clk                            ), //i
    .reset                (reset                          )  //i
  );
  PEWS_1023 pe_mat_0_1 (
    .io_in_r_data         (pe_mat_0_0_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_0_0_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_0_0_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_0_1_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_0_1_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_0_1_io_out_r_stall      ), //o
    .io_in_c_data         (io_in_c_1_data[15:0]           ), //i
    .io_in_c_is_weight    (io_in_c_1_is_weight            ), //i
    .io_out_c_data        (pe_mat_0_1_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_0_1_io_out_c_is_weight  ), //o
    .clk                  (clk                            ), //i
    .reset                (reset                          )  //i
  );
  PEWS_1023 pe_mat_0_2 (
    .io_in_r_data         (pe_mat_0_1_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_0_1_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_0_1_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_0_2_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_0_2_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_0_2_io_out_r_stall      ), //o
    .io_in_c_data         (io_in_c_2_data[15:0]           ), //i
    .io_in_c_is_weight    (io_in_c_2_is_weight            ), //i
    .io_out_c_data        (pe_mat_0_2_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_0_2_io_out_c_is_weight  ), //o
    .clk                  (clk                            ), //i
    .reset                (reset                          )  //i
  );
  PEWS_1023 pe_mat_0_3 (
    .io_in_r_data         (pe_mat_0_2_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_0_2_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_0_2_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_0_3_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_0_3_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_0_3_io_out_r_stall      ), //o
    .io_in_c_data         (io_in_c_3_data[15:0]           ), //i
    .io_in_c_is_weight    (io_in_c_3_is_weight            ), //i
    .io_out_c_data        (pe_mat_0_3_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_0_3_io_out_c_is_weight  ), //o
    .clk                  (clk                            ), //i
    .reset                (reset                          )  //i
  );
  PEWS_1023 pe_mat_0_4 (
    .io_in_r_data         (pe_mat_0_3_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_0_3_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_0_3_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_0_4_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_0_4_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_0_4_io_out_r_stall      ), //o
    .io_in_c_data         (io_in_c_4_data[15:0]           ), //i
    .io_in_c_is_weight    (io_in_c_4_is_weight            ), //i
    .io_out_c_data        (pe_mat_0_4_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_0_4_io_out_c_is_weight  ), //o
    .clk                  (clk                            ), //i
    .reset                (reset                          )  //i
  );
  PEWS_1023 pe_mat_0_5 (
    .io_in_r_data         (pe_mat_0_4_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_0_4_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_0_4_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_0_5_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_0_5_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_0_5_io_out_r_stall      ), //o
    .io_in_c_data         (io_in_c_5_data[15:0]           ), //i
    .io_in_c_is_weight    (io_in_c_5_is_weight            ), //i
    .io_out_c_data        (pe_mat_0_5_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_0_5_io_out_c_is_weight  ), //o
    .clk                  (clk                            ), //i
    .reset                (reset                          )  //i
  );
  PEWS_1023 pe_mat_0_6 (
    .io_in_r_data         (pe_mat_0_5_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_0_5_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_0_5_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_0_6_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_0_6_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_0_6_io_out_r_stall      ), //o
    .io_in_c_data         (io_in_c_6_data[15:0]           ), //i
    .io_in_c_is_weight    (io_in_c_6_is_weight            ), //i
    .io_out_c_data        (pe_mat_0_6_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_0_6_io_out_c_is_weight  ), //o
    .clk                  (clk                            ), //i
    .reset                (reset                          )  //i
  );
  PEWS_1023 pe_mat_0_7 (
    .io_in_r_data         (pe_mat_0_6_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_0_6_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_0_6_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_0_7_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_0_7_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_0_7_io_out_r_stall      ), //o
    .io_in_c_data         (io_in_c_7_data[15:0]           ), //i
    .io_in_c_is_weight    (io_in_c_7_is_weight            ), //i
    .io_out_c_data        (pe_mat_0_7_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_0_7_io_out_c_is_weight  ), //o
    .clk                  (clk                            ), //i
    .reset                (reset                          )  //i
  );
  PEWS_1023 pe_mat_0_8 (
    .io_in_r_data         (pe_mat_0_7_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_0_7_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_0_7_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_0_8_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_0_8_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_0_8_io_out_r_stall      ), //o
    .io_in_c_data         (io_in_c_8_data[15:0]           ), //i
    .io_in_c_is_weight    (io_in_c_8_is_weight            ), //i
    .io_out_c_data        (pe_mat_0_8_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_0_8_io_out_c_is_weight  ), //o
    .clk                  (clk                            ), //i
    .reset                (reset                          )  //i
  );
  PEWS_1023 pe_mat_0_9 (
    .io_in_r_data         (pe_mat_0_8_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_0_8_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_0_8_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_0_9_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_0_9_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_0_9_io_out_r_stall      ), //o
    .io_in_c_data         (io_in_c_9_data[15:0]           ), //i
    .io_in_c_is_weight    (io_in_c_9_is_weight            ), //i
    .io_out_c_data        (pe_mat_0_9_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_0_9_io_out_c_is_weight  ), //o
    .clk                  (clk                            ), //i
    .reset                (reset                          )  //i
  );
  PEWS_1023 pe_mat_0_10 (
    .io_in_r_data         (pe_mat_0_9_io_out_r_data[15:0]  ), //i
    .io_in_r_stop_weight  (pe_mat_0_9_io_out_r_stop_weight ), //i
    .io_in_r_stall        (pe_mat_0_9_io_out_r_stall       ), //i
    .io_out_r_data        (pe_mat_0_10_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_0_10_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_0_10_io_out_r_stall      ), //o
    .io_in_c_data         (io_in_c_10_data[15:0]           ), //i
    .io_in_c_is_weight    (io_in_c_10_is_weight            ), //i
    .io_out_c_data        (pe_mat_0_10_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_0_10_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_0_11 (
    .io_in_r_data         (pe_mat_0_10_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_0_10_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_0_10_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_0_11_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_0_11_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_0_11_io_out_r_stall      ), //o
    .io_in_c_data         (io_in_c_11_data[15:0]           ), //i
    .io_in_c_is_weight    (io_in_c_11_is_weight            ), //i
    .io_out_c_data        (pe_mat_0_11_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_0_11_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_0_12 (
    .io_in_r_data         (pe_mat_0_11_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_0_11_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_0_11_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_0_12_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_0_12_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_0_12_io_out_r_stall      ), //o
    .io_in_c_data         (io_in_c_12_data[15:0]           ), //i
    .io_in_c_is_weight    (io_in_c_12_is_weight            ), //i
    .io_out_c_data        (pe_mat_0_12_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_0_12_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_0_13 (
    .io_in_r_data         (pe_mat_0_12_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_0_12_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_0_12_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_0_13_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_0_13_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_0_13_io_out_r_stall      ), //o
    .io_in_c_data         (io_in_c_13_data[15:0]           ), //i
    .io_in_c_is_weight    (io_in_c_13_is_weight            ), //i
    .io_out_c_data        (pe_mat_0_13_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_0_13_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_0_14 (
    .io_in_r_data         (pe_mat_0_13_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_0_13_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_0_13_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_0_14_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_0_14_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_0_14_io_out_r_stall      ), //o
    .io_in_c_data         (io_in_c_14_data[15:0]           ), //i
    .io_in_c_is_weight    (io_in_c_14_is_weight            ), //i
    .io_out_c_data        (pe_mat_0_14_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_0_14_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_0_15 (
    .io_in_r_data         (pe_mat_0_14_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_0_14_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_0_14_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_0_15_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_0_15_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_0_15_io_out_r_stall      ), //o
    .io_in_c_data         (io_in_c_15_data[15:0]           ), //i
    .io_in_c_is_weight    (io_in_c_15_is_weight            ), //i
    .io_out_c_data        (pe_mat_0_15_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_0_15_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_0_16 (
    .io_in_r_data         (pe_mat_0_15_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_0_15_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_0_15_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_0_16_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_0_16_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_0_16_io_out_r_stall      ), //o
    .io_in_c_data         (io_in_c_16_data[15:0]           ), //i
    .io_in_c_is_weight    (io_in_c_16_is_weight            ), //i
    .io_out_c_data        (pe_mat_0_16_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_0_16_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_0_17 (
    .io_in_r_data         (pe_mat_0_16_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_0_16_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_0_16_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_0_17_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_0_17_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_0_17_io_out_r_stall      ), //o
    .io_in_c_data         (io_in_c_17_data[15:0]           ), //i
    .io_in_c_is_weight    (io_in_c_17_is_weight            ), //i
    .io_out_c_data        (pe_mat_0_17_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_0_17_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_0_18 (
    .io_in_r_data         (pe_mat_0_17_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_0_17_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_0_17_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_0_18_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_0_18_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_0_18_io_out_r_stall      ), //o
    .io_in_c_data         (io_in_c_18_data[15:0]           ), //i
    .io_in_c_is_weight    (io_in_c_18_is_weight            ), //i
    .io_out_c_data        (pe_mat_0_18_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_0_18_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_0_19 (
    .io_in_r_data         (pe_mat_0_18_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_0_18_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_0_18_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_0_19_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_0_19_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_0_19_io_out_r_stall      ), //o
    .io_in_c_data         (io_in_c_19_data[15:0]           ), //i
    .io_in_c_is_weight    (io_in_c_19_is_weight            ), //i
    .io_out_c_data        (pe_mat_0_19_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_0_19_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_0_20 (
    .io_in_r_data         (pe_mat_0_19_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_0_19_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_0_19_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_0_20_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_0_20_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_0_20_io_out_r_stall      ), //o
    .io_in_c_data         (io_in_c_20_data[15:0]           ), //i
    .io_in_c_is_weight    (io_in_c_20_is_weight            ), //i
    .io_out_c_data        (pe_mat_0_20_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_0_20_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_0_21 (
    .io_in_r_data         (pe_mat_0_20_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_0_20_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_0_20_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_0_21_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_0_21_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_0_21_io_out_r_stall      ), //o
    .io_in_c_data         (io_in_c_21_data[15:0]           ), //i
    .io_in_c_is_weight    (io_in_c_21_is_weight            ), //i
    .io_out_c_data        (pe_mat_0_21_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_0_21_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_0_22 (
    .io_in_r_data         (pe_mat_0_21_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_0_21_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_0_21_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_0_22_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_0_22_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_0_22_io_out_r_stall      ), //o
    .io_in_c_data         (io_in_c_22_data[15:0]           ), //i
    .io_in_c_is_weight    (io_in_c_22_is_weight            ), //i
    .io_out_c_data        (pe_mat_0_22_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_0_22_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_0_23 (
    .io_in_r_data         (pe_mat_0_22_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_0_22_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_0_22_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_0_23_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_0_23_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_0_23_io_out_r_stall      ), //o
    .io_in_c_data         (io_in_c_23_data[15:0]           ), //i
    .io_in_c_is_weight    (io_in_c_23_is_weight            ), //i
    .io_out_c_data        (pe_mat_0_23_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_0_23_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_0_24 (
    .io_in_r_data         (pe_mat_0_23_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_0_23_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_0_23_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_0_24_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_0_24_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_0_24_io_out_r_stall      ), //o
    .io_in_c_data         (io_in_c_24_data[15:0]           ), //i
    .io_in_c_is_weight    (io_in_c_24_is_weight            ), //i
    .io_out_c_data        (pe_mat_0_24_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_0_24_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_0_25 (
    .io_in_r_data         (pe_mat_0_24_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_0_24_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_0_24_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_0_25_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_0_25_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_0_25_io_out_r_stall      ), //o
    .io_in_c_data         (io_in_c_25_data[15:0]           ), //i
    .io_in_c_is_weight    (io_in_c_25_is_weight            ), //i
    .io_out_c_data        (pe_mat_0_25_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_0_25_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_0_26 (
    .io_in_r_data         (pe_mat_0_25_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_0_25_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_0_25_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_0_26_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_0_26_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_0_26_io_out_r_stall      ), //o
    .io_in_c_data         (io_in_c_26_data[15:0]           ), //i
    .io_in_c_is_weight    (io_in_c_26_is_weight            ), //i
    .io_out_c_data        (pe_mat_0_26_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_0_26_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_0_27 (
    .io_in_r_data         (pe_mat_0_26_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_0_26_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_0_26_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_0_27_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_0_27_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_0_27_io_out_r_stall      ), //o
    .io_in_c_data         (io_in_c_27_data[15:0]           ), //i
    .io_in_c_is_weight    (io_in_c_27_is_weight            ), //i
    .io_out_c_data        (pe_mat_0_27_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_0_27_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_0_28 (
    .io_in_r_data         (pe_mat_0_27_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_0_27_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_0_27_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_0_28_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_0_28_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_0_28_io_out_r_stall      ), //o
    .io_in_c_data         (io_in_c_28_data[15:0]           ), //i
    .io_in_c_is_weight    (io_in_c_28_is_weight            ), //i
    .io_out_c_data        (pe_mat_0_28_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_0_28_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_0_29 (
    .io_in_r_data         (pe_mat_0_28_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_0_28_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_0_28_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_0_29_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_0_29_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_0_29_io_out_r_stall      ), //o
    .io_in_c_data         (io_in_c_29_data[15:0]           ), //i
    .io_in_c_is_weight    (io_in_c_29_is_weight            ), //i
    .io_out_c_data        (pe_mat_0_29_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_0_29_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_0_30 (
    .io_in_r_data         (pe_mat_0_29_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_0_29_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_0_29_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_0_30_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_0_30_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_0_30_io_out_r_stall      ), //o
    .io_in_c_data         (io_in_c_30_data[15:0]           ), //i
    .io_in_c_is_weight    (io_in_c_30_is_weight            ), //i
    .io_out_c_data        (pe_mat_0_30_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_0_30_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_0_31 (
    .io_in_r_data         (pe_mat_0_30_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_0_30_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_0_30_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_0_31_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_0_31_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_0_31_io_out_r_stall      ), //o
    .io_in_c_data         (io_in_c_31_data[15:0]           ), //i
    .io_in_c_is_weight    (io_in_c_31_is_weight            ), //i
    .io_out_c_data        (pe_mat_0_31_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_0_31_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_1_0 (
    .io_in_r_data         (io_in_r_1_data[15:0]           ), //i
    .io_in_r_stop_weight  (io_in_r_1_stop_weight          ), //i
    .io_in_r_stall        (io_in_r_1_stall                ), //i
    .io_out_r_data        (pe_mat_1_0_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_1_0_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_1_0_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_0_0_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_0_0_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_1_0_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_1_0_io_out_c_is_weight  ), //o
    .clk                  (clk                            ), //i
    .reset                (reset                          )  //i
  );
  PEWS_1023 pe_mat_1_1 (
    .io_in_r_data         (pe_mat_1_0_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_1_0_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_1_0_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_1_1_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_1_1_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_1_1_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_0_1_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_0_1_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_1_1_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_1_1_io_out_c_is_weight  ), //o
    .clk                  (clk                            ), //i
    .reset                (reset                          )  //i
  );
  PEWS_1023 pe_mat_1_2 (
    .io_in_r_data         (pe_mat_1_1_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_1_1_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_1_1_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_1_2_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_1_2_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_1_2_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_0_2_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_0_2_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_1_2_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_1_2_io_out_c_is_weight  ), //o
    .clk                  (clk                            ), //i
    .reset                (reset                          )  //i
  );
  PEWS_1023 pe_mat_1_3 (
    .io_in_r_data         (pe_mat_1_2_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_1_2_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_1_2_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_1_3_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_1_3_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_1_3_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_0_3_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_0_3_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_1_3_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_1_3_io_out_c_is_weight  ), //o
    .clk                  (clk                            ), //i
    .reset                (reset                          )  //i
  );
  PEWS_1023 pe_mat_1_4 (
    .io_in_r_data         (pe_mat_1_3_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_1_3_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_1_3_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_1_4_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_1_4_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_1_4_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_0_4_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_0_4_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_1_4_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_1_4_io_out_c_is_weight  ), //o
    .clk                  (clk                            ), //i
    .reset                (reset                          )  //i
  );
  PEWS_1023 pe_mat_1_5 (
    .io_in_r_data         (pe_mat_1_4_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_1_4_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_1_4_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_1_5_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_1_5_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_1_5_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_0_5_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_0_5_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_1_5_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_1_5_io_out_c_is_weight  ), //o
    .clk                  (clk                            ), //i
    .reset                (reset                          )  //i
  );
  PEWS_1023 pe_mat_1_6 (
    .io_in_r_data         (pe_mat_1_5_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_1_5_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_1_5_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_1_6_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_1_6_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_1_6_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_0_6_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_0_6_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_1_6_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_1_6_io_out_c_is_weight  ), //o
    .clk                  (clk                            ), //i
    .reset                (reset                          )  //i
  );
  PEWS_1023 pe_mat_1_7 (
    .io_in_r_data         (pe_mat_1_6_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_1_6_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_1_6_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_1_7_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_1_7_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_1_7_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_0_7_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_0_7_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_1_7_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_1_7_io_out_c_is_weight  ), //o
    .clk                  (clk                            ), //i
    .reset                (reset                          )  //i
  );
  PEWS_1023 pe_mat_1_8 (
    .io_in_r_data         (pe_mat_1_7_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_1_7_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_1_7_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_1_8_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_1_8_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_1_8_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_0_8_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_0_8_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_1_8_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_1_8_io_out_c_is_weight  ), //o
    .clk                  (clk                            ), //i
    .reset                (reset                          )  //i
  );
  PEWS_1023 pe_mat_1_9 (
    .io_in_r_data         (pe_mat_1_8_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_1_8_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_1_8_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_1_9_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_1_9_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_1_9_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_0_9_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_0_9_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_1_9_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_1_9_io_out_c_is_weight  ), //o
    .clk                  (clk                            ), //i
    .reset                (reset                          )  //i
  );
  PEWS_1023 pe_mat_1_10 (
    .io_in_r_data         (pe_mat_1_9_io_out_r_data[15:0]  ), //i
    .io_in_r_stop_weight  (pe_mat_1_9_io_out_r_stop_weight ), //i
    .io_in_r_stall        (pe_mat_1_9_io_out_r_stall       ), //i
    .io_out_r_data        (pe_mat_1_10_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_1_10_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_1_10_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_0_10_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_0_10_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_1_10_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_1_10_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_1_11 (
    .io_in_r_data         (pe_mat_1_10_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_1_10_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_1_10_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_1_11_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_1_11_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_1_11_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_0_11_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_0_11_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_1_11_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_1_11_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_1_12 (
    .io_in_r_data         (pe_mat_1_11_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_1_11_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_1_11_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_1_12_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_1_12_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_1_12_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_0_12_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_0_12_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_1_12_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_1_12_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_1_13 (
    .io_in_r_data         (pe_mat_1_12_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_1_12_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_1_12_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_1_13_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_1_13_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_1_13_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_0_13_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_0_13_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_1_13_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_1_13_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_1_14 (
    .io_in_r_data         (pe_mat_1_13_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_1_13_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_1_13_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_1_14_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_1_14_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_1_14_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_0_14_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_0_14_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_1_14_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_1_14_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_1_15 (
    .io_in_r_data         (pe_mat_1_14_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_1_14_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_1_14_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_1_15_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_1_15_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_1_15_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_0_15_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_0_15_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_1_15_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_1_15_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_1_16 (
    .io_in_r_data         (pe_mat_1_15_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_1_15_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_1_15_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_1_16_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_1_16_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_1_16_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_0_16_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_0_16_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_1_16_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_1_16_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_1_17 (
    .io_in_r_data         (pe_mat_1_16_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_1_16_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_1_16_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_1_17_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_1_17_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_1_17_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_0_17_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_0_17_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_1_17_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_1_17_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_1_18 (
    .io_in_r_data         (pe_mat_1_17_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_1_17_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_1_17_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_1_18_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_1_18_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_1_18_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_0_18_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_0_18_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_1_18_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_1_18_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_1_19 (
    .io_in_r_data         (pe_mat_1_18_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_1_18_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_1_18_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_1_19_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_1_19_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_1_19_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_0_19_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_0_19_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_1_19_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_1_19_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_1_20 (
    .io_in_r_data         (pe_mat_1_19_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_1_19_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_1_19_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_1_20_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_1_20_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_1_20_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_0_20_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_0_20_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_1_20_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_1_20_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_1_21 (
    .io_in_r_data         (pe_mat_1_20_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_1_20_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_1_20_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_1_21_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_1_21_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_1_21_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_0_21_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_0_21_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_1_21_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_1_21_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_1_22 (
    .io_in_r_data         (pe_mat_1_21_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_1_21_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_1_21_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_1_22_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_1_22_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_1_22_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_0_22_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_0_22_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_1_22_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_1_22_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_1_23 (
    .io_in_r_data         (pe_mat_1_22_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_1_22_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_1_22_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_1_23_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_1_23_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_1_23_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_0_23_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_0_23_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_1_23_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_1_23_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_1_24 (
    .io_in_r_data         (pe_mat_1_23_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_1_23_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_1_23_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_1_24_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_1_24_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_1_24_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_0_24_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_0_24_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_1_24_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_1_24_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_1_25 (
    .io_in_r_data         (pe_mat_1_24_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_1_24_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_1_24_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_1_25_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_1_25_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_1_25_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_0_25_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_0_25_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_1_25_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_1_25_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_1_26 (
    .io_in_r_data         (pe_mat_1_25_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_1_25_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_1_25_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_1_26_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_1_26_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_1_26_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_0_26_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_0_26_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_1_26_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_1_26_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_1_27 (
    .io_in_r_data         (pe_mat_1_26_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_1_26_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_1_26_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_1_27_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_1_27_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_1_27_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_0_27_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_0_27_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_1_27_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_1_27_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_1_28 (
    .io_in_r_data         (pe_mat_1_27_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_1_27_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_1_27_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_1_28_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_1_28_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_1_28_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_0_28_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_0_28_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_1_28_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_1_28_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_1_29 (
    .io_in_r_data         (pe_mat_1_28_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_1_28_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_1_28_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_1_29_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_1_29_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_1_29_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_0_29_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_0_29_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_1_29_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_1_29_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_1_30 (
    .io_in_r_data         (pe_mat_1_29_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_1_29_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_1_29_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_1_30_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_1_30_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_1_30_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_0_30_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_0_30_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_1_30_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_1_30_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_1_31 (
    .io_in_r_data         (pe_mat_1_30_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_1_30_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_1_30_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_1_31_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_1_31_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_1_31_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_0_31_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_0_31_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_1_31_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_1_31_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_2_0 (
    .io_in_r_data         (io_in_r_2_data[15:0]           ), //i
    .io_in_r_stop_weight  (io_in_r_2_stop_weight          ), //i
    .io_in_r_stall        (io_in_r_2_stall                ), //i
    .io_out_r_data        (pe_mat_2_0_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_2_0_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_2_0_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_1_0_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_1_0_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_2_0_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_2_0_io_out_c_is_weight  ), //o
    .clk                  (clk                            ), //i
    .reset                (reset                          )  //i
  );
  PEWS_1023 pe_mat_2_1 (
    .io_in_r_data         (pe_mat_2_0_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_2_0_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_2_0_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_2_1_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_2_1_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_2_1_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_1_1_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_1_1_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_2_1_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_2_1_io_out_c_is_weight  ), //o
    .clk                  (clk                            ), //i
    .reset                (reset                          )  //i
  );
  PEWS_1023 pe_mat_2_2 (
    .io_in_r_data         (pe_mat_2_1_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_2_1_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_2_1_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_2_2_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_2_2_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_2_2_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_1_2_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_1_2_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_2_2_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_2_2_io_out_c_is_weight  ), //o
    .clk                  (clk                            ), //i
    .reset                (reset                          )  //i
  );
  PEWS_1023 pe_mat_2_3 (
    .io_in_r_data         (pe_mat_2_2_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_2_2_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_2_2_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_2_3_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_2_3_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_2_3_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_1_3_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_1_3_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_2_3_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_2_3_io_out_c_is_weight  ), //o
    .clk                  (clk                            ), //i
    .reset                (reset                          )  //i
  );
  PEWS_1023 pe_mat_2_4 (
    .io_in_r_data         (pe_mat_2_3_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_2_3_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_2_3_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_2_4_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_2_4_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_2_4_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_1_4_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_1_4_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_2_4_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_2_4_io_out_c_is_weight  ), //o
    .clk                  (clk                            ), //i
    .reset                (reset                          )  //i
  );
  PEWS_1023 pe_mat_2_5 (
    .io_in_r_data         (pe_mat_2_4_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_2_4_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_2_4_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_2_5_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_2_5_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_2_5_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_1_5_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_1_5_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_2_5_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_2_5_io_out_c_is_weight  ), //o
    .clk                  (clk                            ), //i
    .reset                (reset                          )  //i
  );
  PEWS_1023 pe_mat_2_6 (
    .io_in_r_data         (pe_mat_2_5_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_2_5_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_2_5_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_2_6_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_2_6_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_2_6_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_1_6_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_1_6_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_2_6_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_2_6_io_out_c_is_weight  ), //o
    .clk                  (clk                            ), //i
    .reset                (reset                          )  //i
  );
  PEWS_1023 pe_mat_2_7 (
    .io_in_r_data         (pe_mat_2_6_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_2_6_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_2_6_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_2_7_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_2_7_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_2_7_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_1_7_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_1_7_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_2_7_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_2_7_io_out_c_is_weight  ), //o
    .clk                  (clk                            ), //i
    .reset                (reset                          )  //i
  );
  PEWS_1023 pe_mat_2_8 (
    .io_in_r_data         (pe_mat_2_7_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_2_7_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_2_7_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_2_8_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_2_8_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_2_8_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_1_8_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_1_8_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_2_8_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_2_8_io_out_c_is_weight  ), //o
    .clk                  (clk                            ), //i
    .reset                (reset                          )  //i
  );
  PEWS_1023 pe_mat_2_9 (
    .io_in_r_data         (pe_mat_2_8_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_2_8_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_2_8_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_2_9_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_2_9_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_2_9_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_1_9_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_1_9_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_2_9_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_2_9_io_out_c_is_weight  ), //o
    .clk                  (clk                            ), //i
    .reset                (reset                          )  //i
  );
  PEWS_1023 pe_mat_2_10 (
    .io_in_r_data         (pe_mat_2_9_io_out_r_data[15:0]  ), //i
    .io_in_r_stop_weight  (pe_mat_2_9_io_out_r_stop_weight ), //i
    .io_in_r_stall        (pe_mat_2_9_io_out_r_stall       ), //i
    .io_out_r_data        (pe_mat_2_10_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_2_10_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_2_10_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_1_10_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_1_10_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_2_10_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_2_10_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_2_11 (
    .io_in_r_data         (pe_mat_2_10_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_2_10_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_2_10_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_2_11_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_2_11_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_2_11_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_1_11_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_1_11_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_2_11_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_2_11_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_2_12 (
    .io_in_r_data         (pe_mat_2_11_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_2_11_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_2_11_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_2_12_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_2_12_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_2_12_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_1_12_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_1_12_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_2_12_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_2_12_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_2_13 (
    .io_in_r_data         (pe_mat_2_12_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_2_12_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_2_12_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_2_13_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_2_13_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_2_13_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_1_13_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_1_13_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_2_13_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_2_13_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_2_14 (
    .io_in_r_data         (pe_mat_2_13_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_2_13_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_2_13_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_2_14_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_2_14_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_2_14_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_1_14_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_1_14_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_2_14_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_2_14_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_2_15 (
    .io_in_r_data         (pe_mat_2_14_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_2_14_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_2_14_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_2_15_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_2_15_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_2_15_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_1_15_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_1_15_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_2_15_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_2_15_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_2_16 (
    .io_in_r_data         (pe_mat_2_15_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_2_15_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_2_15_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_2_16_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_2_16_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_2_16_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_1_16_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_1_16_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_2_16_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_2_16_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_2_17 (
    .io_in_r_data         (pe_mat_2_16_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_2_16_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_2_16_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_2_17_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_2_17_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_2_17_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_1_17_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_1_17_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_2_17_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_2_17_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_2_18 (
    .io_in_r_data         (pe_mat_2_17_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_2_17_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_2_17_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_2_18_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_2_18_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_2_18_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_1_18_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_1_18_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_2_18_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_2_18_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_2_19 (
    .io_in_r_data         (pe_mat_2_18_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_2_18_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_2_18_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_2_19_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_2_19_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_2_19_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_1_19_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_1_19_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_2_19_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_2_19_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_2_20 (
    .io_in_r_data         (pe_mat_2_19_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_2_19_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_2_19_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_2_20_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_2_20_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_2_20_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_1_20_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_1_20_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_2_20_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_2_20_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_2_21 (
    .io_in_r_data         (pe_mat_2_20_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_2_20_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_2_20_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_2_21_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_2_21_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_2_21_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_1_21_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_1_21_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_2_21_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_2_21_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_2_22 (
    .io_in_r_data         (pe_mat_2_21_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_2_21_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_2_21_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_2_22_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_2_22_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_2_22_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_1_22_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_1_22_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_2_22_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_2_22_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_2_23 (
    .io_in_r_data         (pe_mat_2_22_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_2_22_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_2_22_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_2_23_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_2_23_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_2_23_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_1_23_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_1_23_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_2_23_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_2_23_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_2_24 (
    .io_in_r_data         (pe_mat_2_23_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_2_23_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_2_23_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_2_24_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_2_24_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_2_24_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_1_24_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_1_24_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_2_24_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_2_24_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_2_25 (
    .io_in_r_data         (pe_mat_2_24_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_2_24_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_2_24_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_2_25_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_2_25_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_2_25_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_1_25_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_1_25_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_2_25_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_2_25_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_2_26 (
    .io_in_r_data         (pe_mat_2_25_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_2_25_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_2_25_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_2_26_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_2_26_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_2_26_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_1_26_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_1_26_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_2_26_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_2_26_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_2_27 (
    .io_in_r_data         (pe_mat_2_26_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_2_26_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_2_26_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_2_27_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_2_27_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_2_27_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_1_27_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_1_27_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_2_27_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_2_27_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_2_28 (
    .io_in_r_data         (pe_mat_2_27_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_2_27_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_2_27_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_2_28_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_2_28_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_2_28_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_1_28_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_1_28_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_2_28_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_2_28_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_2_29 (
    .io_in_r_data         (pe_mat_2_28_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_2_28_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_2_28_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_2_29_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_2_29_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_2_29_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_1_29_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_1_29_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_2_29_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_2_29_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_2_30 (
    .io_in_r_data         (pe_mat_2_29_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_2_29_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_2_29_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_2_30_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_2_30_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_2_30_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_1_30_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_1_30_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_2_30_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_2_30_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_2_31 (
    .io_in_r_data         (pe_mat_2_30_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_2_30_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_2_30_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_2_31_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_2_31_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_2_31_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_1_31_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_1_31_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_2_31_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_2_31_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_3_0 (
    .io_in_r_data         (io_in_r_3_data[15:0]           ), //i
    .io_in_r_stop_weight  (io_in_r_3_stop_weight          ), //i
    .io_in_r_stall        (io_in_r_3_stall                ), //i
    .io_out_r_data        (pe_mat_3_0_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_3_0_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_3_0_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_2_0_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_2_0_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_3_0_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_3_0_io_out_c_is_weight  ), //o
    .clk                  (clk                            ), //i
    .reset                (reset                          )  //i
  );
  PEWS_1023 pe_mat_3_1 (
    .io_in_r_data         (pe_mat_3_0_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_3_0_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_3_0_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_3_1_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_3_1_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_3_1_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_2_1_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_2_1_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_3_1_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_3_1_io_out_c_is_weight  ), //o
    .clk                  (clk                            ), //i
    .reset                (reset                          )  //i
  );
  PEWS_1023 pe_mat_3_2 (
    .io_in_r_data         (pe_mat_3_1_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_3_1_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_3_1_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_3_2_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_3_2_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_3_2_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_2_2_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_2_2_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_3_2_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_3_2_io_out_c_is_weight  ), //o
    .clk                  (clk                            ), //i
    .reset                (reset                          )  //i
  );
  PEWS_1023 pe_mat_3_3 (
    .io_in_r_data         (pe_mat_3_2_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_3_2_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_3_2_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_3_3_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_3_3_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_3_3_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_2_3_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_2_3_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_3_3_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_3_3_io_out_c_is_weight  ), //o
    .clk                  (clk                            ), //i
    .reset                (reset                          )  //i
  );
  PEWS_1023 pe_mat_3_4 (
    .io_in_r_data         (pe_mat_3_3_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_3_3_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_3_3_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_3_4_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_3_4_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_3_4_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_2_4_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_2_4_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_3_4_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_3_4_io_out_c_is_weight  ), //o
    .clk                  (clk                            ), //i
    .reset                (reset                          )  //i
  );
  PEWS_1023 pe_mat_3_5 (
    .io_in_r_data         (pe_mat_3_4_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_3_4_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_3_4_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_3_5_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_3_5_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_3_5_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_2_5_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_2_5_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_3_5_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_3_5_io_out_c_is_weight  ), //o
    .clk                  (clk                            ), //i
    .reset                (reset                          )  //i
  );
  PEWS_1023 pe_mat_3_6 (
    .io_in_r_data         (pe_mat_3_5_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_3_5_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_3_5_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_3_6_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_3_6_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_3_6_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_2_6_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_2_6_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_3_6_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_3_6_io_out_c_is_weight  ), //o
    .clk                  (clk                            ), //i
    .reset                (reset                          )  //i
  );
  PEWS_1023 pe_mat_3_7 (
    .io_in_r_data         (pe_mat_3_6_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_3_6_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_3_6_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_3_7_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_3_7_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_3_7_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_2_7_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_2_7_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_3_7_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_3_7_io_out_c_is_weight  ), //o
    .clk                  (clk                            ), //i
    .reset                (reset                          )  //i
  );
  PEWS_1023 pe_mat_3_8 (
    .io_in_r_data         (pe_mat_3_7_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_3_7_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_3_7_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_3_8_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_3_8_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_3_8_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_2_8_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_2_8_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_3_8_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_3_8_io_out_c_is_weight  ), //o
    .clk                  (clk                            ), //i
    .reset                (reset                          )  //i
  );
  PEWS_1023 pe_mat_3_9 (
    .io_in_r_data         (pe_mat_3_8_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_3_8_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_3_8_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_3_9_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_3_9_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_3_9_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_2_9_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_2_9_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_3_9_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_3_9_io_out_c_is_weight  ), //o
    .clk                  (clk                            ), //i
    .reset                (reset                          )  //i
  );
  PEWS_1023 pe_mat_3_10 (
    .io_in_r_data         (pe_mat_3_9_io_out_r_data[15:0]  ), //i
    .io_in_r_stop_weight  (pe_mat_3_9_io_out_r_stop_weight ), //i
    .io_in_r_stall        (pe_mat_3_9_io_out_r_stall       ), //i
    .io_out_r_data        (pe_mat_3_10_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_3_10_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_3_10_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_2_10_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_2_10_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_3_10_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_3_10_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_3_11 (
    .io_in_r_data         (pe_mat_3_10_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_3_10_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_3_10_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_3_11_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_3_11_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_3_11_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_2_11_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_2_11_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_3_11_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_3_11_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_3_12 (
    .io_in_r_data         (pe_mat_3_11_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_3_11_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_3_11_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_3_12_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_3_12_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_3_12_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_2_12_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_2_12_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_3_12_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_3_12_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_3_13 (
    .io_in_r_data         (pe_mat_3_12_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_3_12_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_3_12_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_3_13_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_3_13_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_3_13_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_2_13_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_2_13_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_3_13_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_3_13_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_3_14 (
    .io_in_r_data         (pe_mat_3_13_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_3_13_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_3_13_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_3_14_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_3_14_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_3_14_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_2_14_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_2_14_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_3_14_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_3_14_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_3_15 (
    .io_in_r_data         (pe_mat_3_14_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_3_14_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_3_14_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_3_15_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_3_15_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_3_15_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_2_15_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_2_15_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_3_15_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_3_15_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_3_16 (
    .io_in_r_data         (pe_mat_3_15_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_3_15_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_3_15_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_3_16_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_3_16_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_3_16_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_2_16_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_2_16_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_3_16_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_3_16_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_3_17 (
    .io_in_r_data         (pe_mat_3_16_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_3_16_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_3_16_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_3_17_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_3_17_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_3_17_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_2_17_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_2_17_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_3_17_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_3_17_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_3_18 (
    .io_in_r_data         (pe_mat_3_17_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_3_17_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_3_17_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_3_18_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_3_18_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_3_18_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_2_18_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_2_18_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_3_18_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_3_18_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_3_19 (
    .io_in_r_data         (pe_mat_3_18_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_3_18_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_3_18_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_3_19_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_3_19_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_3_19_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_2_19_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_2_19_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_3_19_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_3_19_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_3_20 (
    .io_in_r_data         (pe_mat_3_19_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_3_19_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_3_19_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_3_20_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_3_20_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_3_20_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_2_20_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_2_20_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_3_20_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_3_20_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_3_21 (
    .io_in_r_data         (pe_mat_3_20_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_3_20_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_3_20_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_3_21_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_3_21_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_3_21_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_2_21_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_2_21_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_3_21_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_3_21_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_3_22 (
    .io_in_r_data         (pe_mat_3_21_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_3_21_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_3_21_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_3_22_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_3_22_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_3_22_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_2_22_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_2_22_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_3_22_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_3_22_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_3_23 (
    .io_in_r_data         (pe_mat_3_22_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_3_22_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_3_22_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_3_23_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_3_23_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_3_23_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_2_23_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_2_23_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_3_23_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_3_23_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_3_24 (
    .io_in_r_data         (pe_mat_3_23_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_3_23_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_3_23_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_3_24_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_3_24_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_3_24_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_2_24_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_2_24_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_3_24_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_3_24_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_3_25 (
    .io_in_r_data         (pe_mat_3_24_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_3_24_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_3_24_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_3_25_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_3_25_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_3_25_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_2_25_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_2_25_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_3_25_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_3_25_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_3_26 (
    .io_in_r_data         (pe_mat_3_25_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_3_25_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_3_25_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_3_26_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_3_26_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_3_26_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_2_26_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_2_26_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_3_26_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_3_26_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_3_27 (
    .io_in_r_data         (pe_mat_3_26_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_3_26_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_3_26_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_3_27_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_3_27_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_3_27_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_2_27_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_2_27_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_3_27_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_3_27_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_3_28 (
    .io_in_r_data         (pe_mat_3_27_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_3_27_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_3_27_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_3_28_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_3_28_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_3_28_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_2_28_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_2_28_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_3_28_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_3_28_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_3_29 (
    .io_in_r_data         (pe_mat_3_28_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_3_28_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_3_28_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_3_29_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_3_29_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_3_29_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_2_29_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_2_29_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_3_29_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_3_29_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_3_30 (
    .io_in_r_data         (pe_mat_3_29_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_3_29_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_3_29_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_3_30_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_3_30_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_3_30_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_2_30_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_2_30_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_3_30_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_3_30_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_3_31 (
    .io_in_r_data         (pe_mat_3_30_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_3_30_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_3_30_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_3_31_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_3_31_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_3_31_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_2_31_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_2_31_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_3_31_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_3_31_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_4_0 (
    .io_in_r_data         (io_in_r_4_data[15:0]           ), //i
    .io_in_r_stop_weight  (io_in_r_4_stop_weight          ), //i
    .io_in_r_stall        (io_in_r_4_stall                ), //i
    .io_out_r_data        (pe_mat_4_0_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_4_0_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_4_0_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_3_0_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_3_0_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_4_0_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_4_0_io_out_c_is_weight  ), //o
    .clk                  (clk                            ), //i
    .reset                (reset                          )  //i
  );
  PEWS_1023 pe_mat_4_1 (
    .io_in_r_data         (pe_mat_4_0_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_4_0_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_4_0_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_4_1_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_4_1_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_4_1_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_3_1_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_3_1_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_4_1_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_4_1_io_out_c_is_weight  ), //o
    .clk                  (clk                            ), //i
    .reset                (reset                          )  //i
  );
  PEWS_1023 pe_mat_4_2 (
    .io_in_r_data         (pe_mat_4_1_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_4_1_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_4_1_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_4_2_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_4_2_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_4_2_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_3_2_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_3_2_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_4_2_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_4_2_io_out_c_is_weight  ), //o
    .clk                  (clk                            ), //i
    .reset                (reset                          )  //i
  );
  PEWS_1023 pe_mat_4_3 (
    .io_in_r_data         (pe_mat_4_2_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_4_2_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_4_2_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_4_3_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_4_3_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_4_3_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_3_3_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_3_3_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_4_3_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_4_3_io_out_c_is_weight  ), //o
    .clk                  (clk                            ), //i
    .reset                (reset                          )  //i
  );
  PEWS_1023 pe_mat_4_4 (
    .io_in_r_data         (pe_mat_4_3_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_4_3_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_4_3_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_4_4_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_4_4_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_4_4_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_3_4_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_3_4_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_4_4_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_4_4_io_out_c_is_weight  ), //o
    .clk                  (clk                            ), //i
    .reset                (reset                          )  //i
  );
  PEWS_1023 pe_mat_4_5 (
    .io_in_r_data         (pe_mat_4_4_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_4_4_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_4_4_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_4_5_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_4_5_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_4_5_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_3_5_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_3_5_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_4_5_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_4_5_io_out_c_is_weight  ), //o
    .clk                  (clk                            ), //i
    .reset                (reset                          )  //i
  );
  PEWS_1023 pe_mat_4_6 (
    .io_in_r_data         (pe_mat_4_5_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_4_5_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_4_5_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_4_6_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_4_6_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_4_6_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_3_6_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_3_6_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_4_6_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_4_6_io_out_c_is_weight  ), //o
    .clk                  (clk                            ), //i
    .reset                (reset                          )  //i
  );
  PEWS_1023 pe_mat_4_7 (
    .io_in_r_data         (pe_mat_4_6_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_4_6_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_4_6_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_4_7_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_4_7_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_4_7_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_3_7_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_3_7_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_4_7_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_4_7_io_out_c_is_weight  ), //o
    .clk                  (clk                            ), //i
    .reset                (reset                          )  //i
  );
  PEWS_1023 pe_mat_4_8 (
    .io_in_r_data         (pe_mat_4_7_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_4_7_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_4_7_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_4_8_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_4_8_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_4_8_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_3_8_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_3_8_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_4_8_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_4_8_io_out_c_is_weight  ), //o
    .clk                  (clk                            ), //i
    .reset                (reset                          )  //i
  );
  PEWS_1023 pe_mat_4_9 (
    .io_in_r_data         (pe_mat_4_8_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_4_8_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_4_8_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_4_9_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_4_9_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_4_9_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_3_9_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_3_9_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_4_9_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_4_9_io_out_c_is_weight  ), //o
    .clk                  (clk                            ), //i
    .reset                (reset                          )  //i
  );
  PEWS_1023 pe_mat_4_10 (
    .io_in_r_data         (pe_mat_4_9_io_out_r_data[15:0]  ), //i
    .io_in_r_stop_weight  (pe_mat_4_9_io_out_r_stop_weight ), //i
    .io_in_r_stall        (pe_mat_4_9_io_out_r_stall       ), //i
    .io_out_r_data        (pe_mat_4_10_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_4_10_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_4_10_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_3_10_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_3_10_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_4_10_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_4_10_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_4_11 (
    .io_in_r_data         (pe_mat_4_10_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_4_10_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_4_10_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_4_11_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_4_11_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_4_11_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_3_11_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_3_11_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_4_11_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_4_11_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_4_12 (
    .io_in_r_data         (pe_mat_4_11_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_4_11_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_4_11_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_4_12_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_4_12_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_4_12_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_3_12_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_3_12_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_4_12_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_4_12_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_4_13 (
    .io_in_r_data         (pe_mat_4_12_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_4_12_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_4_12_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_4_13_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_4_13_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_4_13_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_3_13_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_3_13_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_4_13_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_4_13_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_4_14 (
    .io_in_r_data         (pe_mat_4_13_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_4_13_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_4_13_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_4_14_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_4_14_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_4_14_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_3_14_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_3_14_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_4_14_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_4_14_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_4_15 (
    .io_in_r_data         (pe_mat_4_14_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_4_14_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_4_14_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_4_15_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_4_15_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_4_15_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_3_15_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_3_15_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_4_15_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_4_15_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_4_16 (
    .io_in_r_data         (pe_mat_4_15_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_4_15_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_4_15_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_4_16_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_4_16_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_4_16_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_3_16_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_3_16_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_4_16_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_4_16_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_4_17 (
    .io_in_r_data         (pe_mat_4_16_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_4_16_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_4_16_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_4_17_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_4_17_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_4_17_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_3_17_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_3_17_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_4_17_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_4_17_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_4_18 (
    .io_in_r_data         (pe_mat_4_17_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_4_17_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_4_17_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_4_18_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_4_18_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_4_18_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_3_18_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_3_18_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_4_18_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_4_18_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_4_19 (
    .io_in_r_data         (pe_mat_4_18_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_4_18_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_4_18_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_4_19_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_4_19_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_4_19_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_3_19_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_3_19_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_4_19_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_4_19_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_4_20 (
    .io_in_r_data         (pe_mat_4_19_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_4_19_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_4_19_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_4_20_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_4_20_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_4_20_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_3_20_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_3_20_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_4_20_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_4_20_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_4_21 (
    .io_in_r_data         (pe_mat_4_20_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_4_20_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_4_20_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_4_21_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_4_21_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_4_21_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_3_21_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_3_21_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_4_21_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_4_21_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_4_22 (
    .io_in_r_data         (pe_mat_4_21_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_4_21_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_4_21_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_4_22_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_4_22_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_4_22_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_3_22_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_3_22_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_4_22_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_4_22_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_4_23 (
    .io_in_r_data         (pe_mat_4_22_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_4_22_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_4_22_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_4_23_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_4_23_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_4_23_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_3_23_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_3_23_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_4_23_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_4_23_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_4_24 (
    .io_in_r_data         (pe_mat_4_23_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_4_23_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_4_23_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_4_24_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_4_24_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_4_24_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_3_24_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_3_24_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_4_24_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_4_24_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_4_25 (
    .io_in_r_data         (pe_mat_4_24_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_4_24_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_4_24_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_4_25_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_4_25_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_4_25_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_3_25_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_3_25_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_4_25_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_4_25_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_4_26 (
    .io_in_r_data         (pe_mat_4_25_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_4_25_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_4_25_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_4_26_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_4_26_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_4_26_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_3_26_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_3_26_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_4_26_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_4_26_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_4_27 (
    .io_in_r_data         (pe_mat_4_26_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_4_26_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_4_26_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_4_27_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_4_27_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_4_27_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_3_27_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_3_27_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_4_27_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_4_27_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_4_28 (
    .io_in_r_data         (pe_mat_4_27_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_4_27_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_4_27_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_4_28_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_4_28_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_4_28_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_3_28_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_3_28_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_4_28_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_4_28_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_4_29 (
    .io_in_r_data         (pe_mat_4_28_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_4_28_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_4_28_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_4_29_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_4_29_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_4_29_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_3_29_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_3_29_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_4_29_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_4_29_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_4_30 (
    .io_in_r_data         (pe_mat_4_29_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_4_29_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_4_29_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_4_30_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_4_30_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_4_30_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_3_30_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_3_30_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_4_30_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_4_30_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_4_31 (
    .io_in_r_data         (pe_mat_4_30_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_4_30_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_4_30_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_4_31_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_4_31_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_4_31_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_3_31_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_3_31_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_4_31_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_4_31_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_5_0 (
    .io_in_r_data         (io_in_r_5_data[15:0]           ), //i
    .io_in_r_stop_weight  (io_in_r_5_stop_weight          ), //i
    .io_in_r_stall        (io_in_r_5_stall                ), //i
    .io_out_r_data        (pe_mat_5_0_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_5_0_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_5_0_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_4_0_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_4_0_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_5_0_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_5_0_io_out_c_is_weight  ), //o
    .clk                  (clk                            ), //i
    .reset                (reset                          )  //i
  );
  PEWS_1023 pe_mat_5_1 (
    .io_in_r_data         (pe_mat_5_0_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_5_0_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_5_0_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_5_1_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_5_1_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_5_1_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_4_1_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_4_1_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_5_1_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_5_1_io_out_c_is_weight  ), //o
    .clk                  (clk                            ), //i
    .reset                (reset                          )  //i
  );
  PEWS_1023 pe_mat_5_2 (
    .io_in_r_data         (pe_mat_5_1_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_5_1_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_5_1_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_5_2_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_5_2_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_5_2_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_4_2_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_4_2_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_5_2_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_5_2_io_out_c_is_weight  ), //o
    .clk                  (clk                            ), //i
    .reset                (reset                          )  //i
  );
  PEWS_1023 pe_mat_5_3 (
    .io_in_r_data         (pe_mat_5_2_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_5_2_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_5_2_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_5_3_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_5_3_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_5_3_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_4_3_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_4_3_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_5_3_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_5_3_io_out_c_is_weight  ), //o
    .clk                  (clk                            ), //i
    .reset                (reset                          )  //i
  );
  PEWS_1023 pe_mat_5_4 (
    .io_in_r_data         (pe_mat_5_3_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_5_3_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_5_3_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_5_4_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_5_4_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_5_4_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_4_4_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_4_4_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_5_4_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_5_4_io_out_c_is_weight  ), //o
    .clk                  (clk                            ), //i
    .reset                (reset                          )  //i
  );
  PEWS_1023 pe_mat_5_5 (
    .io_in_r_data         (pe_mat_5_4_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_5_4_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_5_4_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_5_5_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_5_5_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_5_5_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_4_5_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_4_5_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_5_5_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_5_5_io_out_c_is_weight  ), //o
    .clk                  (clk                            ), //i
    .reset                (reset                          )  //i
  );
  PEWS_1023 pe_mat_5_6 (
    .io_in_r_data         (pe_mat_5_5_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_5_5_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_5_5_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_5_6_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_5_6_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_5_6_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_4_6_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_4_6_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_5_6_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_5_6_io_out_c_is_weight  ), //o
    .clk                  (clk                            ), //i
    .reset                (reset                          )  //i
  );
  PEWS_1023 pe_mat_5_7 (
    .io_in_r_data         (pe_mat_5_6_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_5_6_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_5_6_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_5_7_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_5_7_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_5_7_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_4_7_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_4_7_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_5_7_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_5_7_io_out_c_is_weight  ), //o
    .clk                  (clk                            ), //i
    .reset                (reset                          )  //i
  );
  PEWS_1023 pe_mat_5_8 (
    .io_in_r_data         (pe_mat_5_7_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_5_7_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_5_7_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_5_8_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_5_8_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_5_8_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_4_8_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_4_8_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_5_8_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_5_8_io_out_c_is_weight  ), //o
    .clk                  (clk                            ), //i
    .reset                (reset                          )  //i
  );
  PEWS_1023 pe_mat_5_9 (
    .io_in_r_data         (pe_mat_5_8_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_5_8_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_5_8_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_5_9_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_5_9_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_5_9_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_4_9_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_4_9_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_5_9_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_5_9_io_out_c_is_weight  ), //o
    .clk                  (clk                            ), //i
    .reset                (reset                          )  //i
  );
  PEWS_1023 pe_mat_5_10 (
    .io_in_r_data         (pe_mat_5_9_io_out_r_data[15:0]  ), //i
    .io_in_r_stop_weight  (pe_mat_5_9_io_out_r_stop_weight ), //i
    .io_in_r_stall        (pe_mat_5_9_io_out_r_stall       ), //i
    .io_out_r_data        (pe_mat_5_10_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_5_10_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_5_10_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_4_10_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_4_10_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_5_10_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_5_10_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_5_11 (
    .io_in_r_data         (pe_mat_5_10_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_5_10_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_5_10_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_5_11_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_5_11_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_5_11_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_4_11_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_4_11_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_5_11_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_5_11_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_5_12 (
    .io_in_r_data         (pe_mat_5_11_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_5_11_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_5_11_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_5_12_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_5_12_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_5_12_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_4_12_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_4_12_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_5_12_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_5_12_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_5_13 (
    .io_in_r_data         (pe_mat_5_12_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_5_12_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_5_12_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_5_13_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_5_13_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_5_13_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_4_13_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_4_13_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_5_13_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_5_13_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_5_14 (
    .io_in_r_data         (pe_mat_5_13_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_5_13_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_5_13_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_5_14_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_5_14_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_5_14_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_4_14_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_4_14_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_5_14_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_5_14_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_5_15 (
    .io_in_r_data         (pe_mat_5_14_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_5_14_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_5_14_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_5_15_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_5_15_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_5_15_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_4_15_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_4_15_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_5_15_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_5_15_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_5_16 (
    .io_in_r_data         (pe_mat_5_15_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_5_15_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_5_15_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_5_16_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_5_16_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_5_16_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_4_16_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_4_16_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_5_16_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_5_16_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_5_17 (
    .io_in_r_data         (pe_mat_5_16_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_5_16_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_5_16_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_5_17_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_5_17_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_5_17_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_4_17_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_4_17_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_5_17_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_5_17_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_5_18 (
    .io_in_r_data         (pe_mat_5_17_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_5_17_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_5_17_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_5_18_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_5_18_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_5_18_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_4_18_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_4_18_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_5_18_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_5_18_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_5_19 (
    .io_in_r_data         (pe_mat_5_18_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_5_18_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_5_18_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_5_19_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_5_19_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_5_19_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_4_19_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_4_19_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_5_19_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_5_19_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_5_20 (
    .io_in_r_data         (pe_mat_5_19_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_5_19_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_5_19_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_5_20_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_5_20_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_5_20_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_4_20_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_4_20_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_5_20_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_5_20_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_5_21 (
    .io_in_r_data         (pe_mat_5_20_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_5_20_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_5_20_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_5_21_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_5_21_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_5_21_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_4_21_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_4_21_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_5_21_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_5_21_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_5_22 (
    .io_in_r_data         (pe_mat_5_21_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_5_21_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_5_21_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_5_22_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_5_22_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_5_22_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_4_22_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_4_22_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_5_22_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_5_22_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_5_23 (
    .io_in_r_data         (pe_mat_5_22_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_5_22_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_5_22_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_5_23_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_5_23_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_5_23_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_4_23_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_4_23_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_5_23_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_5_23_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_5_24 (
    .io_in_r_data         (pe_mat_5_23_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_5_23_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_5_23_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_5_24_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_5_24_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_5_24_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_4_24_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_4_24_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_5_24_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_5_24_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_5_25 (
    .io_in_r_data         (pe_mat_5_24_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_5_24_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_5_24_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_5_25_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_5_25_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_5_25_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_4_25_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_4_25_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_5_25_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_5_25_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_5_26 (
    .io_in_r_data         (pe_mat_5_25_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_5_25_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_5_25_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_5_26_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_5_26_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_5_26_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_4_26_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_4_26_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_5_26_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_5_26_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_5_27 (
    .io_in_r_data         (pe_mat_5_26_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_5_26_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_5_26_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_5_27_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_5_27_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_5_27_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_4_27_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_4_27_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_5_27_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_5_27_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_5_28 (
    .io_in_r_data         (pe_mat_5_27_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_5_27_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_5_27_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_5_28_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_5_28_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_5_28_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_4_28_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_4_28_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_5_28_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_5_28_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_5_29 (
    .io_in_r_data         (pe_mat_5_28_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_5_28_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_5_28_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_5_29_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_5_29_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_5_29_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_4_29_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_4_29_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_5_29_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_5_29_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_5_30 (
    .io_in_r_data         (pe_mat_5_29_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_5_29_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_5_29_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_5_30_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_5_30_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_5_30_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_4_30_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_4_30_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_5_30_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_5_30_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_5_31 (
    .io_in_r_data         (pe_mat_5_30_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_5_30_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_5_30_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_5_31_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_5_31_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_5_31_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_4_31_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_4_31_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_5_31_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_5_31_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_6_0 (
    .io_in_r_data         (io_in_r_6_data[15:0]           ), //i
    .io_in_r_stop_weight  (io_in_r_6_stop_weight          ), //i
    .io_in_r_stall        (io_in_r_6_stall                ), //i
    .io_out_r_data        (pe_mat_6_0_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_6_0_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_6_0_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_5_0_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_5_0_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_6_0_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_6_0_io_out_c_is_weight  ), //o
    .clk                  (clk                            ), //i
    .reset                (reset                          )  //i
  );
  PEWS_1023 pe_mat_6_1 (
    .io_in_r_data         (pe_mat_6_0_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_6_0_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_6_0_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_6_1_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_6_1_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_6_1_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_5_1_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_5_1_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_6_1_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_6_1_io_out_c_is_weight  ), //o
    .clk                  (clk                            ), //i
    .reset                (reset                          )  //i
  );
  PEWS_1023 pe_mat_6_2 (
    .io_in_r_data         (pe_mat_6_1_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_6_1_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_6_1_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_6_2_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_6_2_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_6_2_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_5_2_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_5_2_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_6_2_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_6_2_io_out_c_is_weight  ), //o
    .clk                  (clk                            ), //i
    .reset                (reset                          )  //i
  );
  PEWS_1023 pe_mat_6_3 (
    .io_in_r_data         (pe_mat_6_2_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_6_2_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_6_2_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_6_3_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_6_3_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_6_3_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_5_3_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_5_3_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_6_3_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_6_3_io_out_c_is_weight  ), //o
    .clk                  (clk                            ), //i
    .reset                (reset                          )  //i
  );
  PEWS_1023 pe_mat_6_4 (
    .io_in_r_data         (pe_mat_6_3_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_6_3_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_6_3_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_6_4_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_6_4_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_6_4_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_5_4_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_5_4_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_6_4_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_6_4_io_out_c_is_weight  ), //o
    .clk                  (clk                            ), //i
    .reset                (reset                          )  //i
  );
  PEWS_1023 pe_mat_6_5 (
    .io_in_r_data         (pe_mat_6_4_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_6_4_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_6_4_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_6_5_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_6_5_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_6_5_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_5_5_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_5_5_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_6_5_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_6_5_io_out_c_is_weight  ), //o
    .clk                  (clk                            ), //i
    .reset                (reset                          )  //i
  );
  PEWS_1023 pe_mat_6_6 (
    .io_in_r_data         (pe_mat_6_5_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_6_5_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_6_5_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_6_6_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_6_6_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_6_6_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_5_6_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_5_6_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_6_6_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_6_6_io_out_c_is_weight  ), //o
    .clk                  (clk                            ), //i
    .reset                (reset                          )  //i
  );
  PEWS_1023 pe_mat_6_7 (
    .io_in_r_data         (pe_mat_6_6_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_6_6_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_6_6_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_6_7_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_6_7_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_6_7_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_5_7_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_5_7_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_6_7_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_6_7_io_out_c_is_weight  ), //o
    .clk                  (clk                            ), //i
    .reset                (reset                          )  //i
  );
  PEWS_1023 pe_mat_6_8 (
    .io_in_r_data         (pe_mat_6_7_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_6_7_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_6_7_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_6_8_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_6_8_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_6_8_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_5_8_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_5_8_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_6_8_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_6_8_io_out_c_is_weight  ), //o
    .clk                  (clk                            ), //i
    .reset                (reset                          )  //i
  );
  PEWS_1023 pe_mat_6_9 (
    .io_in_r_data         (pe_mat_6_8_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_6_8_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_6_8_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_6_9_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_6_9_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_6_9_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_5_9_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_5_9_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_6_9_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_6_9_io_out_c_is_weight  ), //o
    .clk                  (clk                            ), //i
    .reset                (reset                          )  //i
  );
  PEWS_1023 pe_mat_6_10 (
    .io_in_r_data         (pe_mat_6_9_io_out_r_data[15:0]  ), //i
    .io_in_r_stop_weight  (pe_mat_6_9_io_out_r_stop_weight ), //i
    .io_in_r_stall        (pe_mat_6_9_io_out_r_stall       ), //i
    .io_out_r_data        (pe_mat_6_10_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_6_10_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_6_10_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_5_10_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_5_10_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_6_10_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_6_10_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_6_11 (
    .io_in_r_data         (pe_mat_6_10_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_6_10_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_6_10_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_6_11_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_6_11_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_6_11_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_5_11_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_5_11_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_6_11_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_6_11_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_6_12 (
    .io_in_r_data         (pe_mat_6_11_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_6_11_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_6_11_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_6_12_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_6_12_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_6_12_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_5_12_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_5_12_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_6_12_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_6_12_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_6_13 (
    .io_in_r_data         (pe_mat_6_12_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_6_12_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_6_12_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_6_13_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_6_13_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_6_13_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_5_13_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_5_13_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_6_13_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_6_13_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_6_14 (
    .io_in_r_data         (pe_mat_6_13_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_6_13_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_6_13_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_6_14_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_6_14_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_6_14_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_5_14_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_5_14_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_6_14_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_6_14_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_6_15 (
    .io_in_r_data         (pe_mat_6_14_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_6_14_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_6_14_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_6_15_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_6_15_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_6_15_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_5_15_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_5_15_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_6_15_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_6_15_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_6_16 (
    .io_in_r_data         (pe_mat_6_15_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_6_15_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_6_15_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_6_16_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_6_16_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_6_16_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_5_16_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_5_16_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_6_16_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_6_16_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_6_17 (
    .io_in_r_data         (pe_mat_6_16_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_6_16_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_6_16_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_6_17_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_6_17_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_6_17_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_5_17_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_5_17_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_6_17_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_6_17_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_6_18 (
    .io_in_r_data         (pe_mat_6_17_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_6_17_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_6_17_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_6_18_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_6_18_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_6_18_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_5_18_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_5_18_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_6_18_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_6_18_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_6_19 (
    .io_in_r_data         (pe_mat_6_18_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_6_18_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_6_18_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_6_19_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_6_19_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_6_19_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_5_19_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_5_19_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_6_19_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_6_19_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_6_20 (
    .io_in_r_data         (pe_mat_6_19_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_6_19_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_6_19_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_6_20_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_6_20_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_6_20_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_5_20_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_5_20_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_6_20_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_6_20_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_6_21 (
    .io_in_r_data         (pe_mat_6_20_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_6_20_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_6_20_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_6_21_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_6_21_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_6_21_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_5_21_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_5_21_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_6_21_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_6_21_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_6_22 (
    .io_in_r_data         (pe_mat_6_21_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_6_21_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_6_21_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_6_22_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_6_22_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_6_22_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_5_22_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_5_22_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_6_22_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_6_22_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_6_23 (
    .io_in_r_data         (pe_mat_6_22_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_6_22_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_6_22_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_6_23_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_6_23_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_6_23_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_5_23_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_5_23_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_6_23_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_6_23_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_6_24 (
    .io_in_r_data         (pe_mat_6_23_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_6_23_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_6_23_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_6_24_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_6_24_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_6_24_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_5_24_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_5_24_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_6_24_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_6_24_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_6_25 (
    .io_in_r_data         (pe_mat_6_24_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_6_24_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_6_24_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_6_25_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_6_25_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_6_25_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_5_25_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_5_25_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_6_25_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_6_25_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_6_26 (
    .io_in_r_data         (pe_mat_6_25_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_6_25_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_6_25_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_6_26_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_6_26_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_6_26_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_5_26_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_5_26_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_6_26_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_6_26_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_6_27 (
    .io_in_r_data         (pe_mat_6_26_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_6_26_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_6_26_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_6_27_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_6_27_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_6_27_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_5_27_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_5_27_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_6_27_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_6_27_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_6_28 (
    .io_in_r_data         (pe_mat_6_27_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_6_27_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_6_27_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_6_28_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_6_28_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_6_28_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_5_28_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_5_28_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_6_28_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_6_28_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_6_29 (
    .io_in_r_data         (pe_mat_6_28_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_6_28_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_6_28_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_6_29_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_6_29_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_6_29_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_5_29_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_5_29_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_6_29_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_6_29_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_6_30 (
    .io_in_r_data         (pe_mat_6_29_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_6_29_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_6_29_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_6_30_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_6_30_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_6_30_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_5_30_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_5_30_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_6_30_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_6_30_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_6_31 (
    .io_in_r_data         (pe_mat_6_30_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_6_30_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_6_30_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_6_31_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_6_31_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_6_31_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_5_31_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_5_31_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_6_31_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_6_31_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_7_0 (
    .io_in_r_data         (io_in_r_7_data[15:0]           ), //i
    .io_in_r_stop_weight  (io_in_r_7_stop_weight          ), //i
    .io_in_r_stall        (io_in_r_7_stall                ), //i
    .io_out_r_data        (pe_mat_7_0_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_7_0_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_7_0_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_6_0_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_6_0_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_7_0_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_7_0_io_out_c_is_weight  ), //o
    .clk                  (clk                            ), //i
    .reset                (reset                          )  //i
  );
  PEWS_1023 pe_mat_7_1 (
    .io_in_r_data         (pe_mat_7_0_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_7_0_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_7_0_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_7_1_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_7_1_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_7_1_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_6_1_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_6_1_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_7_1_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_7_1_io_out_c_is_weight  ), //o
    .clk                  (clk                            ), //i
    .reset                (reset                          )  //i
  );
  PEWS_1023 pe_mat_7_2 (
    .io_in_r_data         (pe_mat_7_1_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_7_1_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_7_1_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_7_2_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_7_2_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_7_2_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_6_2_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_6_2_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_7_2_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_7_2_io_out_c_is_weight  ), //o
    .clk                  (clk                            ), //i
    .reset                (reset                          )  //i
  );
  PEWS_1023 pe_mat_7_3 (
    .io_in_r_data         (pe_mat_7_2_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_7_2_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_7_2_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_7_3_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_7_3_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_7_3_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_6_3_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_6_3_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_7_3_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_7_3_io_out_c_is_weight  ), //o
    .clk                  (clk                            ), //i
    .reset                (reset                          )  //i
  );
  PEWS_1023 pe_mat_7_4 (
    .io_in_r_data         (pe_mat_7_3_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_7_3_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_7_3_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_7_4_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_7_4_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_7_4_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_6_4_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_6_4_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_7_4_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_7_4_io_out_c_is_weight  ), //o
    .clk                  (clk                            ), //i
    .reset                (reset                          )  //i
  );
  PEWS_1023 pe_mat_7_5 (
    .io_in_r_data         (pe_mat_7_4_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_7_4_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_7_4_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_7_5_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_7_5_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_7_5_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_6_5_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_6_5_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_7_5_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_7_5_io_out_c_is_weight  ), //o
    .clk                  (clk                            ), //i
    .reset                (reset                          )  //i
  );
  PEWS_1023 pe_mat_7_6 (
    .io_in_r_data         (pe_mat_7_5_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_7_5_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_7_5_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_7_6_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_7_6_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_7_6_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_6_6_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_6_6_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_7_6_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_7_6_io_out_c_is_weight  ), //o
    .clk                  (clk                            ), //i
    .reset                (reset                          )  //i
  );
  PEWS_1023 pe_mat_7_7 (
    .io_in_r_data         (pe_mat_7_6_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_7_6_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_7_6_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_7_7_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_7_7_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_7_7_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_6_7_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_6_7_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_7_7_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_7_7_io_out_c_is_weight  ), //o
    .clk                  (clk                            ), //i
    .reset                (reset                          )  //i
  );
  PEWS_1023 pe_mat_7_8 (
    .io_in_r_data         (pe_mat_7_7_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_7_7_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_7_7_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_7_8_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_7_8_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_7_8_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_6_8_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_6_8_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_7_8_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_7_8_io_out_c_is_weight  ), //o
    .clk                  (clk                            ), //i
    .reset                (reset                          )  //i
  );
  PEWS_1023 pe_mat_7_9 (
    .io_in_r_data         (pe_mat_7_8_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_7_8_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_7_8_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_7_9_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_7_9_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_7_9_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_6_9_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_6_9_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_7_9_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_7_9_io_out_c_is_weight  ), //o
    .clk                  (clk                            ), //i
    .reset                (reset                          )  //i
  );
  PEWS_1023 pe_mat_7_10 (
    .io_in_r_data         (pe_mat_7_9_io_out_r_data[15:0]  ), //i
    .io_in_r_stop_weight  (pe_mat_7_9_io_out_r_stop_weight ), //i
    .io_in_r_stall        (pe_mat_7_9_io_out_r_stall       ), //i
    .io_out_r_data        (pe_mat_7_10_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_7_10_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_7_10_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_6_10_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_6_10_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_7_10_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_7_10_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_7_11 (
    .io_in_r_data         (pe_mat_7_10_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_7_10_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_7_10_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_7_11_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_7_11_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_7_11_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_6_11_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_6_11_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_7_11_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_7_11_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_7_12 (
    .io_in_r_data         (pe_mat_7_11_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_7_11_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_7_11_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_7_12_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_7_12_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_7_12_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_6_12_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_6_12_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_7_12_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_7_12_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_7_13 (
    .io_in_r_data         (pe_mat_7_12_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_7_12_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_7_12_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_7_13_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_7_13_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_7_13_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_6_13_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_6_13_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_7_13_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_7_13_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_7_14 (
    .io_in_r_data         (pe_mat_7_13_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_7_13_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_7_13_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_7_14_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_7_14_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_7_14_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_6_14_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_6_14_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_7_14_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_7_14_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_7_15 (
    .io_in_r_data         (pe_mat_7_14_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_7_14_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_7_14_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_7_15_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_7_15_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_7_15_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_6_15_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_6_15_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_7_15_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_7_15_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_7_16 (
    .io_in_r_data         (pe_mat_7_15_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_7_15_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_7_15_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_7_16_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_7_16_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_7_16_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_6_16_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_6_16_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_7_16_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_7_16_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_7_17 (
    .io_in_r_data         (pe_mat_7_16_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_7_16_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_7_16_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_7_17_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_7_17_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_7_17_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_6_17_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_6_17_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_7_17_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_7_17_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_7_18 (
    .io_in_r_data         (pe_mat_7_17_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_7_17_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_7_17_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_7_18_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_7_18_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_7_18_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_6_18_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_6_18_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_7_18_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_7_18_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_7_19 (
    .io_in_r_data         (pe_mat_7_18_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_7_18_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_7_18_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_7_19_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_7_19_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_7_19_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_6_19_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_6_19_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_7_19_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_7_19_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_7_20 (
    .io_in_r_data         (pe_mat_7_19_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_7_19_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_7_19_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_7_20_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_7_20_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_7_20_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_6_20_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_6_20_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_7_20_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_7_20_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_7_21 (
    .io_in_r_data         (pe_mat_7_20_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_7_20_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_7_20_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_7_21_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_7_21_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_7_21_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_6_21_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_6_21_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_7_21_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_7_21_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_7_22 (
    .io_in_r_data         (pe_mat_7_21_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_7_21_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_7_21_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_7_22_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_7_22_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_7_22_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_6_22_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_6_22_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_7_22_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_7_22_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_7_23 (
    .io_in_r_data         (pe_mat_7_22_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_7_22_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_7_22_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_7_23_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_7_23_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_7_23_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_6_23_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_6_23_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_7_23_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_7_23_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_7_24 (
    .io_in_r_data         (pe_mat_7_23_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_7_23_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_7_23_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_7_24_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_7_24_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_7_24_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_6_24_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_6_24_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_7_24_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_7_24_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_7_25 (
    .io_in_r_data         (pe_mat_7_24_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_7_24_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_7_24_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_7_25_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_7_25_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_7_25_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_6_25_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_6_25_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_7_25_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_7_25_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_7_26 (
    .io_in_r_data         (pe_mat_7_25_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_7_25_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_7_25_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_7_26_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_7_26_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_7_26_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_6_26_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_6_26_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_7_26_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_7_26_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_7_27 (
    .io_in_r_data         (pe_mat_7_26_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_7_26_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_7_26_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_7_27_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_7_27_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_7_27_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_6_27_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_6_27_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_7_27_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_7_27_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_7_28 (
    .io_in_r_data         (pe_mat_7_27_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_7_27_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_7_27_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_7_28_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_7_28_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_7_28_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_6_28_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_6_28_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_7_28_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_7_28_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_7_29 (
    .io_in_r_data         (pe_mat_7_28_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_7_28_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_7_28_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_7_29_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_7_29_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_7_29_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_6_29_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_6_29_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_7_29_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_7_29_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_7_30 (
    .io_in_r_data         (pe_mat_7_29_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_7_29_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_7_29_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_7_30_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_7_30_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_7_30_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_6_30_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_6_30_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_7_30_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_7_30_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_7_31 (
    .io_in_r_data         (pe_mat_7_30_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_7_30_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_7_30_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_7_31_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_7_31_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_7_31_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_6_31_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_6_31_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_7_31_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_7_31_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_8_0 (
    .io_in_r_data         (io_in_r_8_data[15:0]           ), //i
    .io_in_r_stop_weight  (io_in_r_8_stop_weight          ), //i
    .io_in_r_stall        (io_in_r_8_stall                ), //i
    .io_out_r_data        (pe_mat_8_0_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_8_0_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_8_0_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_7_0_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_7_0_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_8_0_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_8_0_io_out_c_is_weight  ), //o
    .clk                  (clk                            ), //i
    .reset                (reset                          )  //i
  );
  PEWS_1023 pe_mat_8_1 (
    .io_in_r_data         (pe_mat_8_0_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_8_0_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_8_0_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_8_1_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_8_1_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_8_1_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_7_1_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_7_1_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_8_1_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_8_1_io_out_c_is_weight  ), //o
    .clk                  (clk                            ), //i
    .reset                (reset                          )  //i
  );
  PEWS_1023 pe_mat_8_2 (
    .io_in_r_data         (pe_mat_8_1_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_8_1_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_8_1_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_8_2_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_8_2_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_8_2_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_7_2_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_7_2_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_8_2_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_8_2_io_out_c_is_weight  ), //o
    .clk                  (clk                            ), //i
    .reset                (reset                          )  //i
  );
  PEWS_1023 pe_mat_8_3 (
    .io_in_r_data         (pe_mat_8_2_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_8_2_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_8_2_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_8_3_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_8_3_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_8_3_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_7_3_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_7_3_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_8_3_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_8_3_io_out_c_is_weight  ), //o
    .clk                  (clk                            ), //i
    .reset                (reset                          )  //i
  );
  PEWS_1023 pe_mat_8_4 (
    .io_in_r_data         (pe_mat_8_3_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_8_3_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_8_3_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_8_4_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_8_4_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_8_4_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_7_4_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_7_4_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_8_4_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_8_4_io_out_c_is_weight  ), //o
    .clk                  (clk                            ), //i
    .reset                (reset                          )  //i
  );
  PEWS_1023 pe_mat_8_5 (
    .io_in_r_data         (pe_mat_8_4_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_8_4_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_8_4_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_8_5_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_8_5_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_8_5_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_7_5_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_7_5_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_8_5_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_8_5_io_out_c_is_weight  ), //o
    .clk                  (clk                            ), //i
    .reset                (reset                          )  //i
  );
  PEWS_1023 pe_mat_8_6 (
    .io_in_r_data         (pe_mat_8_5_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_8_5_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_8_5_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_8_6_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_8_6_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_8_6_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_7_6_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_7_6_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_8_6_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_8_6_io_out_c_is_weight  ), //o
    .clk                  (clk                            ), //i
    .reset                (reset                          )  //i
  );
  PEWS_1023 pe_mat_8_7 (
    .io_in_r_data         (pe_mat_8_6_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_8_6_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_8_6_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_8_7_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_8_7_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_8_7_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_7_7_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_7_7_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_8_7_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_8_7_io_out_c_is_weight  ), //o
    .clk                  (clk                            ), //i
    .reset                (reset                          )  //i
  );
  PEWS_1023 pe_mat_8_8 (
    .io_in_r_data         (pe_mat_8_7_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_8_7_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_8_7_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_8_8_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_8_8_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_8_8_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_7_8_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_7_8_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_8_8_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_8_8_io_out_c_is_weight  ), //o
    .clk                  (clk                            ), //i
    .reset                (reset                          )  //i
  );
  PEWS_1023 pe_mat_8_9 (
    .io_in_r_data         (pe_mat_8_8_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_8_8_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_8_8_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_8_9_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_8_9_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_8_9_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_7_9_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_7_9_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_8_9_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_8_9_io_out_c_is_weight  ), //o
    .clk                  (clk                            ), //i
    .reset                (reset                          )  //i
  );
  PEWS_1023 pe_mat_8_10 (
    .io_in_r_data         (pe_mat_8_9_io_out_r_data[15:0]  ), //i
    .io_in_r_stop_weight  (pe_mat_8_9_io_out_r_stop_weight ), //i
    .io_in_r_stall        (pe_mat_8_9_io_out_r_stall       ), //i
    .io_out_r_data        (pe_mat_8_10_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_8_10_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_8_10_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_7_10_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_7_10_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_8_10_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_8_10_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_8_11 (
    .io_in_r_data         (pe_mat_8_10_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_8_10_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_8_10_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_8_11_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_8_11_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_8_11_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_7_11_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_7_11_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_8_11_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_8_11_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_8_12 (
    .io_in_r_data         (pe_mat_8_11_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_8_11_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_8_11_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_8_12_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_8_12_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_8_12_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_7_12_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_7_12_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_8_12_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_8_12_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_8_13 (
    .io_in_r_data         (pe_mat_8_12_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_8_12_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_8_12_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_8_13_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_8_13_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_8_13_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_7_13_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_7_13_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_8_13_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_8_13_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_8_14 (
    .io_in_r_data         (pe_mat_8_13_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_8_13_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_8_13_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_8_14_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_8_14_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_8_14_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_7_14_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_7_14_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_8_14_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_8_14_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_8_15 (
    .io_in_r_data         (pe_mat_8_14_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_8_14_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_8_14_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_8_15_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_8_15_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_8_15_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_7_15_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_7_15_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_8_15_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_8_15_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_8_16 (
    .io_in_r_data         (pe_mat_8_15_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_8_15_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_8_15_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_8_16_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_8_16_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_8_16_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_7_16_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_7_16_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_8_16_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_8_16_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_8_17 (
    .io_in_r_data         (pe_mat_8_16_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_8_16_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_8_16_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_8_17_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_8_17_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_8_17_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_7_17_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_7_17_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_8_17_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_8_17_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_8_18 (
    .io_in_r_data         (pe_mat_8_17_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_8_17_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_8_17_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_8_18_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_8_18_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_8_18_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_7_18_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_7_18_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_8_18_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_8_18_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_8_19 (
    .io_in_r_data         (pe_mat_8_18_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_8_18_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_8_18_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_8_19_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_8_19_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_8_19_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_7_19_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_7_19_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_8_19_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_8_19_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_8_20 (
    .io_in_r_data         (pe_mat_8_19_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_8_19_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_8_19_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_8_20_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_8_20_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_8_20_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_7_20_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_7_20_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_8_20_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_8_20_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_8_21 (
    .io_in_r_data         (pe_mat_8_20_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_8_20_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_8_20_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_8_21_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_8_21_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_8_21_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_7_21_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_7_21_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_8_21_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_8_21_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_8_22 (
    .io_in_r_data         (pe_mat_8_21_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_8_21_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_8_21_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_8_22_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_8_22_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_8_22_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_7_22_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_7_22_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_8_22_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_8_22_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_8_23 (
    .io_in_r_data         (pe_mat_8_22_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_8_22_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_8_22_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_8_23_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_8_23_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_8_23_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_7_23_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_7_23_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_8_23_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_8_23_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_8_24 (
    .io_in_r_data         (pe_mat_8_23_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_8_23_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_8_23_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_8_24_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_8_24_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_8_24_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_7_24_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_7_24_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_8_24_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_8_24_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_8_25 (
    .io_in_r_data         (pe_mat_8_24_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_8_24_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_8_24_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_8_25_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_8_25_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_8_25_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_7_25_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_7_25_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_8_25_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_8_25_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_8_26 (
    .io_in_r_data         (pe_mat_8_25_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_8_25_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_8_25_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_8_26_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_8_26_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_8_26_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_7_26_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_7_26_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_8_26_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_8_26_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_8_27 (
    .io_in_r_data         (pe_mat_8_26_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_8_26_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_8_26_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_8_27_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_8_27_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_8_27_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_7_27_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_7_27_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_8_27_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_8_27_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_8_28 (
    .io_in_r_data         (pe_mat_8_27_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_8_27_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_8_27_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_8_28_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_8_28_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_8_28_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_7_28_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_7_28_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_8_28_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_8_28_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_8_29 (
    .io_in_r_data         (pe_mat_8_28_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_8_28_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_8_28_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_8_29_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_8_29_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_8_29_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_7_29_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_7_29_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_8_29_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_8_29_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_8_30 (
    .io_in_r_data         (pe_mat_8_29_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_8_29_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_8_29_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_8_30_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_8_30_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_8_30_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_7_30_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_7_30_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_8_30_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_8_30_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_8_31 (
    .io_in_r_data         (pe_mat_8_30_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_8_30_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_8_30_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_8_31_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_8_31_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_8_31_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_7_31_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_7_31_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_8_31_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_8_31_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_9_0 (
    .io_in_r_data         (io_in_r_9_data[15:0]           ), //i
    .io_in_r_stop_weight  (io_in_r_9_stop_weight          ), //i
    .io_in_r_stall        (io_in_r_9_stall                ), //i
    .io_out_r_data        (pe_mat_9_0_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_9_0_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_9_0_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_8_0_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_8_0_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_9_0_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_9_0_io_out_c_is_weight  ), //o
    .clk                  (clk                            ), //i
    .reset                (reset                          )  //i
  );
  PEWS_1023 pe_mat_9_1 (
    .io_in_r_data         (pe_mat_9_0_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_9_0_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_9_0_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_9_1_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_9_1_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_9_1_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_8_1_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_8_1_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_9_1_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_9_1_io_out_c_is_weight  ), //o
    .clk                  (clk                            ), //i
    .reset                (reset                          )  //i
  );
  PEWS_1023 pe_mat_9_2 (
    .io_in_r_data         (pe_mat_9_1_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_9_1_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_9_1_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_9_2_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_9_2_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_9_2_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_8_2_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_8_2_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_9_2_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_9_2_io_out_c_is_weight  ), //o
    .clk                  (clk                            ), //i
    .reset                (reset                          )  //i
  );
  PEWS_1023 pe_mat_9_3 (
    .io_in_r_data         (pe_mat_9_2_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_9_2_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_9_2_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_9_3_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_9_3_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_9_3_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_8_3_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_8_3_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_9_3_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_9_3_io_out_c_is_weight  ), //o
    .clk                  (clk                            ), //i
    .reset                (reset                          )  //i
  );
  PEWS_1023 pe_mat_9_4 (
    .io_in_r_data         (pe_mat_9_3_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_9_3_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_9_3_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_9_4_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_9_4_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_9_4_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_8_4_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_8_4_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_9_4_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_9_4_io_out_c_is_weight  ), //o
    .clk                  (clk                            ), //i
    .reset                (reset                          )  //i
  );
  PEWS_1023 pe_mat_9_5 (
    .io_in_r_data         (pe_mat_9_4_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_9_4_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_9_4_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_9_5_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_9_5_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_9_5_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_8_5_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_8_5_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_9_5_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_9_5_io_out_c_is_weight  ), //o
    .clk                  (clk                            ), //i
    .reset                (reset                          )  //i
  );
  PEWS_1023 pe_mat_9_6 (
    .io_in_r_data         (pe_mat_9_5_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_9_5_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_9_5_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_9_6_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_9_6_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_9_6_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_8_6_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_8_6_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_9_6_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_9_6_io_out_c_is_weight  ), //o
    .clk                  (clk                            ), //i
    .reset                (reset                          )  //i
  );
  PEWS_1023 pe_mat_9_7 (
    .io_in_r_data         (pe_mat_9_6_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_9_6_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_9_6_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_9_7_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_9_7_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_9_7_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_8_7_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_8_7_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_9_7_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_9_7_io_out_c_is_weight  ), //o
    .clk                  (clk                            ), //i
    .reset                (reset                          )  //i
  );
  PEWS_1023 pe_mat_9_8 (
    .io_in_r_data         (pe_mat_9_7_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_9_7_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_9_7_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_9_8_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_9_8_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_9_8_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_8_8_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_8_8_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_9_8_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_9_8_io_out_c_is_weight  ), //o
    .clk                  (clk                            ), //i
    .reset                (reset                          )  //i
  );
  PEWS_1023 pe_mat_9_9 (
    .io_in_r_data         (pe_mat_9_8_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_9_8_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_9_8_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_9_9_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_9_9_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_9_9_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_8_9_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_8_9_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_9_9_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_9_9_io_out_c_is_weight  ), //o
    .clk                  (clk                            ), //i
    .reset                (reset                          )  //i
  );
  PEWS_1023 pe_mat_9_10 (
    .io_in_r_data         (pe_mat_9_9_io_out_r_data[15:0]  ), //i
    .io_in_r_stop_weight  (pe_mat_9_9_io_out_r_stop_weight ), //i
    .io_in_r_stall        (pe_mat_9_9_io_out_r_stall       ), //i
    .io_out_r_data        (pe_mat_9_10_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_9_10_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_9_10_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_8_10_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_8_10_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_9_10_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_9_10_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_9_11 (
    .io_in_r_data         (pe_mat_9_10_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_9_10_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_9_10_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_9_11_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_9_11_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_9_11_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_8_11_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_8_11_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_9_11_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_9_11_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_9_12 (
    .io_in_r_data         (pe_mat_9_11_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_9_11_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_9_11_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_9_12_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_9_12_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_9_12_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_8_12_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_8_12_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_9_12_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_9_12_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_9_13 (
    .io_in_r_data         (pe_mat_9_12_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_9_12_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_9_12_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_9_13_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_9_13_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_9_13_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_8_13_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_8_13_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_9_13_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_9_13_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_9_14 (
    .io_in_r_data         (pe_mat_9_13_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_9_13_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_9_13_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_9_14_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_9_14_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_9_14_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_8_14_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_8_14_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_9_14_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_9_14_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_9_15 (
    .io_in_r_data         (pe_mat_9_14_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_9_14_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_9_14_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_9_15_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_9_15_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_9_15_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_8_15_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_8_15_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_9_15_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_9_15_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_9_16 (
    .io_in_r_data         (pe_mat_9_15_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_9_15_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_9_15_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_9_16_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_9_16_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_9_16_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_8_16_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_8_16_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_9_16_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_9_16_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_9_17 (
    .io_in_r_data         (pe_mat_9_16_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_9_16_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_9_16_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_9_17_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_9_17_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_9_17_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_8_17_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_8_17_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_9_17_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_9_17_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_9_18 (
    .io_in_r_data         (pe_mat_9_17_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_9_17_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_9_17_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_9_18_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_9_18_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_9_18_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_8_18_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_8_18_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_9_18_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_9_18_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_9_19 (
    .io_in_r_data         (pe_mat_9_18_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_9_18_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_9_18_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_9_19_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_9_19_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_9_19_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_8_19_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_8_19_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_9_19_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_9_19_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_9_20 (
    .io_in_r_data         (pe_mat_9_19_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_9_19_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_9_19_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_9_20_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_9_20_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_9_20_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_8_20_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_8_20_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_9_20_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_9_20_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_9_21 (
    .io_in_r_data         (pe_mat_9_20_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_9_20_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_9_20_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_9_21_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_9_21_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_9_21_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_8_21_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_8_21_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_9_21_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_9_21_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_9_22 (
    .io_in_r_data         (pe_mat_9_21_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_9_21_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_9_21_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_9_22_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_9_22_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_9_22_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_8_22_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_8_22_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_9_22_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_9_22_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_9_23 (
    .io_in_r_data         (pe_mat_9_22_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_9_22_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_9_22_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_9_23_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_9_23_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_9_23_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_8_23_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_8_23_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_9_23_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_9_23_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_9_24 (
    .io_in_r_data         (pe_mat_9_23_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_9_23_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_9_23_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_9_24_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_9_24_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_9_24_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_8_24_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_8_24_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_9_24_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_9_24_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_9_25 (
    .io_in_r_data         (pe_mat_9_24_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_9_24_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_9_24_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_9_25_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_9_25_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_9_25_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_8_25_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_8_25_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_9_25_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_9_25_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_9_26 (
    .io_in_r_data         (pe_mat_9_25_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_9_25_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_9_25_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_9_26_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_9_26_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_9_26_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_8_26_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_8_26_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_9_26_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_9_26_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_9_27 (
    .io_in_r_data         (pe_mat_9_26_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_9_26_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_9_26_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_9_27_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_9_27_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_9_27_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_8_27_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_8_27_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_9_27_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_9_27_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_9_28 (
    .io_in_r_data         (pe_mat_9_27_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_9_27_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_9_27_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_9_28_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_9_28_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_9_28_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_8_28_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_8_28_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_9_28_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_9_28_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_9_29 (
    .io_in_r_data         (pe_mat_9_28_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_9_28_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_9_28_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_9_29_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_9_29_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_9_29_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_8_29_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_8_29_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_9_29_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_9_29_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_9_30 (
    .io_in_r_data         (pe_mat_9_29_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_9_29_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_9_29_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_9_30_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_9_30_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_9_30_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_8_30_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_8_30_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_9_30_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_9_30_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_9_31 (
    .io_in_r_data         (pe_mat_9_30_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_9_30_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_9_30_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_9_31_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_9_31_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_9_31_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_8_31_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_8_31_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_9_31_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_9_31_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_10_0 (
    .io_in_r_data         (io_in_r_10_data[15:0]           ), //i
    .io_in_r_stop_weight  (io_in_r_10_stop_weight          ), //i
    .io_in_r_stall        (io_in_r_10_stall                ), //i
    .io_out_r_data        (pe_mat_10_0_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_10_0_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_10_0_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_9_0_io_out_c_data[15:0]  ), //i
    .io_in_c_is_weight    (pe_mat_9_0_io_out_c_is_weight   ), //i
    .io_out_c_data        (pe_mat_10_0_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_10_0_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_10_1 (
    .io_in_r_data         (pe_mat_10_0_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_10_0_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_10_0_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_10_1_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_10_1_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_10_1_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_9_1_io_out_c_data[15:0]  ), //i
    .io_in_c_is_weight    (pe_mat_9_1_io_out_c_is_weight   ), //i
    .io_out_c_data        (pe_mat_10_1_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_10_1_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_10_2 (
    .io_in_r_data         (pe_mat_10_1_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_10_1_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_10_1_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_10_2_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_10_2_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_10_2_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_9_2_io_out_c_data[15:0]  ), //i
    .io_in_c_is_weight    (pe_mat_9_2_io_out_c_is_weight   ), //i
    .io_out_c_data        (pe_mat_10_2_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_10_2_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_10_3 (
    .io_in_r_data         (pe_mat_10_2_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_10_2_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_10_2_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_10_3_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_10_3_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_10_3_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_9_3_io_out_c_data[15:0]  ), //i
    .io_in_c_is_weight    (pe_mat_9_3_io_out_c_is_weight   ), //i
    .io_out_c_data        (pe_mat_10_3_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_10_3_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_10_4 (
    .io_in_r_data         (pe_mat_10_3_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_10_3_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_10_3_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_10_4_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_10_4_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_10_4_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_9_4_io_out_c_data[15:0]  ), //i
    .io_in_c_is_weight    (pe_mat_9_4_io_out_c_is_weight   ), //i
    .io_out_c_data        (pe_mat_10_4_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_10_4_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_10_5 (
    .io_in_r_data         (pe_mat_10_4_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_10_4_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_10_4_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_10_5_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_10_5_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_10_5_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_9_5_io_out_c_data[15:0]  ), //i
    .io_in_c_is_weight    (pe_mat_9_5_io_out_c_is_weight   ), //i
    .io_out_c_data        (pe_mat_10_5_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_10_5_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_10_6 (
    .io_in_r_data         (pe_mat_10_5_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_10_5_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_10_5_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_10_6_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_10_6_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_10_6_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_9_6_io_out_c_data[15:0]  ), //i
    .io_in_c_is_weight    (pe_mat_9_6_io_out_c_is_weight   ), //i
    .io_out_c_data        (pe_mat_10_6_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_10_6_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_10_7 (
    .io_in_r_data         (pe_mat_10_6_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_10_6_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_10_6_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_10_7_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_10_7_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_10_7_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_9_7_io_out_c_data[15:0]  ), //i
    .io_in_c_is_weight    (pe_mat_9_7_io_out_c_is_weight   ), //i
    .io_out_c_data        (pe_mat_10_7_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_10_7_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_10_8 (
    .io_in_r_data         (pe_mat_10_7_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_10_7_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_10_7_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_10_8_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_10_8_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_10_8_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_9_8_io_out_c_data[15:0]  ), //i
    .io_in_c_is_weight    (pe_mat_9_8_io_out_c_is_weight   ), //i
    .io_out_c_data        (pe_mat_10_8_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_10_8_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_10_9 (
    .io_in_r_data         (pe_mat_10_8_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_10_8_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_10_8_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_10_9_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_10_9_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_10_9_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_9_9_io_out_c_data[15:0]  ), //i
    .io_in_c_is_weight    (pe_mat_9_9_io_out_c_is_weight   ), //i
    .io_out_c_data        (pe_mat_10_9_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_10_9_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_10_10 (
    .io_in_r_data         (pe_mat_10_9_io_out_r_data[15:0]  ), //i
    .io_in_r_stop_weight  (pe_mat_10_9_io_out_r_stop_weight ), //i
    .io_in_r_stall        (pe_mat_10_9_io_out_r_stall       ), //i
    .io_out_r_data        (pe_mat_10_10_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_10_10_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_10_10_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_9_10_io_out_c_data[15:0]  ), //i
    .io_in_c_is_weight    (pe_mat_9_10_io_out_c_is_weight   ), //i
    .io_out_c_data        (pe_mat_10_10_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_10_10_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_10_11 (
    .io_in_r_data         (pe_mat_10_10_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_10_10_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_10_10_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_10_11_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_10_11_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_10_11_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_9_11_io_out_c_data[15:0]  ), //i
    .io_in_c_is_weight    (pe_mat_9_11_io_out_c_is_weight   ), //i
    .io_out_c_data        (pe_mat_10_11_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_10_11_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_10_12 (
    .io_in_r_data         (pe_mat_10_11_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_10_11_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_10_11_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_10_12_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_10_12_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_10_12_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_9_12_io_out_c_data[15:0]  ), //i
    .io_in_c_is_weight    (pe_mat_9_12_io_out_c_is_weight   ), //i
    .io_out_c_data        (pe_mat_10_12_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_10_12_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_10_13 (
    .io_in_r_data         (pe_mat_10_12_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_10_12_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_10_12_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_10_13_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_10_13_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_10_13_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_9_13_io_out_c_data[15:0]  ), //i
    .io_in_c_is_weight    (pe_mat_9_13_io_out_c_is_weight   ), //i
    .io_out_c_data        (pe_mat_10_13_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_10_13_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_10_14 (
    .io_in_r_data         (pe_mat_10_13_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_10_13_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_10_13_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_10_14_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_10_14_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_10_14_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_9_14_io_out_c_data[15:0]  ), //i
    .io_in_c_is_weight    (pe_mat_9_14_io_out_c_is_weight   ), //i
    .io_out_c_data        (pe_mat_10_14_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_10_14_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_10_15 (
    .io_in_r_data         (pe_mat_10_14_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_10_14_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_10_14_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_10_15_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_10_15_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_10_15_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_9_15_io_out_c_data[15:0]  ), //i
    .io_in_c_is_weight    (pe_mat_9_15_io_out_c_is_weight   ), //i
    .io_out_c_data        (pe_mat_10_15_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_10_15_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_10_16 (
    .io_in_r_data         (pe_mat_10_15_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_10_15_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_10_15_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_10_16_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_10_16_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_10_16_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_9_16_io_out_c_data[15:0]  ), //i
    .io_in_c_is_weight    (pe_mat_9_16_io_out_c_is_weight   ), //i
    .io_out_c_data        (pe_mat_10_16_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_10_16_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_10_17 (
    .io_in_r_data         (pe_mat_10_16_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_10_16_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_10_16_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_10_17_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_10_17_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_10_17_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_9_17_io_out_c_data[15:0]  ), //i
    .io_in_c_is_weight    (pe_mat_9_17_io_out_c_is_weight   ), //i
    .io_out_c_data        (pe_mat_10_17_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_10_17_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_10_18 (
    .io_in_r_data         (pe_mat_10_17_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_10_17_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_10_17_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_10_18_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_10_18_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_10_18_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_9_18_io_out_c_data[15:0]  ), //i
    .io_in_c_is_weight    (pe_mat_9_18_io_out_c_is_weight   ), //i
    .io_out_c_data        (pe_mat_10_18_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_10_18_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_10_19 (
    .io_in_r_data         (pe_mat_10_18_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_10_18_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_10_18_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_10_19_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_10_19_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_10_19_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_9_19_io_out_c_data[15:0]  ), //i
    .io_in_c_is_weight    (pe_mat_9_19_io_out_c_is_weight   ), //i
    .io_out_c_data        (pe_mat_10_19_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_10_19_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_10_20 (
    .io_in_r_data         (pe_mat_10_19_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_10_19_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_10_19_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_10_20_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_10_20_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_10_20_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_9_20_io_out_c_data[15:0]  ), //i
    .io_in_c_is_weight    (pe_mat_9_20_io_out_c_is_weight   ), //i
    .io_out_c_data        (pe_mat_10_20_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_10_20_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_10_21 (
    .io_in_r_data         (pe_mat_10_20_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_10_20_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_10_20_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_10_21_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_10_21_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_10_21_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_9_21_io_out_c_data[15:0]  ), //i
    .io_in_c_is_weight    (pe_mat_9_21_io_out_c_is_weight   ), //i
    .io_out_c_data        (pe_mat_10_21_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_10_21_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_10_22 (
    .io_in_r_data         (pe_mat_10_21_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_10_21_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_10_21_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_10_22_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_10_22_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_10_22_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_9_22_io_out_c_data[15:0]  ), //i
    .io_in_c_is_weight    (pe_mat_9_22_io_out_c_is_weight   ), //i
    .io_out_c_data        (pe_mat_10_22_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_10_22_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_10_23 (
    .io_in_r_data         (pe_mat_10_22_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_10_22_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_10_22_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_10_23_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_10_23_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_10_23_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_9_23_io_out_c_data[15:0]  ), //i
    .io_in_c_is_weight    (pe_mat_9_23_io_out_c_is_weight   ), //i
    .io_out_c_data        (pe_mat_10_23_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_10_23_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_10_24 (
    .io_in_r_data         (pe_mat_10_23_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_10_23_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_10_23_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_10_24_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_10_24_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_10_24_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_9_24_io_out_c_data[15:0]  ), //i
    .io_in_c_is_weight    (pe_mat_9_24_io_out_c_is_weight   ), //i
    .io_out_c_data        (pe_mat_10_24_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_10_24_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_10_25 (
    .io_in_r_data         (pe_mat_10_24_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_10_24_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_10_24_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_10_25_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_10_25_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_10_25_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_9_25_io_out_c_data[15:0]  ), //i
    .io_in_c_is_weight    (pe_mat_9_25_io_out_c_is_weight   ), //i
    .io_out_c_data        (pe_mat_10_25_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_10_25_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_10_26 (
    .io_in_r_data         (pe_mat_10_25_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_10_25_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_10_25_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_10_26_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_10_26_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_10_26_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_9_26_io_out_c_data[15:0]  ), //i
    .io_in_c_is_weight    (pe_mat_9_26_io_out_c_is_weight   ), //i
    .io_out_c_data        (pe_mat_10_26_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_10_26_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_10_27 (
    .io_in_r_data         (pe_mat_10_26_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_10_26_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_10_26_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_10_27_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_10_27_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_10_27_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_9_27_io_out_c_data[15:0]  ), //i
    .io_in_c_is_weight    (pe_mat_9_27_io_out_c_is_weight   ), //i
    .io_out_c_data        (pe_mat_10_27_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_10_27_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_10_28 (
    .io_in_r_data         (pe_mat_10_27_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_10_27_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_10_27_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_10_28_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_10_28_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_10_28_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_9_28_io_out_c_data[15:0]  ), //i
    .io_in_c_is_weight    (pe_mat_9_28_io_out_c_is_weight   ), //i
    .io_out_c_data        (pe_mat_10_28_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_10_28_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_10_29 (
    .io_in_r_data         (pe_mat_10_28_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_10_28_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_10_28_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_10_29_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_10_29_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_10_29_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_9_29_io_out_c_data[15:0]  ), //i
    .io_in_c_is_weight    (pe_mat_9_29_io_out_c_is_weight   ), //i
    .io_out_c_data        (pe_mat_10_29_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_10_29_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_10_30 (
    .io_in_r_data         (pe_mat_10_29_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_10_29_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_10_29_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_10_30_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_10_30_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_10_30_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_9_30_io_out_c_data[15:0]  ), //i
    .io_in_c_is_weight    (pe_mat_9_30_io_out_c_is_weight   ), //i
    .io_out_c_data        (pe_mat_10_30_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_10_30_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_10_31 (
    .io_in_r_data         (pe_mat_10_30_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_10_30_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_10_30_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_10_31_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_10_31_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_10_31_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_9_31_io_out_c_data[15:0]  ), //i
    .io_in_c_is_weight    (pe_mat_9_31_io_out_c_is_weight   ), //i
    .io_out_c_data        (pe_mat_10_31_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_10_31_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_11_0 (
    .io_in_r_data         (io_in_r_11_data[15:0]           ), //i
    .io_in_r_stop_weight  (io_in_r_11_stop_weight          ), //i
    .io_in_r_stall        (io_in_r_11_stall                ), //i
    .io_out_r_data        (pe_mat_11_0_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_11_0_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_11_0_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_10_0_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_10_0_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_11_0_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_11_0_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_11_1 (
    .io_in_r_data         (pe_mat_11_0_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_11_0_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_11_0_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_11_1_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_11_1_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_11_1_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_10_1_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_10_1_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_11_1_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_11_1_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_11_2 (
    .io_in_r_data         (pe_mat_11_1_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_11_1_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_11_1_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_11_2_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_11_2_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_11_2_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_10_2_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_10_2_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_11_2_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_11_2_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_11_3 (
    .io_in_r_data         (pe_mat_11_2_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_11_2_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_11_2_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_11_3_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_11_3_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_11_3_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_10_3_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_10_3_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_11_3_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_11_3_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_11_4 (
    .io_in_r_data         (pe_mat_11_3_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_11_3_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_11_3_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_11_4_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_11_4_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_11_4_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_10_4_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_10_4_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_11_4_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_11_4_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_11_5 (
    .io_in_r_data         (pe_mat_11_4_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_11_4_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_11_4_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_11_5_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_11_5_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_11_5_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_10_5_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_10_5_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_11_5_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_11_5_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_11_6 (
    .io_in_r_data         (pe_mat_11_5_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_11_5_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_11_5_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_11_6_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_11_6_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_11_6_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_10_6_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_10_6_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_11_6_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_11_6_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_11_7 (
    .io_in_r_data         (pe_mat_11_6_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_11_6_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_11_6_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_11_7_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_11_7_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_11_7_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_10_7_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_10_7_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_11_7_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_11_7_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_11_8 (
    .io_in_r_data         (pe_mat_11_7_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_11_7_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_11_7_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_11_8_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_11_8_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_11_8_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_10_8_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_10_8_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_11_8_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_11_8_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_11_9 (
    .io_in_r_data         (pe_mat_11_8_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_11_8_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_11_8_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_11_9_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_11_9_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_11_9_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_10_9_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_10_9_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_11_9_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_11_9_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_11_10 (
    .io_in_r_data         (pe_mat_11_9_io_out_r_data[15:0]  ), //i
    .io_in_r_stop_weight  (pe_mat_11_9_io_out_r_stop_weight ), //i
    .io_in_r_stall        (pe_mat_11_9_io_out_r_stall       ), //i
    .io_out_r_data        (pe_mat_11_10_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_11_10_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_11_10_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_10_10_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_10_10_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_11_10_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_11_10_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_11_11 (
    .io_in_r_data         (pe_mat_11_10_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_11_10_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_11_10_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_11_11_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_11_11_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_11_11_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_10_11_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_10_11_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_11_11_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_11_11_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_11_12 (
    .io_in_r_data         (pe_mat_11_11_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_11_11_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_11_11_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_11_12_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_11_12_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_11_12_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_10_12_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_10_12_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_11_12_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_11_12_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_11_13 (
    .io_in_r_data         (pe_mat_11_12_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_11_12_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_11_12_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_11_13_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_11_13_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_11_13_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_10_13_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_10_13_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_11_13_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_11_13_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_11_14 (
    .io_in_r_data         (pe_mat_11_13_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_11_13_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_11_13_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_11_14_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_11_14_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_11_14_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_10_14_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_10_14_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_11_14_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_11_14_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_11_15 (
    .io_in_r_data         (pe_mat_11_14_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_11_14_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_11_14_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_11_15_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_11_15_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_11_15_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_10_15_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_10_15_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_11_15_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_11_15_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_11_16 (
    .io_in_r_data         (pe_mat_11_15_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_11_15_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_11_15_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_11_16_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_11_16_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_11_16_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_10_16_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_10_16_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_11_16_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_11_16_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_11_17 (
    .io_in_r_data         (pe_mat_11_16_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_11_16_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_11_16_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_11_17_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_11_17_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_11_17_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_10_17_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_10_17_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_11_17_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_11_17_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_11_18 (
    .io_in_r_data         (pe_mat_11_17_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_11_17_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_11_17_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_11_18_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_11_18_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_11_18_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_10_18_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_10_18_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_11_18_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_11_18_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_11_19 (
    .io_in_r_data         (pe_mat_11_18_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_11_18_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_11_18_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_11_19_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_11_19_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_11_19_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_10_19_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_10_19_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_11_19_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_11_19_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_11_20 (
    .io_in_r_data         (pe_mat_11_19_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_11_19_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_11_19_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_11_20_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_11_20_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_11_20_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_10_20_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_10_20_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_11_20_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_11_20_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_11_21 (
    .io_in_r_data         (pe_mat_11_20_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_11_20_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_11_20_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_11_21_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_11_21_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_11_21_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_10_21_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_10_21_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_11_21_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_11_21_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_11_22 (
    .io_in_r_data         (pe_mat_11_21_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_11_21_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_11_21_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_11_22_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_11_22_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_11_22_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_10_22_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_10_22_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_11_22_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_11_22_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_11_23 (
    .io_in_r_data         (pe_mat_11_22_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_11_22_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_11_22_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_11_23_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_11_23_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_11_23_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_10_23_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_10_23_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_11_23_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_11_23_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_11_24 (
    .io_in_r_data         (pe_mat_11_23_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_11_23_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_11_23_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_11_24_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_11_24_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_11_24_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_10_24_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_10_24_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_11_24_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_11_24_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_11_25 (
    .io_in_r_data         (pe_mat_11_24_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_11_24_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_11_24_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_11_25_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_11_25_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_11_25_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_10_25_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_10_25_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_11_25_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_11_25_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_11_26 (
    .io_in_r_data         (pe_mat_11_25_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_11_25_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_11_25_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_11_26_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_11_26_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_11_26_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_10_26_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_10_26_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_11_26_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_11_26_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_11_27 (
    .io_in_r_data         (pe_mat_11_26_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_11_26_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_11_26_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_11_27_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_11_27_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_11_27_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_10_27_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_10_27_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_11_27_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_11_27_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_11_28 (
    .io_in_r_data         (pe_mat_11_27_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_11_27_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_11_27_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_11_28_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_11_28_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_11_28_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_10_28_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_10_28_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_11_28_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_11_28_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_11_29 (
    .io_in_r_data         (pe_mat_11_28_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_11_28_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_11_28_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_11_29_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_11_29_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_11_29_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_10_29_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_10_29_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_11_29_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_11_29_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_11_30 (
    .io_in_r_data         (pe_mat_11_29_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_11_29_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_11_29_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_11_30_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_11_30_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_11_30_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_10_30_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_10_30_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_11_30_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_11_30_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_11_31 (
    .io_in_r_data         (pe_mat_11_30_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_11_30_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_11_30_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_11_31_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_11_31_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_11_31_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_10_31_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_10_31_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_11_31_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_11_31_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_12_0 (
    .io_in_r_data         (io_in_r_12_data[15:0]           ), //i
    .io_in_r_stop_weight  (io_in_r_12_stop_weight          ), //i
    .io_in_r_stall        (io_in_r_12_stall                ), //i
    .io_out_r_data        (pe_mat_12_0_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_12_0_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_12_0_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_11_0_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_11_0_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_12_0_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_12_0_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_12_1 (
    .io_in_r_data         (pe_mat_12_0_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_12_0_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_12_0_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_12_1_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_12_1_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_12_1_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_11_1_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_11_1_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_12_1_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_12_1_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_12_2 (
    .io_in_r_data         (pe_mat_12_1_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_12_1_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_12_1_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_12_2_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_12_2_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_12_2_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_11_2_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_11_2_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_12_2_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_12_2_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_12_3 (
    .io_in_r_data         (pe_mat_12_2_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_12_2_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_12_2_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_12_3_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_12_3_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_12_3_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_11_3_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_11_3_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_12_3_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_12_3_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_12_4 (
    .io_in_r_data         (pe_mat_12_3_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_12_3_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_12_3_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_12_4_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_12_4_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_12_4_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_11_4_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_11_4_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_12_4_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_12_4_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_12_5 (
    .io_in_r_data         (pe_mat_12_4_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_12_4_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_12_4_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_12_5_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_12_5_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_12_5_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_11_5_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_11_5_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_12_5_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_12_5_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_12_6 (
    .io_in_r_data         (pe_mat_12_5_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_12_5_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_12_5_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_12_6_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_12_6_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_12_6_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_11_6_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_11_6_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_12_6_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_12_6_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_12_7 (
    .io_in_r_data         (pe_mat_12_6_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_12_6_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_12_6_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_12_7_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_12_7_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_12_7_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_11_7_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_11_7_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_12_7_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_12_7_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_12_8 (
    .io_in_r_data         (pe_mat_12_7_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_12_7_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_12_7_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_12_8_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_12_8_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_12_8_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_11_8_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_11_8_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_12_8_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_12_8_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_12_9 (
    .io_in_r_data         (pe_mat_12_8_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_12_8_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_12_8_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_12_9_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_12_9_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_12_9_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_11_9_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_11_9_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_12_9_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_12_9_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_12_10 (
    .io_in_r_data         (pe_mat_12_9_io_out_r_data[15:0]  ), //i
    .io_in_r_stop_weight  (pe_mat_12_9_io_out_r_stop_weight ), //i
    .io_in_r_stall        (pe_mat_12_9_io_out_r_stall       ), //i
    .io_out_r_data        (pe_mat_12_10_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_12_10_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_12_10_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_11_10_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_11_10_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_12_10_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_12_10_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_12_11 (
    .io_in_r_data         (pe_mat_12_10_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_12_10_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_12_10_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_12_11_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_12_11_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_12_11_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_11_11_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_11_11_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_12_11_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_12_11_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_12_12 (
    .io_in_r_data         (pe_mat_12_11_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_12_11_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_12_11_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_12_12_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_12_12_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_12_12_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_11_12_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_11_12_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_12_12_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_12_12_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_12_13 (
    .io_in_r_data         (pe_mat_12_12_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_12_12_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_12_12_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_12_13_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_12_13_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_12_13_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_11_13_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_11_13_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_12_13_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_12_13_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_12_14 (
    .io_in_r_data         (pe_mat_12_13_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_12_13_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_12_13_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_12_14_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_12_14_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_12_14_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_11_14_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_11_14_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_12_14_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_12_14_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_12_15 (
    .io_in_r_data         (pe_mat_12_14_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_12_14_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_12_14_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_12_15_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_12_15_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_12_15_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_11_15_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_11_15_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_12_15_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_12_15_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_12_16 (
    .io_in_r_data         (pe_mat_12_15_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_12_15_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_12_15_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_12_16_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_12_16_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_12_16_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_11_16_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_11_16_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_12_16_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_12_16_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_12_17 (
    .io_in_r_data         (pe_mat_12_16_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_12_16_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_12_16_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_12_17_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_12_17_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_12_17_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_11_17_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_11_17_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_12_17_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_12_17_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_12_18 (
    .io_in_r_data         (pe_mat_12_17_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_12_17_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_12_17_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_12_18_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_12_18_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_12_18_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_11_18_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_11_18_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_12_18_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_12_18_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_12_19 (
    .io_in_r_data         (pe_mat_12_18_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_12_18_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_12_18_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_12_19_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_12_19_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_12_19_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_11_19_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_11_19_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_12_19_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_12_19_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_12_20 (
    .io_in_r_data         (pe_mat_12_19_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_12_19_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_12_19_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_12_20_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_12_20_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_12_20_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_11_20_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_11_20_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_12_20_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_12_20_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_12_21 (
    .io_in_r_data         (pe_mat_12_20_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_12_20_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_12_20_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_12_21_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_12_21_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_12_21_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_11_21_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_11_21_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_12_21_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_12_21_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_12_22 (
    .io_in_r_data         (pe_mat_12_21_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_12_21_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_12_21_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_12_22_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_12_22_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_12_22_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_11_22_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_11_22_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_12_22_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_12_22_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_12_23 (
    .io_in_r_data         (pe_mat_12_22_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_12_22_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_12_22_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_12_23_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_12_23_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_12_23_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_11_23_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_11_23_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_12_23_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_12_23_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_12_24 (
    .io_in_r_data         (pe_mat_12_23_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_12_23_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_12_23_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_12_24_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_12_24_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_12_24_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_11_24_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_11_24_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_12_24_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_12_24_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_12_25 (
    .io_in_r_data         (pe_mat_12_24_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_12_24_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_12_24_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_12_25_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_12_25_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_12_25_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_11_25_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_11_25_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_12_25_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_12_25_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_12_26 (
    .io_in_r_data         (pe_mat_12_25_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_12_25_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_12_25_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_12_26_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_12_26_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_12_26_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_11_26_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_11_26_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_12_26_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_12_26_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_12_27 (
    .io_in_r_data         (pe_mat_12_26_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_12_26_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_12_26_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_12_27_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_12_27_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_12_27_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_11_27_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_11_27_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_12_27_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_12_27_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_12_28 (
    .io_in_r_data         (pe_mat_12_27_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_12_27_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_12_27_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_12_28_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_12_28_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_12_28_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_11_28_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_11_28_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_12_28_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_12_28_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_12_29 (
    .io_in_r_data         (pe_mat_12_28_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_12_28_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_12_28_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_12_29_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_12_29_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_12_29_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_11_29_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_11_29_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_12_29_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_12_29_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_12_30 (
    .io_in_r_data         (pe_mat_12_29_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_12_29_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_12_29_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_12_30_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_12_30_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_12_30_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_11_30_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_11_30_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_12_30_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_12_30_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_12_31 (
    .io_in_r_data         (pe_mat_12_30_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_12_30_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_12_30_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_12_31_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_12_31_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_12_31_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_11_31_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_11_31_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_12_31_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_12_31_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_13_0 (
    .io_in_r_data         (io_in_r_13_data[15:0]           ), //i
    .io_in_r_stop_weight  (io_in_r_13_stop_weight          ), //i
    .io_in_r_stall        (io_in_r_13_stall                ), //i
    .io_out_r_data        (pe_mat_13_0_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_13_0_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_13_0_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_12_0_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_12_0_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_13_0_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_13_0_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_13_1 (
    .io_in_r_data         (pe_mat_13_0_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_13_0_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_13_0_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_13_1_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_13_1_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_13_1_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_12_1_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_12_1_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_13_1_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_13_1_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_13_2 (
    .io_in_r_data         (pe_mat_13_1_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_13_1_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_13_1_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_13_2_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_13_2_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_13_2_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_12_2_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_12_2_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_13_2_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_13_2_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_13_3 (
    .io_in_r_data         (pe_mat_13_2_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_13_2_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_13_2_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_13_3_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_13_3_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_13_3_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_12_3_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_12_3_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_13_3_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_13_3_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_13_4 (
    .io_in_r_data         (pe_mat_13_3_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_13_3_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_13_3_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_13_4_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_13_4_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_13_4_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_12_4_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_12_4_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_13_4_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_13_4_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_13_5 (
    .io_in_r_data         (pe_mat_13_4_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_13_4_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_13_4_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_13_5_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_13_5_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_13_5_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_12_5_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_12_5_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_13_5_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_13_5_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_13_6 (
    .io_in_r_data         (pe_mat_13_5_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_13_5_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_13_5_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_13_6_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_13_6_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_13_6_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_12_6_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_12_6_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_13_6_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_13_6_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_13_7 (
    .io_in_r_data         (pe_mat_13_6_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_13_6_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_13_6_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_13_7_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_13_7_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_13_7_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_12_7_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_12_7_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_13_7_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_13_7_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_13_8 (
    .io_in_r_data         (pe_mat_13_7_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_13_7_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_13_7_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_13_8_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_13_8_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_13_8_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_12_8_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_12_8_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_13_8_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_13_8_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_13_9 (
    .io_in_r_data         (pe_mat_13_8_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_13_8_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_13_8_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_13_9_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_13_9_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_13_9_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_12_9_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_12_9_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_13_9_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_13_9_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_13_10 (
    .io_in_r_data         (pe_mat_13_9_io_out_r_data[15:0]  ), //i
    .io_in_r_stop_weight  (pe_mat_13_9_io_out_r_stop_weight ), //i
    .io_in_r_stall        (pe_mat_13_9_io_out_r_stall       ), //i
    .io_out_r_data        (pe_mat_13_10_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_13_10_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_13_10_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_12_10_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_12_10_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_13_10_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_13_10_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_13_11 (
    .io_in_r_data         (pe_mat_13_10_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_13_10_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_13_10_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_13_11_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_13_11_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_13_11_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_12_11_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_12_11_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_13_11_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_13_11_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_13_12 (
    .io_in_r_data         (pe_mat_13_11_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_13_11_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_13_11_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_13_12_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_13_12_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_13_12_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_12_12_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_12_12_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_13_12_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_13_12_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_13_13 (
    .io_in_r_data         (pe_mat_13_12_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_13_12_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_13_12_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_13_13_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_13_13_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_13_13_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_12_13_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_12_13_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_13_13_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_13_13_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_13_14 (
    .io_in_r_data         (pe_mat_13_13_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_13_13_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_13_13_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_13_14_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_13_14_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_13_14_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_12_14_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_12_14_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_13_14_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_13_14_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_13_15 (
    .io_in_r_data         (pe_mat_13_14_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_13_14_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_13_14_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_13_15_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_13_15_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_13_15_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_12_15_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_12_15_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_13_15_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_13_15_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_13_16 (
    .io_in_r_data         (pe_mat_13_15_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_13_15_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_13_15_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_13_16_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_13_16_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_13_16_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_12_16_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_12_16_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_13_16_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_13_16_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_13_17 (
    .io_in_r_data         (pe_mat_13_16_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_13_16_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_13_16_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_13_17_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_13_17_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_13_17_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_12_17_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_12_17_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_13_17_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_13_17_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_13_18 (
    .io_in_r_data         (pe_mat_13_17_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_13_17_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_13_17_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_13_18_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_13_18_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_13_18_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_12_18_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_12_18_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_13_18_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_13_18_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_13_19 (
    .io_in_r_data         (pe_mat_13_18_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_13_18_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_13_18_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_13_19_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_13_19_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_13_19_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_12_19_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_12_19_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_13_19_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_13_19_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_13_20 (
    .io_in_r_data         (pe_mat_13_19_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_13_19_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_13_19_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_13_20_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_13_20_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_13_20_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_12_20_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_12_20_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_13_20_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_13_20_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_13_21 (
    .io_in_r_data         (pe_mat_13_20_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_13_20_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_13_20_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_13_21_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_13_21_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_13_21_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_12_21_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_12_21_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_13_21_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_13_21_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_13_22 (
    .io_in_r_data         (pe_mat_13_21_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_13_21_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_13_21_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_13_22_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_13_22_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_13_22_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_12_22_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_12_22_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_13_22_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_13_22_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_13_23 (
    .io_in_r_data         (pe_mat_13_22_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_13_22_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_13_22_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_13_23_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_13_23_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_13_23_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_12_23_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_12_23_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_13_23_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_13_23_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_13_24 (
    .io_in_r_data         (pe_mat_13_23_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_13_23_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_13_23_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_13_24_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_13_24_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_13_24_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_12_24_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_12_24_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_13_24_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_13_24_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_13_25 (
    .io_in_r_data         (pe_mat_13_24_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_13_24_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_13_24_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_13_25_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_13_25_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_13_25_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_12_25_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_12_25_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_13_25_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_13_25_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_13_26 (
    .io_in_r_data         (pe_mat_13_25_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_13_25_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_13_25_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_13_26_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_13_26_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_13_26_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_12_26_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_12_26_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_13_26_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_13_26_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_13_27 (
    .io_in_r_data         (pe_mat_13_26_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_13_26_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_13_26_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_13_27_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_13_27_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_13_27_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_12_27_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_12_27_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_13_27_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_13_27_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_13_28 (
    .io_in_r_data         (pe_mat_13_27_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_13_27_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_13_27_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_13_28_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_13_28_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_13_28_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_12_28_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_12_28_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_13_28_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_13_28_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_13_29 (
    .io_in_r_data         (pe_mat_13_28_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_13_28_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_13_28_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_13_29_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_13_29_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_13_29_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_12_29_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_12_29_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_13_29_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_13_29_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_13_30 (
    .io_in_r_data         (pe_mat_13_29_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_13_29_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_13_29_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_13_30_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_13_30_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_13_30_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_12_30_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_12_30_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_13_30_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_13_30_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_13_31 (
    .io_in_r_data         (pe_mat_13_30_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_13_30_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_13_30_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_13_31_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_13_31_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_13_31_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_12_31_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_12_31_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_13_31_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_13_31_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_14_0 (
    .io_in_r_data         (io_in_r_14_data[15:0]           ), //i
    .io_in_r_stop_weight  (io_in_r_14_stop_weight          ), //i
    .io_in_r_stall        (io_in_r_14_stall                ), //i
    .io_out_r_data        (pe_mat_14_0_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_14_0_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_14_0_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_13_0_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_13_0_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_14_0_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_14_0_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_14_1 (
    .io_in_r_data         (pe_mat_14_0_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_14_0_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_14_0_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_14_1_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_14_1_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_14_1_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_13_1_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_13_1_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_14_1_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_14_1_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_14_2 (
    .io_in_r_data         (pe_mat_14_1_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_14_1_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_14_1_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_14_2_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_14_2_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_14_2_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_13_2_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_13_2_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_14_2_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_14_2_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_14_3 (
    .io_in_r_data         (pe_mat_14_2_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_14_2_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_14_2_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_14_3_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_14_3_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_14_3_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_13_3_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_13_3_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_14_3_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_14_3_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_14_4 (
    .io_in_r_data         (pe_mat_14_3_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_14_3_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_14_3_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_14_4_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_14_4_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_14_4_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_13_4_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_13_4_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_14_4_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_14_4_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_14_5 (
    .io_in_r_data         (pe_mat_14_4_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_14_4_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_14_4_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_14_5_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_14_5_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_14_5_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_13_5_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_13_5_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_14_5_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_14_5_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_14_6 (
    .io_in_r_data         (pe_mat_14_5_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_14_5_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_14_5_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_14_6_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_14_6_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_14_6_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_13_6_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_13_6_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_14_6_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_14_6_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_14_7 (
    .io_in_r_data         (pe_mat_14_6_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_14_6_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_14_6_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_14_7_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_14_7_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_14_7_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_13_7_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_13_7_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_14_7_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_14_7_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_14_8 (
    .io_in_r_data         (pe_mat_14_7_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_14_7_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_14_7_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_14_8_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_14_8_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_14_8_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_13_8_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_13_8_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_14_8_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_14_8_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_14_9 (
    .io_in_r_data         (pe_mat_14_8_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_14_8_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_14_8_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_14_9_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_14_9_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_14_9_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_13_9_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_13_9_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_14_9_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_14_9_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_14_10 (
    .io_in_r_data         (pe_mat_14_9_io_out_r_data[15:0]  ), //i
    .io_in_r_stop_weight  (pe_mat_14_9_io_out_r_stop_weight ), //i
    .io_in_r_stall        (pe_mat_14_9_io_out_r_stall       ), //i
    .io_out_r_data        (pe_mat_14_10_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_14_10_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_14_10_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_13_10_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_13_10_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_14_10_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_14_10_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_14_11 (
    .io_in_r_data         (pe_mat_14_10_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_14_10_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_14_10_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_14_11_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_14_11_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_14_11_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_13_11_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_13_11_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_14_11_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_14_11_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_14_12 (
    .io_in_r_data         (pe_mat_14_11_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_14_11_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_14_11_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_14_12_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_14_12_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_14_12_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_13_12_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_13_12_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_14_12_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_14_12_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_14_13 (
    .io_in_r_data         (pe_mat_14_12_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_14_12_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_14_12_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_14_13_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_14_13_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_14_13_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_13_13_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_13_13_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_14_13_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_14_13_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_14_14 (
    .io_in_r_data         (pe_mat_14_13_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_14_13_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_14_13_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_14_14_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_14_14_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_14_14_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_13_14_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_13_14_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_14_14_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_14_14_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_14_15 (
    .io_in_r_data         (pe_mat_14_14_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_14_14_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_14_14_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_14_15_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_14_15_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_14_15_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_13_15_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_13_15_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_14_15_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_14_15_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_14_16 (
    .io_in_r_data         (pe_mat_14_15_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_14_15_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_14_15_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_14_16_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_14_16_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_14_16_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_13_16_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_13_16_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_14_16_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_14_16_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_14_17 (
    .io_in_r_data         (pe_mat_14_16_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_14_16_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_14_16_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_14_17_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_14_17_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_14_17_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_13_17_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_13_17_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_14_17_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_14_17_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_14_18 (
    .io_in_r_data         (pe_mat_14_17_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_14_17_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_14_17_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_14_18_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_14_18_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_14_18_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_13_18_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_13_18_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_14_18_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_14_18_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_14_19 (
    .io_in_r_data         (pe_mat_14_18_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_14_18_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_14_18_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_14_19_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_14_19_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_14_19_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_13_19_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_13_19_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_14_19_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_14_19_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_14_20 (
    .io_in_r_data         (pe_mat_14_19_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_14_19_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_14_19_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_14_20_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_14_20_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_14_20_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_13_20_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_13_20_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_14_20_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_14_20_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_14_21 (
    .io_in_r_data         (pe_mat_14_20_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_14_20_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_14_20_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_14_21_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_14_21_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_14_21_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_13_21_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_13_21_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_14_21_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_14_21_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_14_22 (
    .io_in_r_data         (pe_mat_14_21_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_14_21_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_14_21_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_14_22_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_14_22_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_14_22_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_13_22_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_13_22_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_14_22_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_14_22_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_14_23 (
    .io_in_r_data         (pe_mat_14_22_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_14_22_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_14_22_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_14_23_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_14_23_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_14_23_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_13_23_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_13_23_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_14_23_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_14_23_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_14_24 (
    .io_in_r_data         (pe_mat_14_23_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_14_23_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_14_23_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_14_24_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_14_24_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_14_24_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_13_24_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_13_24_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_14_24_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_14_24_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_14_25 (
    .io_in_r_data         (pe_mat_14_24_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_14_24_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_14_24_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_14_25_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_14_25_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_14_25_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_13_25_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_13_25_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_14_25_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_14_25_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_14_26 (
    .io_in_r_data         (pe_mat_14_25_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_14_25_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_14_25_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_14_26_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_14_26_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_14_26_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_13_26_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_13_26_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_14_26_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_14_26_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_14_27 (
    .io_in_r_data         (pe_mat_14_26_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_14_26_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_14_26_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_14_27_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_14_27_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_14_27_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_13_27_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_13_27_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_14_27_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_14_27_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_14_28 (
    .io_in_r_data         (pe_mat_14_27_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_14_27_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_14_27_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_14_28_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_14_28_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_14_28_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_13_28_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_13_28_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_14_28_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_14_28_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_14_29 (
    .io_in_r_data         (pe_mat_14_28_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_14_28_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_14_28_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_14_29_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_14_29_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_14_29_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_13_29_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_13_29_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_14_29_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_14_29_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_14_30 (
    .io_in_r_data         (pe_mat_14_29_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_14_29_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_14_29_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_14_30_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_14_30_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_14_30_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_13_30_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_13_30_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_14_30_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_14_30_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_14_31 (
    .io_in_r_data         (pe_mat_14_30_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_14_30_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_14_30_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_14_31_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_14_31_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_14_31_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_13_31_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_13_31_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_14_31_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_14_31_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_15_0 (
    .io_in_r_data         (io_in_r_15_data[15:0]           ), //i
    .io_in_r_stop_weight  (io_in_r_15_stop_weight          ), //i
    .io_in_r_stall        (io_in_r_15_stall                ), //i
    .io_out_r_data        (pe_mat_15_0_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_15_0_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_15_0_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_14_0_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_14_0_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_15_0_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_15_0_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_15_1 (
    .io_in_r_data         (pe_mat_15_0_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_15_0_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_15_0_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_15_1_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_15_1_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_15_1_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_14_1_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_14_1_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_15_1_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_15_1_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_15_2 (
    .io_in_r_data         (pe_mat_15_1_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_15_1_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_15_1_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_15_2_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_15_2_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_15_2_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_14_2_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_14_2_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_15_2_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_15_2_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_15_3 (
    .io_in_r_data         (pe_mat_15_2_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_15_2_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_15_2_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_15_3_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_15_3_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_15_3_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_14_3_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_14_3_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_15_3_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_15_3_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_15_4 (
    .io_in_r_data         (pe_mat_15_3_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_15_3_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_15_3_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_15_4_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_15_4_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_15_4_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_14_4_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_14_4_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_15_4_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_15_4_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_15_5 (
    .io_in_r_data         (pe_mat_15_4_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_15_4_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_15_4_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_15_5_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_15_5_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_15_5_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_14_5_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_14_5_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_15_5_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_15_5_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_15_6 (
    .io_in_r_data         (pe_mat_15_5_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_15_5_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_15_5_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_15_6_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_15_6_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_15_6_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_14_6_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_14_6_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_15_6_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_15_6_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_15_7 (
    .io_in_r_data         (pe_mat_15_6_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_15_6_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_15_6_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_15_7_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_15_7_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_15_7_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_14_7_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_14_7_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_15_7_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_15_7_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_15_8 (
    .io_in_r_data         (pe_mat_15_7_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_15_7_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_15_7_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_15_8_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_15_8_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_15_8_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_14_8_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_14_8_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_15_8_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_15_8_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_15_9 (
    .io_in_r_data         (pe_mat_15_8_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_15_8_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_15_8_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_15_9_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_15_9_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_15_9_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_14_9_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_14_9_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_15_9_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_15_9_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_15_10 (
    .io_in_r_data         (pe_mat_15_9_io_out_r_data[15:0]  ), //i
    .io_in_r_stop_weight  (pe_mat_15_9_io_out_r_stop_weight ), //i
    .io_in_r_stall        (pe_mat_15_9_io_out_r_stall       ), //i
    .io_out_r_data        (pe_mat_15_10_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_15_10_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_15_10_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_14_10_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_14_10_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_15_10_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_15_10_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_15_11 (
    .io_in_r_data         (pe_mat_15_10_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_15_10_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_15_10_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_15_11_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_15_11_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_15_11_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_14_11_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_14_11_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_15_11_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_15_11_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_15_12 (
    .io_in_r_data         (pe_mat_15_11_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_15_11_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_15_11_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_15_12_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_15_12_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_15_12_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_14_12_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_14_12_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_15_12_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_15_12_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_15_13 (
    .io_in_r_data         (pe_mat_15_12_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_15_12_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_15_12_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_15_13_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_15_13_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_15_13_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_14_13_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_14_13_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_15_13_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_15_13_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_15_14 (
    .io_in_r_data         (pe_mat_15_13_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_15_13_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_15_13_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_15_14_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_15_14_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_15_14_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_14_14_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_14_14_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_15_14_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_15_14_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_15_15 (
    .io_in_r_data         (pe_mat_15_14_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_15_14_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_15_14_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_15_15_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_15_15_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_15_15_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_14_15_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_14_15_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_15_15_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_15_15_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_15_16 (
    .io_in_r_data         (pe_mat_15_15_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_15_15_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_15_15_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_15_16_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_15_16_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_15_16_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_14_16_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_14_16_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_15_16_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_15_16_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_15_17 (
    .io_in_r_data         (pe_mat_15_16_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_15_16_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_15_16_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_15_17_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_15_17_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_15_17_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_14_17_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_14_17_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_15_17_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_15_17_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_15_18 (
    .io_in_r_data         (pe_mat_15_17_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_15_17_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_15_17_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_15_18_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_15_18_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_15_18_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_14_18_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_14_18_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_15_18_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_15_18_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_15_19 (
    .io_in_r_data         (pe_mat_15_18_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_15_18_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_15_18_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_15_19_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_15_19_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_15_19_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_14_19_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_14_19_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_15_19_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_15_19_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_15_20 (
    .io_in_r_data         (pe_mat_15_19_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_15_19_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_15_19_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_15_20_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_15_20_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_15_20_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_14_20_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_14_20_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_15_20_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_15_20_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_15_21 (
    .io_in_r_data         (pe_mat_15_20_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_15_20_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_15_20_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_15_21_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_15_21_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_15_21_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_14_21_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_14_21_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_15_21_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_15_21_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_15_22 (
    .io_in_r_data         (pe_mat_15_21_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_15_21_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_15_21_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_15_22_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_15_22_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_15_22_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_14_22_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_14_22_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_15_22_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_15_22_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_15_23 (
    .io_in_r_data         (pe_mat_15_22_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_15_22_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_15_22_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_15_23_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_15_23_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_15_23_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_14_23_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_14_23_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_15_23_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_15_23_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_15_24 (
    .io_in_r_data         (pe_mat_15_23_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_15_23_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_15_23_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_15_24_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_15_24_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_15_24_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_14_24_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_14_24_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_15_24_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_15_24_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_15_25 (
    .io_in_r_data         (pe_mat_15_24_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_15_24_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_15_24_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_15_25_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_15_25_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_15_25_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_14_25_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_14_25_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_15_25_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_15_25_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_15_26 (
    .io_in_r_data         (pe_mat_15_25_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_15_25_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_15_25_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_15_26_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_15_26_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_15_26_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_14_26_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_14_26_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_15_26_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_15_26_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_15_27 (
    .io_in_r_data         (pe_mat_15_26_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_15_26_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_15_26_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_15_27_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_15_27_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_15_27_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_14_27_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_14_27_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_15_27_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_15_27_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_15_28 (
    .io_in_r_data         (pe_mat_15_27_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_15_27_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_15_27_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_15_28_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_15_28_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_15_28_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_14_28_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_14_28_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_15_28_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_15_28_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_15_29 (
    .io_in_r_data         (pe_mat_15_28_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_15_28_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_15_28_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_15_29_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_15_29_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_15_29_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_14_29_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_14_29_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_15_29_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_15_29_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_15_30 (
    .io_in_r_data         (pe_mat_15_29_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_15_29_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_15_29_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_15_30_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_15_30_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_15_30_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_14_30_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_14_30_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_15_30_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_15_30_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_15_31 (
    .io_in_r_data         (pe_mat_15_30_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_15_30_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_15_30_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_15_31_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_15_31_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_15_31_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_14_31_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_14_31_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_15_31_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_15_31_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_16_0 (
    .io_in_r_data         (io_in_r_16_data[15:0]           ), //i
    .io_in_r_stop_weight  (io_in_r_16_stop_weight          ), //i
    .io_in_r_stall        (io_in_r_16_stall                ), //i
    .io_out_r_data        (pe_mat_16_0_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_16_0_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_16_0_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_15_0_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_15_0_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_16_0_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_16_0_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_16_1 (
    .io_in_r_data         (pe_mat_16_0_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_16_0_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_16_0_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_16_1_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_16_1_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_16_1_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_15_1_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_15_1_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_16_1_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_16_1_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_16_2 (
    .io_in_r_data         (pe_mat_16_1_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_16_1_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_16_1_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_16_2_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_16_2_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_16_2_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_15_2_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_15_2_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_16_2_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_16_2_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_16_3 (
    .io_in_r_data         (pe_mat_16_2_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_16_2_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_16_2_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_16_3_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_16_3_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_16_3_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_15_3_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_15_3_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_16_3_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_16_3_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_16_4 (
    .io_in_r_data         (pe_mat_16_3_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_16_3_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_16_3_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_16_4_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_16_4_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_16_4_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_15_4_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_15_4_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_16_4_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_16_4_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_16_5 (
    .io_in_r_data         (pe_mat_16_4_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_16_4_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_16_4_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_16_5_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_16_5_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_16_5_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_15_5_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_15_5_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_16_5_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_16_5_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_16_6 (
    .io_in_r_data         (pe_mat_16_5_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_16_5_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_16_5_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_16_6_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_16_6_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_16_6_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_15_6_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_15_6_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_16_6_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_16_6_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_16_7 (
    .io_in_r_data         (pe_mat_16_6_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_16_6_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_16_6_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_16_7_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_16_7_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_16_7_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_15_7_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_15_7_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_16_7_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_16_7_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_16_8 (
    .io_in_r_data         (pe_mat_16_7_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_16_7_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_16_7_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_16_8_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_16_8_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_16_8_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_15_8_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_15_8_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_16_8_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_16_8_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_16_9 (
    .io_in_r_data         (pe_mat_16_8_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_16_8_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_16_8_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_16_9_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_16_9_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_16_9_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_15_9_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_15_9_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_16_9_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_16_9_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_16_10 (
    .io_in_r_data         (pe_mat_16_9_io_out_r_data[15:0]  ), //i
    .io_in_r_stop_weight  (pe_mat_16_9_io_out_r_stop_weight ), //i
    .io_in_r_stall        (pe_mat_16_9_io_out_r_stall       ), //i
    .io_out_r_data        (pe_mat_16_10_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_16_10_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_16_10_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_15_10_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_15_10_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_16_10_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_16_10_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_16_11 (
    .io_in_r_data         (pe_mat_16_10_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_16_10_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_16_10_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_16_11_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_16_11_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_16_11_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_15_11_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_15_11_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_16_11_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_16_11_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_16_12 (
    .io_in_r_data         (pe_mat_16_11_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_16_11_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_16_11_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_16_12_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_16_12_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_16_12_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_15_12_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_15_12_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_16_12_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_16_12_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_16_13 (
    .io_in_r_data         (pe_mat_16_12_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_16_12_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_16_12_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_16_13_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_16_13_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_16_13_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_15_13_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_15_13_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_16_13_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_16_13_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_16_14 (
    .io_in_r_data         (pe_mat_16_13_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_16_13_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_16_13_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_16_14_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_16_14_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_16_14_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_15_14_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_15_14_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_16_14_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_16_14_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_16_15 (
    .io_in_r_data         (pe_mat_16_14_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_16_14_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_16_14_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_16_15_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_16_15_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_16_15_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_15_15_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_15_15_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_16_15_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_16_15_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_16_16 (
    .io_in_r_data         (pe_mat_16_15_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_16_15_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_16_15_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_16_16_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_16_16_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_16_16_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_15_16_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_15_16_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_16_16_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_16_16_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_16_17 (
    .io_in_r_data         (pe_mat_16_16_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_16_16_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_16_16_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_16_17_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_16_17_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_16_17_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_15_17_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_15_17_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_16_17_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_16_17_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_16_18 (
    .io_in_r_data         (pe_mat_16_17_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_16_17_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_16_17_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_16_18_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_16_18_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_16_18_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_15_18_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_15_18_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_16_18_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_16_18_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_16_19 (
    .io_in_r_data         (pe_mat_16_18_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_16_18_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_16_18_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_16_19_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_16_19_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_16_19_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_15_19_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_15_19_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_16_19_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_16_19_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_16_20 (
    .io_in_r_data         (pe_mat_16_19_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_16_19_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_16_19_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_16_20_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_16_20_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_16_20_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_15_20_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_15_20_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_16_20_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_16_20_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_16_21 (
    .io_in_r_data         (pe_mat_16_20_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_16_20_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_16_20_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_16_21_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_16_21_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_16_21_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_15_21_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_15_21_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_16_21_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_16_21_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_16_22 (
    .io_in_r_data         (pe_mat_16_21_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_16_21_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_16_21_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_16_22_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_16_22_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_16_22_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_15_22_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_15_22_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_16_22_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_16_22_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_16_23 (
    .io_in_r_data         (pe_mat_16_22_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_16_22_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_16_22_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_16_23_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_16_23_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_16_23_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_15_23_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_15_23_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_16_23_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_16_23_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_16_24 (
    .io_in_r_data         (pe_mat_16_23_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_16_23_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_16_23_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_16_24_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_16_24_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_16_24_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_15_24_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_15_24_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_16_24_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_16_24_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_16_25 (
    .io_in_r_data         (pe_mat_16_24_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_16_24_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_16_24_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_16_25_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_16_25_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_16_25_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_15_25_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_15_25_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_16_25_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_16_25_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_16_26 (
    .io_in_r_data         (pe_mat_16_25_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_16_25_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_16_25_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_16_26_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_16_26_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_16_26_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_15_26_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_15_26_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_16_26_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_16_26_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_16_27 (
    .io_in_r_data         (pe_mat_16_26_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_16_26_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_16_26_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_16_27_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_16_27_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_16_27_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_15_27_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_15_27_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_16_27_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_16_27_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_16_28 (
    .io_in_r_data         (pe_mat_16_27_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_16_27_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_16_27_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_16_28_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_16_28_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_16_28_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_15_28_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_15_28_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_16_28_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_16_28_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_16_29 (
    .io_in_r_data         (pe_mat_16_28_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_16_28_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_16_28_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_16_29_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_16_29_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_16_29_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_15_29_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_15_29_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_16_29_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_16_29_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_16_30 (
    .io_in_r_data         (pe_mat_16_29_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_16_29_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_16_29_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_16_30_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_16_30_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_16_30_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_15_30_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_15_30_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_16_30_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_16_30_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_16_31 (
    .io_in_r_data         (pe_mat_16_30_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_16_30_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_16_30_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_16_31_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_16_31_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_16_31_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_15_31_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_15_31_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_16_31_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_16_31_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_17_0 (
    .io_in_r_data         (io_in_r_17_data[15:0]           ), //i
    .io_in_r_stop_weight  (io_in_r_17_stop_weight          ), //i
    .io_in_r_stall        (io_in_r_17_stall                ), //i
    .io_out_r_data        (pe_mat_17_0_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_17_0_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_17_0_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_16_0_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_16_0_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_17_0_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_17_0_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_17_1 (
    .io_in_r_data         (pe_mat_17_0_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_17_0_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_17_0_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_17_1_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_17_1_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_17_1_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_16_1_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_16_1_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_17_1_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_17_1_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_17_2 (
    .io_in_r_data         (pe_mat_17_1_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_17_1_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_17_1_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_17_2_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_17_2_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_17_2_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_16_2_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_16_2_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_17_2_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_17_2_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_17_3 (
    .io_in_r_data         (pe_mat_17_2_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_17_2_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_17_2_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_17_3_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_17_3_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_17_3_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_16_3_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_16_3_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_17_3_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_17_3_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_17_4 (
    .io_in_r_data         (pe_mat_17_3_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_17_3_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_17_3_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_17_4_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_17_4_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_17_4_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_16_4_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_16_4_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_17_4_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_17_4_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_17_5 (
    .io_in_r_data         (pe_mat_17_4_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_17_4_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_17_4_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_17_5_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_17_5_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_17_5_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_16_5_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_16_5_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_17_5_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_17_5_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_17_6 (
    .io_in_r_data         (pe_mat_17_5_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_17_5_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_17_5_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_17_6_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_17_6_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_17_6_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_16_6_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_16_6_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_17_6_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_17_6_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_17_7 (
    .io_in_r_data         (pe_mat_17_6_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_17_6_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_17_6_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_17_7_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_17_7_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_17_7_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_16_7_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_16_7_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_17_7_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_17_7_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_17_8 (
    .io_in_r_data         (pe_mat_17_7_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_17_7_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_17_7_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_17_8_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_17_8_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_17_8_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_16_8_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_16_8_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_17_8_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_17_8_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_17_9 (
    .io_in_r_data         (pe_mat_17_8_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_17_8_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_17_8_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_17_9_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_17_9_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_17_9_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_16_9_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_16_9_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_17_9_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_17_9_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_17_10 (
    .io_in_r_data         (pe_mat_17_9_io_out_r_data[15:0]  ), //i
    .io_in_r_stop_weight  (pe_mat_17_9_io_out_r_stop_weight ), //i
    .io_in_r_stall        (pe_mat_17_9_io_out_r_stall       ), //i
    .io_out_r_data        (pe_mat_17_10_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_17_10_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_17_10_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_16_10_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_16_10_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_17_10_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_17_10_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_17_11 (
    .io_in_r_data         (pe_mat_17_10_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_17_10_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_17_10_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_17_11_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_17_11_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_17_11_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_16_11_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_16_11_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_17_11_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_17_11_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_17_12 (
    .io_in_r_data         (pe_mat_17_11_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_17_11_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_17_11_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_17_12_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_17_12_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_17_12_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_16_12_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_16_12_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_17_12_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_17_12_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_17_13 (
    .io_in_r_data         (pe_mat_17_12_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_17_12_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_17_12_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_17_13_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_17_13_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_17_13_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_16_13_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_16_13_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_17_13_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_17_13_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_17_14 (
    .io_in_r_data         (pe_mat_17_13_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_17_13_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_17_13_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_17_14_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_17_14_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_17_14_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_16_14_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_16_14_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_17_14_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_17_14_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_17_15 (
    .io_in_r_data         (pe_mat_17_14_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_17_14_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_17_14_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_17_15_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_17_15_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_17_15_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_16_15_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_16_15_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_17_15_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_17_15_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_17_16 (
    .io_in_r_data         (pe_mat_17_15_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_17_15_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_17_15_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_17_16_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_17_16_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_17_16_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_16_16_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_16_16_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_17_16_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_17_16_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_17_17 (
    .io_in_r_data         (pe_mat_17_16_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_17_16_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_17_16_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_17_17_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_17_17_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_17_17_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_16_17_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_16_17_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_17_17_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_17_17_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_17_18 (
    .io_in_r_data         (pe_mat_17_17_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_17_17_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_17_17_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_17_18_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_17_18_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_17_18_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_16_18_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_16_18_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_17_18_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_17_18_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_17_19 (
    .io_in_r_data         (pe_mat_17_18_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_17_18_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_17_18_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_17_19_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_17_19_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_17_19_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_16_19_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_16_19_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_17_19_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_17_19_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_17_20 (
    .io_in_r_data         (pe_mat_17_19_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_17_19_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_17_19_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_17_20_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_17_20_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_17_20_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_16_20_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_16_20_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_17_20_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_17_20_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_17_21 (
    .io_in_r_data         (pe_mat_17_20_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_17_20_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_17_20_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_17_21_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_17_21_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_17_21_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_16_21_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_16_21_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_17_21_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_17_21_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_17_22 (
    .io_in_r_data         (pe_mat_17_21_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_17_21_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_17_21_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_17_22_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_17_22_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_17_22_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_16_22_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_16_22_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_17_22_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_17_22_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_17_23 (
    .io_in_r_data         (pe_mat_17_22_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_17_22_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_17_22_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_17_23_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_17_23_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_17_23_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_16_23_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_16_23_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_17_23_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_17_23_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_17_24 (
    .io_in_r_data         (pe_mat_17_23_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_17_23_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_17_23_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_17_24_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_17_24_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_17_24_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_16_24_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_16_24_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_17_24_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_17_24_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_17_25 (
    .io_in_r_data         (pe_mat_17_24_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_17_24_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_17_24_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_17_25_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_17_25_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_17_25_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_16_25_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_16_25_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_17_25_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_17_25_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_17_26 (
    .io_in_r_data         (pe_mat_17_25_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_17_25_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_17_25_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_17_26_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_17_26_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_17_26_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_16_26_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_16_26_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_17_26_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_17_26_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_17_27 (
    .io_in_r_data         (pe_mat_17_26_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_17_26_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_17_26_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_17_27_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_17_27_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_17_27_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_16_27_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_16_27_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_17_27_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_17_27_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_17_28 (
    .io_in_r_data         (pe_mat_17_27_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_17_27_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_17_27_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_17_28_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_17_28_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_17_28_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_16_28_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_16_28_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_17_28_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_17_28_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_17_29 (
    .io_in_r_data         (pe_mat_17_28_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_17_28_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_17_28_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_17_29_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_17_29_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_17_29_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_16_29_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_16_29_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_17_29_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_17_29_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_17_30 (
    .io_in_r_data         (pe_mat_17_29_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_17_29_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_17_29_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_17_30_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_17_30_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_17_30_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_16_30_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_16_30_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_17_30_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_17_30_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_17_31 (
    .io_in_r_data         (pe_mat_17_30_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_17_30_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_17_30_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_17_31_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_17_31_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_17_31_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_16_31_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_16_31_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_17_31_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_17_31_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_18_0 (
    .io_in_r_data         (io_in_r_18_data[15:0]           ), //i
    .io_in_r_stop_weight  (io_in_r_18_stop_weight          ), //i
    .io_in_r_stall        (io_in_r_18_stall                ), //i
    .io_out_r_data        (pe_mat_18_0_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_18_0_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_18_0_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_17_0_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_17_0_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_18_0_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_18_0_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_18_1 (
    .io_in_r_data         (pe_mat_18_0_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_18_0_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_18_0_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_18_1_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_18_1_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_18_1_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_17_1_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_17_1_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_18_1_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_18_1_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_18_2 (
    .io_in_r_data         (pe_mat_18_1_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_18_1_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_18_1_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_18_2_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_18_2_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_18_2_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_17_2_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_17_2_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_18_2_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_18_2_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_18_3 (
    .io_in_r_data         (pe_mat_18_2_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_18_2_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_18_2_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_18_3_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_18_3_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_18_3_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_17_3_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_17_3_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_18_3_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_18_3_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_18_4 (
    .io_in_r_data         (pe_mat_18_3_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_18_3_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_18_3_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_18_4_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_18_4_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_18_4_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_17_4_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_17_4_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_18_4_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_18_4_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_18_5 (
    .io_in_r_data         (pe_mat_18_4_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_18_4_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_18_4_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_18_5_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_18_5_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_18_5_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_17_5_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_17_5_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_18_5_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_18_5_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_18_6 (
    .io_in_r_data         (pe_mat_18_5_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_18_5_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_18_5_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_18_6_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_18_6_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_18_6_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_17_6_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_17_6_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_18_6_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_18_6_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_18_7 (
    .io_in_r_data         (pe_mat_18_6_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_18_6_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_18_6_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_18_7_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_18_7_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_18_7_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_17_7_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_17_7_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_18_7_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_18_7_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_18_8 (
    .io_in_r_data         (pe_mat_18_7_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_18_7_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_18_7_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_18_8_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_18_8_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_18_8_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_17_8_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_17_8_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_18_8_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_18_8_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_18_9 (
    .io_in_r_data         (pe_mat_18_8_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_18_8_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_18_8_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_18_9_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_18_9_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_18_9_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_17_9_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_17_9_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_18_9_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_18_9_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_18_10 (
    .io_in_r_data         (pe_mat_18_9_io_out_r_data[15:0]  ), //i
    .io_in_r_stop_weight  (pe_mat_18_9_io_out_r_stop_weight ), //i
    .io_in_r_stall        (pe_mat_18_9_io_out_r_stall       ), //i
    .io_out_r_data        (pe_mat_18_10_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_18_10_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_18_10_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_17_10_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_17_10_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_18_10_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_18_10_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_18_11 (
    .io_in_r_data         (pe_mat_18_10_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_18_10_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_18_10_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_18_11_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_18_11_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_18_11_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_17_11_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_17_11_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_18_11_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_18_11_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_18_12 (
    .io_in_r_data         (pe_mat_18_11_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_18_11_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_18_11_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_18_12_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_18_12_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_18_12_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_17_12_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_17_12_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_18_12_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_18_12_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_18_13 (
    .io_in_r_data         (pe_mat_18_12_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_18_12_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_18_12_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_18_13_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_18_13_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_18_13_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_17_13_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_17_13_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_18_13_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_18_13_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_18_14 (
    .io_in_r_data         (pe_mat_18_13_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_18_13_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_18_13_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_18_14_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_18_14_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_18_14_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_17_14_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_17_14_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_18_14_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_18_14_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_18_15 (
    .io_in_r_data         (pe_mat_18_14_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_18_14_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_18_14_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_18_15_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_18_15_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_18_15_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_17_15_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_17_15_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_18_15_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_18_15_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_18_16 (
    .io_in_r_data         (pe_mat_18_15_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_18_15_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_18_15_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_18_16_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_18_16_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_18_16_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_17_16_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_17_16_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_18_16_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_18_16_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_18_17 (
    .io_in_r_data         (pe_mat_18_16_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_18_16_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_18_16_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_18_17_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_18_17_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_18_17_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_17_17_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_17_17_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_18_17_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_18_17_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_18_18 (
    .io_in_r_data         (pe_mat_18_17_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_18_17_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_18_17_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_18_18_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_18_18_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_18_18_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_17_18_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_17_18_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_18_18_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_18_18_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_18_19 (
    .io_in_r_data         (pe_mat_18_18_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_18_18_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_18_18_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_18_19_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_18_19_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_18_19_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_17_19_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_17_19_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_18_19_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_18_19_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_18_20 (
    .io_in_r_data         (pe_mat_18_19_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_18_19_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_18_19_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_18_20_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_18_20_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_18_20_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_17_20_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_17_20_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_18_20_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_18_20_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_18_21 (
    .io_in_r_data         (pe_mat_18_20_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_18_20_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_18_20_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_18_21_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_18_21_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_18_21_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_17_21_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_17_21_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_18_21_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_18_21_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_18_22 (
    .io_in_r_data         (pe_mat_18_21_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_18_21_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_18_21_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_18_22_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_18_22_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_18_22_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_17_22_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_17_22_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_18_22_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_18_22_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_18_23 (
    .io_in_r_data         (pe_mat_18_22_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_18_22_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_18_22_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_18_23_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_18_23_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_18_23_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_17_23_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_17_23_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_18_23_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_18_23_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_18_24 (
    .io_in_r_data         (pe_mat_18_23_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_18_23_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_18_23_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_18_24_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_18_24_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_18_24_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_17_24_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_17_24_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_18_24_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_18_24_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_18_25 (
    .io_in_r_data         (pe_mat_18_24_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_18_24_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_18_24_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_18_25_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_18_25_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_18_25_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_17_25_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_17_25_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_18_25_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_18_25_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_18_26 (
    .io_in_r_data         (pe_mat_18_25_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_18_25_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_18_25_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_18_26_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_18_26_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_18_26_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_17_26_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_17_26_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_18_26_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_18_26_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_18_27 (
    .io_in_r_data         (pe_mat_18_26_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_18_26_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_18_26_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_18_27_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_18_27_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_18_27_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_17_27_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_17_27_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_18_27_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_18_27_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_18_28 (
    .io_in_r_data         (pe_mat_18_27_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_18_27_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_18_27_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_18_28_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_18_28_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_18_28_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_17_28_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_17_28_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_18_28_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_18_28_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_18_29 (
    .io_in_r_data         (pe_mat_18_28_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_18_28_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_18_28_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_18_29_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_18_29_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_18_29_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_17_29_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_17_29_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_18_29_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_18_29_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_18_30 (
    .io_in_r_data         (pe_mat_18_29_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_18_29_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_18_29_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_18_30_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_18_30_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_18_30_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_17_30_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_17_30_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_18_30_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_18_30_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_18_31 (
    .io_in_r_data         (pe_mat_18_30_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_18_30_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_18_30_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_18_31_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_18_31_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_18_31_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_17_31_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_17_31_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_18_31_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_18_31_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_19_0 (
    .io_in_r_data         (io_in_r_19_data[15:0]           ), //i
    .io_in_r_stop_weight  (io_in_r_19_stop_weight          ), //i
    .io_in_r_stall        (io_in_r_19_stall                ), //i
    .io_out_r_data        (pe_mat_19_0_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_19_0_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_19_0_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_18_0_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_18_0_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_19_0_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_19_0_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_19_1 (
    .io_in_r_data         (pe_mat_19_0_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_19_0_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_19_0_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_19_1_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_19_1_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_19_1_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_18_1_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_18_1_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_19_1_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_19_1_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_19_2 (
    .io_in_r_data         (pe_mat_19_1_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_19_1_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_19_1_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_19_2_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_19_2_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_19_2_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_18_2_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_18_2_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_19_2_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_19_2_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_19_3 (
    .io_in_r_data         (pe_mat_19_2_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_19_2_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_19_2_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_19_3_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_19_3_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_19_3_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_18_3_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_18_3_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_19_3_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_19_3_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_19_4 (
    .io_in_r_data         (pe_mat_19_3_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_19_3_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_19_3_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_19_4_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_19_4_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_19_4_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_18_4_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_18_4_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_19_4_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_19_4_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_19_5 (
    .io_in_r_data         (pe_mat_19_4_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_19_4_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_19_4_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_19_5_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_19_5_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_19_5_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_18_5_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_18_5_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_19_5_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_19_5_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_19_6 (
    .io_in_r_data         (pe_mat_19_5_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_19_5_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_19_5_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_19_6_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_19_6_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_19_6_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_18_6_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_18_6_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_19_6_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_19_6_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_19_7 (
    .io_in_r_data         (pe_mat_19_6_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_19_6_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_19_6_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_19_7_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_19_7_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_19_7_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_18_7_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_18_7_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_19_7_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_19_7_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_19_8 (
    .io_in_r_data         (pe_mat_19_7_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_19_7_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_19_7_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_19_8_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_19_8_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_19_8_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_18_8_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_18_8_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_19_8_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_19_8_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_19_9 (
    .io_in_r_data         (pe_mat_19_8_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_19_8_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_19_8_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_19_9_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_19_9_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_19_9_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_18_9_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_18_9_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_19_9_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_19_9_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_19_10 (
    .io_in_r_data         (pe_mat_19_9_io_out_r_data[15:0]  ), //i
    .io_in_r_stop_weight  (pe_mat_19_9_io_out_r_stop_weight ), //i
    .io_in_r_stall        (pe_mat_19_9_io_out_r_stall       ), //i
    .io_out_r_data        (pe_mat_19_10_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_19_10_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_19_10_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_18_10_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_18_10_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_19_10_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_19_10_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_19_11 (
    .io_in_r_data         (pe_mat_19_10_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_19_10_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_19_10_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_19_11_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_19_11_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_19_11_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_18_11_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_18_11_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_19_11_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_19_11_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_19_12 (
    .io_in_r_data         (pe_mat_19_11_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_19_11_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_19_11_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_19_12_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_19_12_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_19_12_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_18_12_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_18_12_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_19_12_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_19_12_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_19_13 (
    .io_in_r_data         (pe_mat_19_12_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_19_12_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_19_12_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_19_13_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_19_13_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_19_13_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_18_13_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_18_13_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_19_13_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_19_13_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_19_14 (
    .io_in_r_data         (pe_mat_19_13_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_19_13_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_19_13_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_19_14_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_19_14_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_19_14_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_18_14_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_18_14_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_19_14_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_19_14_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_19_15 (
    .io_in_r_data         (pe_mat_19_14_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_19_14_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_19_14_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_19_15_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_19_15_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_19_15_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_18_15_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_18_15_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_19_15_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_19_15_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_19_16 (
    .io_in_r_data         (pe_mat_19_15_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_19_15_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_19_15_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_19_16_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_19_16_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_19_16_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_18_16_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_18_16_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_19_16_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_19_16_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_19_17 (
    .io_in_r_data         (pe_mat_19_16_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_19_16_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_19_16_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_19_17_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_19_17_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_19_17_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_18_17_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_18_17_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_19_17_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_19_17_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_19_18 (
    .io_in_r_data         (pe_mat_19_17_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_19_17_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_19_17_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_19_18_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_19_18_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_19_18_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_18_18_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_18_18_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_19_18_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_19_18_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_19_19 (
    .io_in_r_data         (pe_mat_19_18_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_19_18_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_19_18_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_19_19_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_19_19_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_19_19_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_18_19_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_18_19_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_19_19_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_19_19_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_19_20 (
    .io_in_r_data         (pe_mat_19_19_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_19_19_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_19_19_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_19_20_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_19_20_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_19_20_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_18_20_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_18_20_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_19_20_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_19_20_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_19_21 (
    .io_in_r_data         (pe_mat_19_20_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_19_20_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_19_20_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_19_21_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_19_21_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_19_21_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_18_21_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_18_21_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_19_21_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_19_21_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_19_22 (
    .io_in_r_data         (pe_mat_19_21_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_19_21_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_19_21_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_19_22_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_19_22_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_19_22_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_18_22_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_18_22_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_19_22_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_19_22_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_19_23 (
    .io_in_r_data         (pe_mat_19_22_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_19_22_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_19_22_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_19_23_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_19_23_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_19_23_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_18_23_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_18_23_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_19_23_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_19_23_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_19_24 (
    .io_in_r_data         (pe_mat_19_23_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_19_23_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_19_23_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_19_24_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_19_24_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_19_24_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_18_24_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_18_24_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_19_24_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_19_24_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_19_25 (
    .io_in_r_data         (pe_mat_19_24_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_19_24_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_19_24_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_19_25_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_19_25_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_19_25_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_18_25_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_18_25_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_19_25_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_19_25_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_19_26 (
    .io_in_r_data         (pe_mat_19_25_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_19_25_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_19_25_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_19_26_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_19_26_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_19_26_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_18_26_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_18_26_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_19_26_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_19_26_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_19_27 (
    .io_in_r_data         (pe_mat_19_26_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_19_26_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_19_26_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_19_27_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_19_27_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_19_27_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_18_27_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_18_27_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_19_27_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_19_27_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_19_28 (
    .io_in_r_data         (pe_mat_19_27_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_19_27_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_19_27_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_19_28_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_19_28_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_19_28_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_18_28_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_18_28_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_19_28_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_19_28_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_19_29 (
    .io_in_r_data         (pe_mat_19_28_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_19_28_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_19_28_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_19_29_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_19_29_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_19_29_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_18_29_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_18_29_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_19_29_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_19_29_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_19_30 (
    .io_in_r_data         (pe_mat_19_29_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_19_29_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_19_29_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_19_30_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_19_30_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_19_30_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_18_30_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_18_30_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_19_30_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_19_30_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_19_31 (
    .io_in_r_data         (pe_mat_19_30_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_19_30_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_19_30_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_19_31_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_19_31_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_19_31_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_18_31_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_18_31_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_19_31_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_19_31_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_20_0 (
    .io_in_r_data         (io_in_r_20_data[15:0]           ), //i
    .io_in_r_stop_weight  (io_in_r_20_stop_weight          ), //i
    .io_in_r_stall        (io_in_r_20_stall                ), //i
    .io_out_r_data        (pe_mat_20_0_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_20_0_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_20_0_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_19_0_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_19_0_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_20_0_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_20_0_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_20_1 (
    .io_in_r_data         (pe_mat_20_0_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_20_0_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_20_0_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_20_1_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_20_1_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_20_1_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_19_1_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_19_1_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_20_1_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_20_1_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_20_2 (
    .io_in_r_data         (pe_mat_20_1_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_20_1_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_20_1_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_20_2_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_20_2_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_20_2_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_19_2_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_19_2_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_20_2_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_20_2_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_20_3 (
    .io_in_r_data         (pe_mat_20_2_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_20_2_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_20_2_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_20_3_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_20_3_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_20_3_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_19_3_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_19_3_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_20_3_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_20_3_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_20_4 (
    .io_in_r_data         (pe_mat_20_3_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_20_3_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_20_3_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_20_4_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_20_4_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_20_4_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_19_4_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_19_4_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_20_4_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_20_4_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_20_5 (
    .io_in_r_data         (pe_mat_20_4_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_20_4_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_20_4_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_20_5_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_20_5_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_20_5_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_19_5_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_19_5_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_20_5_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_20_5_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_20_6 (
    .io_in_r_data         (pe_mat_20_5_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_20_5_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_20_5_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_20_6_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_20_6_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_20_6_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_19_6_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_19_6_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_20_6_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_20_6_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_20_7 (
    .io_in_r_data         (pe_mat_20_6_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_20_6_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_20_6_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_20_7_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_20_7_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_20_7_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_19_7_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_19_7_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_20_7_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_20_7_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_20_8 (
    .io_in_r_data         (pe_mat_20_7_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_20_7_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_20_7_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_20_8_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_20_8_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_20_8_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_19_8_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_19_8_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_20_8_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_20_8_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_20_9 (
    .io_in_r_data         (pe_mat_20_8_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_20_8_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_20_8_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_20_9_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_20_9_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_20_9_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_19_9_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_19_9_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_20_9_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_20_9_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_20_10 (
    .io_in_r_data         (pe_mat_20_9_io_out_r_data[15:0]  ), //i
    .io_in_r_stop_weight  (pe_mat_20_9_io_out_r_stop_weight ), //i
    .io_in_r_stall        (pe_mat_20_9_io_out_r_stall       ), //i
    .io_out_r_data        (pe_mat_20_10_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_20_10_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_20_10_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_19_10_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_19_10_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_20_10_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_20_10_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_20_11 (
    .io_in_r_data         (pe_mat_20_10_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_20_10_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_20_10_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_20_11_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_20_11_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_20_11_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_19_11_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_19_11_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_20_11_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_20_11_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_20_12 (
    .io_in_r_data         (pe_mat_20_11_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_20_11_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_20_11_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_20_12_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_20_12_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_20_12_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_19_12_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_19_12_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_20_12_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_20_12_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_20_13 (
    .io_in_r_data         (pe_mat_20_12_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_20_12_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_20_12_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_20_13_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_20_13_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_20_13_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_19_13_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_19_13_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_20_13_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_20_13_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_20_14 (
    .io_in_r_data         (pe_mat_20_13_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_20_13_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_20_13_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_20_14_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_20_14_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_20_14_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_19_14_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_19_14_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_20_14_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_20_14_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_20_15 (
    .io_in_r_data         (pe_mat_20_14_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_20_14_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_20_14_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_20_15_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_20_15_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_20_15_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_19_15_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_19_15_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_20_15_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_20_15_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_20_16 (
    .io_in_r_data         (pe_mat_20_15_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_20_15_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_20_15_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_20_16_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_20_16_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_20_16_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_19_16_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_19_16_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_20_16_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_20_16_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_20_17 (
    .io_in_r_data         (pe_mat_20_16_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_20_16_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_20_16_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_20_17_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_20_17_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_20_17_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_19_17_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_19_17_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_20_17_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_20_17_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_20_18 (
    .io_in_r_data         (pe_mat_20_17_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_20_17_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_20_17_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_20_18_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_20_18_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_20_18_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_19_18_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_19_18_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_20_18_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_20_18_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_20_19 (
    .io_in_r_data         (pe_mat_20_18_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_20_18_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_20_18_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_20_19_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_20_19_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_20_19_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_19_19_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_19_19_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_20_19_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_20_19_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_20_20 (
    .io_in_r_data         (pe_mat_20_19_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_20_19_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_20_19_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_20_20_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_20_20_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_20_20_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_19_20_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_19_20_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_20_20_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_20_20_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_20_21 (
    .io_in_r_data         (pe_mat_20_20_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_20_20_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_20_20_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_20_21_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_20_21_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_20_21_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_19_21_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_19_21_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_20_21_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_20_21_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_20_22 (
    .io_in_r_data         (pe_mat_20_21_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_20_21_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_20_21_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_20_22_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_20_22_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_20_22_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_19_22_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_19_22_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_20_22_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_20_22_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_20_23 (
    .io_in_r_data         (pe_mat_20_22_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_20_22_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_20_22_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_20_23_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_20_23_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_20_23_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_19_23_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_19_23_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_20_23_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_20_23_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_20_24 (
    .io_in_r_data         (pe_mat_20_23_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_20_23_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_20_23_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_20_24_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_20_24_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_20_24_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_19_24_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_19_24_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_20_24_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_20_24_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_20_25 (
    .io_in_r_data         (pe_mat_20_24_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_20_24_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_20_24_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_20_25_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_20_25_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_20_25_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_19_25_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_19_25_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_20_25_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_20_25_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_20_26 (
    .io_in_r_data         (pe_mat_20_25_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_20_25_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_20_25_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_20_26_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_20_26_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_20_26_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_19_26_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_19_26_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_20_26_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_20_26_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_20_27 (
    .io_in_r_data         (pe_mat_20_26_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_20_26_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_20_26_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_20_27_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_20_27_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_20_27_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_19_27_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_19_27_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_20_27_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_20_27_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_20_28 (
    .io_in_r_data         (pe_mat_20_27_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_20_27_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_20_27_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_20_28_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_20_28_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_20_28_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_19_28_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_19_28_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_20_28_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_20_28_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_20_29 (
    .io_in_r_data         (pe_mat_20_28_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_20_28_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_20_28_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_20_29_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_20_29_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_20_29_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_19_29_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_19_29_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_20_29_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_20_29_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_20_30 (
    .io_in_r_data         (pe_mat_20_29_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_20_29_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_20_29_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_20_30_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_20_30_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_20_30_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_19_30_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_19_30_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_20_30_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_20_30_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_20_31 (
    .io_in_r_data         (pe_mat_20_30_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_20_30_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_20_30_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_20_31_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_20_31_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_20_31_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_19_31_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_19_31_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_20_31_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_20_31_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_21_0 (
    .io_in_r_data         (io_in_r_21_data[15:0]           ), //i
    .io_in_r_stop_weight  (io_in_r_21_stop_weight          ), //i
    .io_in_r_stall        (io_in_r_21_stall                ), //i
    .io_out_r_data        (pe_mat_21_0_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_21_0_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_21_0_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_20_0_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_20_0_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_21_0_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_21_0_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_21_1 (
    .io_in_r_data         (pe_mat_21_0_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_21_0_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_21_0_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_21_1_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_21_1_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_21_1_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_20_1_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_20_1_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_21_1_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_21_1_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_21_2 (
    .io_in_r_data         (pe_mat_21_1_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_21_1_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_21_1_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_21_2_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_21_2_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_21_2_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_20_2_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_20_2_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_21_2_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_21_2_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_21_3 (
    .io_in_r_data         (pe_mat_21_2_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_21_2_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_21_2_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_21_3_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_21_3_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_21_3_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_20_3_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_20_3_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_21_3_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_21_3_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_21_4 (
    .io_in_r_data         (pe_mat_21_3_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_21_3_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_21_3_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_21_4_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_21_4_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_21_4_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_20_4_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_20_4_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_21_4_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_21_4_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_21_5 (
    .io_in_r_data         (pe_mat_21_4_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_21_4_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_21_4_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_21_5_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_21_5_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_21_5_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_20_5_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_20_5_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_21_5_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_21_5_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_21_6 (
    .io_in_r_data         (pe_mat_21_5_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_21_5_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_21_5_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_21_6_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_21_6_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_21_6_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_20_6_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_20_6_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_21_6_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_21_6_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_21_7 (
    .io_in_r_data         (pe_mat_21_6_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_21_6_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_21_6_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_21_7_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_21_7_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_21_7_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_20_7_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_20_7_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_21_7_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_21_7_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_21_8 (
    .io_in_r_data         (pe_mat_21_7_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_21_7_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_21_7_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_21_8_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_21_8_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_21_8_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_20_8_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_20_8_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_21_8_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_21_8_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_21_9 (
    .io_in_r_data         (pe_mat_21_8_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_21_8_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_21_8_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_21_9_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_21_9_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_21_9_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_20_9_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_20_9_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_21_9_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_21_9_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_21_10 (
    .io_in_r_data         (pe_mat_21_9_io_out_r_data[15:0]  ), //i
    .io_in_r_stop_weight  (pe_mat_21_9_io_out_r_stop_weight ), //i
    .io_in_r_stall        (pe_mat_21_9_io_out_r_stall       ), //i
    .io_out_r_data        (pe_mat_21_10_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_21_10_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_21_10_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_20_10_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_20_10_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_21_10_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_21_10_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_21_11 (
    .io_in_r_data         (pe_mat_21_10_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_21_10_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_21_10_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_21_11_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_21_11_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_21_11_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_20_11_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_20_11_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_21_11_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_21_11_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_21_12 (
    .io_in_r_data         (pe_mat_21_11_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_21_11_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_21_11_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_21_12_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_21_12_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_21_12_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_20_12_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_20_12_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_21_12_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_21_12_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_21_13 (
    .io_in_r_data         (pe_mat_21_12_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_21_12_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_21_12_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_21_13_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_21_13_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_21_13_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_20_13_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_20_13_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_21_13_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_21_13_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_21_14 (
    .io_in_r_data         (pe_mat_21_13_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_21_13_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_21_13_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_21_14_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_21_14_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_21_14_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_20_14_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_20_14_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_21_14_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_21_14_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_21_15 (
    .io_in_r_data         (pe_mat_21_14_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_21_14_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_21_14_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_21_15_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_21_15_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_21_15_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_20_15_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_20_15_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_21_15_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_21_15_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_21_16 (
    .io_in_r_data         (pe_mat_21_15_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_21_15_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_21_15_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_21_16_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_21_16_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_21_16_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_20_16_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_20_16_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_21_16_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_21_16_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_21_17 (
    .io_in_r_data         (pe_mat_21_16_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_21_16_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_21_16_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_21_17_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_21_17_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_21_17_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_20_17_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_20_17_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_21_17_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_21_17_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_21_18 (
    .io_in_r_data         (pe_mat_21_17_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_21_17_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_21_17_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_21_18_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_21_18_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_21_18_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_20_18_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_20_18_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_21_18_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_21_18_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_21_19 (
    .io_in_r_data         (pe_mat_21_18_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_21_18_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_21_18_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_21_19_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_21_19_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_21_19_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_20_19_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_20_19_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_21_19_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_21_19_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_21_20 (
    .io_in_r_data         (pe_mat_21_19_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_21_19_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_21_19_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_21_20_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_21_20_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_21_20_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_20_20_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_20_20_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_21_20_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_21_20_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_21_21 (
    .io_in_r_data         (pe_mat_21_20_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_21_20_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_21_20_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_21_21_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_21_21_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_21_21_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_20_21_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_20_21_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_21_21_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_21_21_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_21_22 (
    .io_in_r_data         (pe_mat_21_21_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_21_21_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_21_21_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_21_22_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_21_22_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_21_22_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_20_22_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_20_22_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_21_22_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_21_22_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_21_23 (
    .io_in_r_data         (pe_mat_21_22_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_21_22_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_21_22_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_21_23_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_21_23_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_21_23_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_20_23_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_20_23_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_21_23_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_21_23_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_21_24 (
    .io_in_r_data         (pe_mat_21_23_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_21_23_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_21_23_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_21_24_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_21_24_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_21_24_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_20_24_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_20_24_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_21_24_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_21_24_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_21_25 (
    .io_in_r_data         (pe_mat_21_24_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_21_24_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_21_24_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_21_25_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_21_25_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_21_25_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_20_25_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_20_25_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_21_25_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_21_25_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_21_26 (
    .io_in_r_data         (pe_mat_21_25_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_21_25_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_21_25_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_21_26_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_21_26_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_21_26_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_20_26_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_20_26_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_21_26_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_21_26_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_21_27 (
    .io_in_r_data         (pe_mat_21_26_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_21_26_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_21_26_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_21_27_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_21_27_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_21_27_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_20_27_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_20_27_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_21_27_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_21_27_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_21_28 (
    .io_in_r_data         (pe_mat_21_27_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_21_27_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_21_27_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_21_28_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_21_28_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_21_28_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_20_28_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_20_28_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_21_28_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_21_28_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_21_29 (
    .io_in_r_data         (pe_mat_21_28_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_21_28_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_21_28_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_21_29_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_21_29_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_21_29_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_20_29_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_20_29_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_21_29_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_21_29_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_21_30 (
    .io_in_r_data         (pe_mat_21_29_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_21_29_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_21_29_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_21_30_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_21_30_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_21_30_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_20_30_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_20_30_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_21_30_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_21_30_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_21_31 (
    .io_in_r_data         (pe_mat_21_30_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_21_30_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_21_30_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_21_31_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_21_31_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_21_31_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_20_31_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_20_31_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_21_31_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_21_31_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_22_0 (
    .io_in_r_data         (io_in_r_22_data[15:0]           ), //i
    .io_in_r_stop_weight  (io_in_r_22_stop_weight          ), //i
    .io_in_r_stall        (io_in_r_22_stall                ), //i
    .io_out_r_data        (pe_mat_22_0_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_22_0_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_22_0_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_21_0_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_21_0_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_22_0_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_22_0_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_22_1 (
    .io_in_r_data         (pe_mat_22_0_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_22_0_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_22_0_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_22_1_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_22_1_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_22_1_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_21_1_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_21_1_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_22_1_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_22_1_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_22_2 (
    .io_in_r_data         (pe_mat_22_1_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_22_1_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_22_1_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_22_2_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_22_2_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_22_2_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_21_2_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_21_2_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_22_2_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_22_2_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_22_3 (
    .io_in_r_data         (pe_mat_22_2_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_22_2_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_22_2_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_22_3_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_22_3_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_22_3_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_21_3_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_21_3_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_22_3_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_22_3_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_22_4 (
    .io_in_r_data         (pe_mat_22_3_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_22_3_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_22_3_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_22_4_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_22_4_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_22_4_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_21_4_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_21_4_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_22_4_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_22_4_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_22_5 (
    .io_in_r_data         (pe_mat_22_4_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_22_4_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_22_4_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_22_5_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_22_5_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_22_5_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_21_5_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_21_5_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_22_5_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_22_5_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_22_6 (
    .io_in_r_data         (pe_mat_22_5_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_22_5_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_22_5_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_22_6_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_22_6_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_22_6_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_21_6_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_21_6_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_22_6_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_22_6_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_22_7 (
    .io_in_r_data         (pe_mat_22_6_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_22_6_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_22_6_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_22_7_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_22_7_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_22_7_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_21_7_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_21_7_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_22_7_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_22_7_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_22_8 (
    .io_in_r_data         (pe_mat_22_7_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_22_7_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_22_7_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_22_8_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_22_8_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_22_8_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_21_8_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_21_8_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_22_8_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_22_8_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_22_9 (
    .io_in_r_data         (pe_mat_22_8_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_22_8_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_22_8_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_22_9_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_22_9_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_22_9_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_21_9_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_21_9_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_22_9_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_22_9_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_22_10 (
    .io_in_r_data         (pe_mat_22_9_io_out_r_data[15:0]  ), //i
    .io_in_r_stop_weight  (pe_mat_22_9_io_out_r_stop_weight ), //i
    .io_in_r_stall        (pe_mat_22_9_io_out_r_stall       ), //i
    .io_out_r_data        (pe_mat_22_10_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_22_10_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_22_10_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_21_10_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_21_10_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_22_10_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_22_10_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_22_11 (
    .io_in_r_data         (pe_mat_22_10_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_22_10_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_22_10_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_22_11_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_22_11_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_22_11_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_21_11_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_21_11_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_22_11_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_22_11_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_22_12 (
    .io_in_r_data         (pe_mat_22_11_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_22_11_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_22_11_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_22_12_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_22_12_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_22_12_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_21_12_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_21_12_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_22_12_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_22_12_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_22_13 (
    .io_in_r_data         (pe_mat_22_12_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_22_12_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_22_12_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_22_13_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_22_13_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_22_13_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_21_13_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_21_13_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_22_13_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_22_13_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_22_14 (
    .io_in_r_data         (pe_mat_22_13_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_22_13_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_22_13_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_22_14_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_22_14_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_22_14_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_21_14_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_21_14_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_22_14_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_22_14_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_22_15 (
    .io_in_r_data         (pe_mat_22_14_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_22_14_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_22_14_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_22_15_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_22_15_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_22_15_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_21_15_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_21_15_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_22_15_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_22_15_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_22_16 (
    .io_in_r_data         (pe_mat_22_15_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_22_15_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_22_15_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_22_16_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_22_16_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_22_16_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_21_16_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_21_16_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_22_16_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_22_16_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_22_17 (
    .io_in_r_data         (pe_mat_22_16_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_22_16_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_22_16_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_22_17_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_22_17_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_22_17_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_21_17_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_21_17_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_22_17_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_22_17_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_22_18 (
    .io_in_r_data         (pe_mat_22_17_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_22_17_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_22_17_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_22_18_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_22_18_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_22_18_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_21_18_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_21_18_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_22_18_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_22_18_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_22_19 (
    .io_in_r_data         (pe_mat_22_18_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_22_18_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_22_18_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_22_19_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_22_19_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_22_19_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_21_19_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_21_19_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_22_19_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_22_19_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_22_20 (
    .io_in_r_data         (pe_mat_22_19_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_22_19_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_22_19_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_22_20_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_22_20_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_22_20_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_21_20_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_21_20_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_22_20_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_22_20_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_22_21 (
    .io_in_r_data         (pe_mat_22_20_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_22_20_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_22_20_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_22_21_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_22_21_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_22_21_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_21_21_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_21_21_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_22_21_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_22_21_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_22_22 (
    .io_in_r_data         (pe_mat_22_21_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_22_21_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_22_21_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_22_22_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_22_22_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_22_22_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_21_22_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_21_22_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_22_22_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_22_22_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_22_23 (
    .io_in_r_data         (pe_mat_22_22_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_22_22_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_22_22_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_22_23_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_22_23_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_22_23_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_21_23_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_21_23_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_22_23_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_22_23_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_22_24 (
    .io_in_r_data         (pe_mat_22_23_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_22_23_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_22_23_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_22_24_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_22_24_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_22_24_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_21_24_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_21_24_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_22_24_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_22_24_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_22_25 (
    .io_in_r_data         (pe_mat_22_24_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_22_24_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_22_24_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_22_25_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_22_25_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_22_25_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_21_25_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_21_25_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_22_25_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_22_25_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_22_26 (
    .io_in_r_data         (pe_mat_22_25_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_22_25_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_22_25_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_22_26_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_22_26_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_22_26_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_21_26_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_21_26_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_22_26_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_22_26_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_22_27 (
    .io_in_r_data         (pe_mat_22_26_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_22_26_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_22_26_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_22_27_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_22_27_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_22_27_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_21_27_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_21_27_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_22_27_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_22_27_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_22_28 (
    .io_in_r_data         (pe_mat_22_27_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_22_27_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_22_27_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_22_28_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_22_28_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_22_28_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_21_28_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_21_28_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_22_28_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_22_28_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_22_29 (
    .io_in_r_data         (pe_mat_22_28_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_22_28_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_22_28_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_22_29_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_22_29_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_22_29_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_21_29_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_21_29_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_22_29_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_22_29_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_22_30 (
    .io_in_r_data         (pe_mat_22_29_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_22_29_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_22_29_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_22_30_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_22_30_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_22_30_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_21_30_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_21_30_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_22_30_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_22_30_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_22_31 (
    .io_in_r_data         (pe_mat_22_30_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_22_30_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_22_30_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_22_31_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_22_31_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_22_31_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_21_31_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_21_31_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_22_31_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_22_31_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_23_0 (
    .io_in_r_data         (io_in_r_23_data[15:0]           ), //i
    .io_in_r_stop_weight  (io_in_r_23_stop_weight          ), //i
    .io_in_r_stall        (io_in_r_23_stall                ), //i
    .io_out_r_data        (pe_mat_23_0_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_23_0_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_23_0_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_22_0_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_22_0_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_23_0_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_23_0_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_23_1 (
    .io_in_r_data         (pe_mat_23_0_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_23_0_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_23_0_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_23_1_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_23_1_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_23_1_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_22_1_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_22_1_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_23_1_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_23_1_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_23_2 (
    .io_in_r_data         (pe_mat_23_1_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_23_1_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_23_1_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_23_2_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_23_2_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_23_2_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_22_2_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_22_2_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_23_2_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_23_2_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_23_3 (
    .io_in_r_data         (pe_mat_23_2_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_23_2_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_23_2_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_23_3_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_23_3_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_23_3_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_22_3_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_22_3_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_23_3_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_23_3_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_23_4 (
    .io_in_r_data         (pe_mat_23_3_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_23_3_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_23_3_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_23_4_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_23_4_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_23_4_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_22_4_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_22_4_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_23_4_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_23_4_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_23_5 (
    .io_in_r_data         (pe_mat_23_4_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_23_4_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_23_4_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_23_5_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_23_5_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_23_5_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_22_5_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_22_5_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_23_5_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_23_5_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_23_6 (
    .io_in_r_data         (pe_mat_23_5_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_23_5_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_23_5_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_23_6_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_23_6_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_23_6_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_22_6_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_22_6_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_23_6_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_23_6_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_23_7 (
    .io_in_r_data         (pe_mat_23_6_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_23_6_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_23_6_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_23_7_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_23_7_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_23_7_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_22_7_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_22_7_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_23_7_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_23_7_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_23_8 (
    .io_in_r_data         (pe_mat_23_7_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_23_7_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_23_7_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_23_8_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_23_8_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_23_8_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_22_8_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_22_8_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_23_8_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_23_8_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_23_9 (
    .io_in_r_data         (pe_mat_23_8_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_23_8_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_23_8_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_23_9_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_23_9_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_23_9_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_22_9_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_22_9_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_23_9_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_23_9_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_23_10 (
    .io_in_r_data         (pe_mat_23_9_io_out_r_data[15:0]  ), //i
    .io_in_r_stop_weight  (pe_mat_23_9_io_out_r_stop_weight ), //i
    .io_in_r_stall        (pe_mat_23_9_io_out_r_stall       ), //i
    .io_out_r_data        (pe_mat_23_10_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_23_10_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_23_10_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_22_10_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_22_10_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_23_10_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_23_10_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_23_11 (
    .io_in_r_data         (pe_mat_23_10_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_23_10_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_23_10_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_23_11_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_23_11_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_23_11_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_22_11_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_22_11_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_23_11_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_23_11_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_23_12 (
    .io_in_r_data         (pe_mat_23_11_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_23_11_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_23_11_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_23_12_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_23_12_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_23_12_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_22_12_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_22_12_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_23_12_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_23_12_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_23_13 (
    .io_in_r_data         (pe_mat_23_12_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_23_12_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_23_12_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_23_13_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_23_13_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_23_13_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_22_13_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_22_13_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_23_13_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_23_13_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_23_14 (
    .io_in_r_data         (pe_mat_23_13_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_23_13_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_23_13_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_23_14_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_23_14_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_23_14_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_22_14_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_22_14_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_23_14_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_23_14_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_23_15 (
    .io_in_r_data         (pe_mat_23_14_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_23_14_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_23_14_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_23_15_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_23_15_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_23_15_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_22_15_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_22_15_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_23_15_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_23_15_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_23_16 (
    .io_in_r_data         (pe_mat_23_15_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_23_15_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_23_15_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_23_16_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_23_16_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_23_16_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_22_16_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_22_16_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_23_16_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_23_16_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_23_17 (
    .io_in_r_data         (pe_mat_23_16_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_23_16_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_23_16_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_23_17_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_23_17_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_23_17_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_22_17_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_22_17_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_23_17_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_23_17_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_23_18 (
    .io_in_r_data         (pe_mat_23_17_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_23_17_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_23_17_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_23_18_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_23_18_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_23_18_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_22_18_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_22_18_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_23_18_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_23_18_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_23_19 (
    .io_in_r_data         (pe_mat_23_18_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_23_18_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_23_18_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_23_19_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_23_19_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_23_19_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_22_19_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_22_19_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_23_19_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_23_19_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_23_20 (
    .io_in_r_data         (pe_mat_23_19_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_23_19_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_23_19_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_23_20_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_23_20_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_23_20_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_22_20_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_22_20_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_23_20_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_23_20_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_23_21 (
    .io_in_r_data         (pe_mat_23_20_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_23_20_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_23_20_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_23_21_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_23_21_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_23_21_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_22_21_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_22_21_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_23_21_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_23_21_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_23_22 (
    .io_in_r_data         (pe_mat_23_21_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_23_21_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_23_21_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_23_22_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_23_22_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_23_22_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_22_22_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_22_22_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_23_22_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_23_22_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_23_23 (
    .io_in_r_data         (pe_mat_23_22_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_23_22_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_23_22_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_23_23_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_23_23_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_23_23_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_22_23_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_22_23_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_23_23_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_23_23_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_23_24 (
    .io_in_r_data         (pe_mat_23_23_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_23_23_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_23_23_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_23_24_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_23_24_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_23_24_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_22_24_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_22_24_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_23_24_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_23_24_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_23_25 (
    .io_in_r_data         (pe_mat_23_24_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_23_24_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_23_24_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_23_25_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_23_25_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_23_25_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_22_25_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_22_25_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_23_25_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_23_25_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_23_26 (
    .io_in_r_data         (pe_mat_23_25_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_23_25_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_23_25_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_23_26_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_23_26_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_23_26_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_22_26_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_22_26_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_23_26_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_23_26_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_23_27 (
    .io_in_r_data         (pe_mat_23_26_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_23_26_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_23_26_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_23_27_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_23_27_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_23_27_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_22_27_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_22_27_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_23_27_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_23_27_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_23_28 (
    .io_in_r_data         (pe_mat_23_27_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_23_27_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_23_27_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_23_28_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_23_28_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_23_28_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_22_28_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_22_28_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_23_28_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_23_28_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_23_29 (
    .io_in_r_data         (pe_mat_23_28_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_23_28_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_23_28_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_23_29_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_23_29_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_23_29_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_22_29_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_22_29_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_23_29_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_23_29_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_23_30 (
    .io_in_r_data         (pe_mat_23_29_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_23_29_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_23_29_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_23_30_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_23_30_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_23_30_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_22_30_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_22_30_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_23_30_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_23_30_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_23_31 (
    .io_in_r_data         (pe_mat_23_30_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_23_30_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_23_30_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_23_31_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_23_31_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_23_31_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_22_31_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_22_31_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_23_31_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_23_31_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_24_0 (
    .io_in_r_data         (io_in_r_24_data[15:0]           ), //i
    .io_in_r_stop_weight  (io_in_r_24_stop_weight          ), //i
    .io_in_r_stall        (io_in_r_24_stall                ), //i
    .io_out_r_data        (pe_mat_24_0_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_24_0_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_24_0_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_23_0_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_23_0_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_24_0_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_24_0_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_24_1 (
    .io_in_r_data         (pe_mat_24_0_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_24_0_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_24_0_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_24_1_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_24_1_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_24_1_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_23_1_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_23_1_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_24_1_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_24_1_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_24_2 (
    .io_in_r_data         (pe_mat_24_1_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_24_1_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_24_1_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_24_2_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_24_2_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_24_2_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_23_2_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_23_2_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_24_2_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_24_2_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_24_3 (
    .io_in_r_data         (pe_mat_24_2_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_24_2_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_24_2_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_24_3_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_24_3_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_24_3_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_23_3_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_23_3_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_24_3_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_24_3_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_24_4 (
    .io_in_r_data         (pe_mat_24_3_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_24_3_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_24_3_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_24_4_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_24_4_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_24_4_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_23_4_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_23_4_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_24_4_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_24_4_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_24_5 (
    .io_in_r_data         (pe_mat_24_4_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_24_4_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_24_4_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_24_5_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_24_5_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_24_5_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_23_5_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_23_5_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_24_5_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_24_5_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_24_6 (
    .io_in_r_data         (pe_mat_24_5_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_24_5_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_24_5_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_24_6_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_24_6_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_24_6_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_23_6_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_23_6_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_24_6_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_24_6_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_24_7 (
    .io_in_r_data         (pe_mat_24_6_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_24_6_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_24_6_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_24_7_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_24_7_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_24_7_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_23_7_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_23_7_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_24_7_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_24_7_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_24_8 (
    .io_in_r_data         (pe_mat_24_7_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_24_7_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_24_7_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_24_8_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_24_8_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_24_8_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_23_8_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_23_8_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_24_8_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_24_8_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_24_9 (
    .io_in_r_data         (pe_mat_24_8_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_24_8_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_24_8_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_24_9_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_24_9_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_24_9_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_23_9_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_23_9_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_24_9_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_24_9_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_24_10 (
    .io_in_r_data         (pe_mat_24_9_io_out_r_data[15:0]  ), //i
    .io_in_r_stop_weight  (pe_mat_24_9_io_out_r_stop_weight ), //i
    .io_in_r_stall        (pe_mat_24_9_io_out_r_stall       ), //i
    .io_out_r_data        (pe_mat_24_10_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_24_10_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_24_10_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_23_10_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_23_10_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_24_10_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_24_10_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_24_11 (
    .io_in_r_data         (pe_mat_24_10_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_24_10_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_24_10_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_24_11_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_24_11_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_24_11_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_23_11_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_23_11_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_24_11_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_24_11_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_24_12 (
    .io_in_r_data         (pe_mat_24_11_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_24_11_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_24_11_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_24_12_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_24_12_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_24_12_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_23_12_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_23_12_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_24_12_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_24_12_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_24_13 (
    .io_in_r_data         (pe_mat_24_12_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_24_12_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_24_12_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_24_13_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_24_13_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_24_13_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_23_13_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_23_13_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_24_13_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_24_13_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_24_14 (
    .io_in_r_data         (pe_mat_24_13_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_24_13_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_24_13_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_24_14_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_24_14_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_24_14_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_23_14_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_23_14_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_24_14_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_24_14_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_24_15 (
    .io_in_r_data         (pe_mat_24_14_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_24_14_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_24_14_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_24_15_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_24_15_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_24_15_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_23_15_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_23_15_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_24_15_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_24_15_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_24_16 (
    .io_in_r_data         (pe_mat_24_15_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_24_15_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_24_15_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_24_16_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_24_16_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_24_16_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_23_16_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_23_16_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_24_16_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_24_16_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_24_17 (
    .io_in_r_data         (pe_mat_24_16_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_24_16_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_24_16_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_24_17_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_24_17_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_24_17_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_23_17_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_23_17_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_24_17_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_24_17_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_24_18 (
    .io_in_r_data         (pe_mat_24_17_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_24_17_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_24_17_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_24_18_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_24_18_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_24_18_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_23_18_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_23_18_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_24_18_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_24_18_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_24_19 (
    .io_in_r_data         (pe_mat_24_18_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_24_18_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_24_18_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_24_19_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_24_19_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_24_19_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_23_19_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_23_19_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_24_19_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_24_19_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_24_20 (
    .io_in_r_data         (pe_mat_24_19_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_24_19_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_24_19_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_24_20_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_24_20_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_24_20_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_23_20_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_23_20_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_24_20_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_24_20_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_24_21 (
    .io_in_r_data         (pe_mat_24_20_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_24_20_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_24_20_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_24_21_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_24_21_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_24_21_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_23_21_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_23_21_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_24_21_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_24_21_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_24_22 (
    .io_in_r_data         (pe_mat_24_21_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_24_21_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_24_21_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_24_22_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_24_22_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_24_22_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_23_22_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_23_22_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_24_22_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_24_22_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_24_23 (
    .io_in_r_data         (pe_mat_24_22_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_24_22_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_24_22_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_24_23_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_24_23_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_24_23_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_23_23_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_23_23_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_24_23_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_24_23_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_24_24 (
    .io_in_r_data         (pe_mat_24_23_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_24_23_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_24_23_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_24_24_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_24_24_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_24_24_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_23_24_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_23_24_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_24_24_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_24_24_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_24_25 (
    .io_in_r_data         (pe_mat_24_24_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_24_24_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_24_24_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_24_25_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_24_25_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_24_25_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_23_25_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_23_25_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_24_25_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_24_25_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_24_26 (
    .io_in_r_data         (pe_mat_24_25_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_24_25_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_24_25_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_24_26_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_24_26_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_24_26_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_23_26_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_23_26_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_24_26_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_24_26_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_24_27 (
    .io_in_r_data         (pe_mat_24_26_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_24_26_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_24_26_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_24_27_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_24_27_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_24_27_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_23_27_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_23_27_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_24_27_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_24_27_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_24_28 (
    .io_in_r_data         (pe_mat_24_27_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_24_27_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_24_27_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_24_28_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_24_28_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_24_28_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_23_28_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_23_28_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_24_28_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_24_28_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_24_29 (
    .io_in_r_data         (pe_mat_24_28_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_24_28_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_24_28_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_24_29_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_24_29_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_24_29_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_23_29_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_23_29_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_24_29_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_24_29_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_24_30 (
    .io_in_r_data         (pe_mat_24_29_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_24_29_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_24_29_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_24_30_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_24_30_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_24_30_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_23_30_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_23_30_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_24_30_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_24_30_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_24_31 (
    .io_in_r_data         (pe_mat_24_30_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_24_30_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_24_30_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_24_31_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_24_31_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_24_31_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_23_31_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_23_31_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_24_31_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_24_31_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_25_0 (
    .io_in_r_data         (io_in_r_25_data[15:0]           ), //i
    .io_in_r_stop_weight  (io_in_r_25_stop_weight          ), //i
    .io_in_r_stall        (io_in_r_25_stall                ), //i
    .io_out_r_data        (pe_mat_25_0_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_25_0_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_25_0_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_24_0_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_24_0_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_25_0_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_25_0_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_25_1 (
    .io_in_r_data         (pe_mat_25_0_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_25_0_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_25_0_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_25_1_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_25_1_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_25_1_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_24_1_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_24_1_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_25_1_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_25_1_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_25_2 (
    .io_in_r_data         (pe_mat_25_1_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_25_1_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_25_1_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_25_2_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_25_2_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_25_2_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_24_2_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_24_2_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_25_2_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_25_2_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_25_3 (
    .io_in_r_data         (pe_mat_25_2_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_25_2_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_25_2_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_25_3_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_25_3_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_25_3_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_24_3_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_24_3_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_25_3_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_25_3_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_25_4 (
    .io_in_r_data         (pe_mat_25_3_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_25_3_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_25_3_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_25_4_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_25_4_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_25_4_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_24_4_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_24_4_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_25_4_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_25_4_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_25_5 (
    .io_in_r_data         (pe_mat_25_4_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_25_4_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_25_4_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_25_5_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_25_5_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_25_5_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_24_5_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_24_5_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_25_5_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_25_5_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_25_6 (
    .io_in_r_data         (pe_mat_25_5_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_25_5_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_25_5_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_25_6_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_25_6_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_25_6_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_24_6_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_24_6_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_25_6_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_25_6_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_25_7 (
    .io_in_r_data         (pe_mat_25_6_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_25_6_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_25_6_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_25_7_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_25_7_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_25_7_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_24_7_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_24_7_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_25_7_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_25_7_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_25_8 (
    .io_in_r_data         (pe_mat_25_7_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_25_7_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_25_7_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_25_8_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_25_8_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_25_8_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_24_8_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_24_8_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_25_8_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_25_8_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_25_9 (
    .io_in_r_data         (pe_mat_25_8_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_25_8_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_25_8_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_25_9_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_25_9_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_25_9_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_24_9_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_24_9_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_25_9_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_25_9_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_25_10 (
    .io_in_r_data         (pe_mat_25_9_io_out_r_data[15:0]  ), //i
    .io_in_r_stop_weight  (pe_mat_25_9_io_out_r_stop_weight ), //i
    .io_in_r_stall        (pe_mat_25_9_io_out_r_stall       ), //i
    .io_out_r_data        (pe_mat_25_10_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_25_10_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_25_10_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_24_10_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_24_10_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_25_10_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_25_10_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_25_11 (
    .io_in_r_data         (pe_mat_25_10_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_25_10_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_25_10_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_25_11_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_25_11_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_25_11_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_24_11_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_24_11_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_25_11_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_25_11_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_25_12 (
    .io_in_r_data         (pe_mat_25_11_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_25_11_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_25_11_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_25_12_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_25_12_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_25_12_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_24_12_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_24_12_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_25_12_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_25_12_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_25_13 (
    .io_in_r_data         (pe_mat_25_12_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_25_12_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_25_12_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_25_13_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_25_13_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_25_13_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_24_13_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_24_13_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_25_13_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_25_13_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_25_14 (
    .io_in_r_data         (pe_mat_25_13_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_25_13_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_25_13_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_25_14_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_25_14_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_25_14_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_24_14_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_24_14_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_25_14_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_25_14_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_25_15 (
    .io_in_r_data         (pe_mat_25_14_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_25_14_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_25_14_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_25_15_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_25_15_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_25_15_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_24_15_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_24_15_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_25_15_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_25_15_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_25_16 (
    .io_in_r_data         (pe_mat_25_15_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_25_15_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_25_15_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_25_16_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_25_16_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_25_16_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_24_16_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_24_16_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_25_16_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_25_16_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_25_17 (
    .io_in_r_data         (pe_mat_25_16_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_25_16_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_25_16_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_25_17_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_25_17_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_25_17_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_24_17_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_24_17_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_25_17_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_25_17_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_25_18 (
    .io_in_r_data         (pe_mat_25_17_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_25_17_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_25_17_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_25_18_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_25_18_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_25_18_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_24_18_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_24_18_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_25_18_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_25_18_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_25_19 (
    .io_in_r_data         (pe_mat_25_18_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_25_18_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_25_18_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_25_19_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_25_19_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_25_19_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_24_19_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_24_19_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_25_19_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_25_19_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_25_20 (
    .io_in_r_data         (pe_mat_25_19_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_25_19_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_25_19_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_25_20_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_25_20_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_25_20_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_24_20_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_24_20_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_25_20_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_25_20_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_25_21 (
    .io_in_r_data         (pe_mat_25_20_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_25_20_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_25_20_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_25_21_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_25_21_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_25_21_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_24_21_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_24_21_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_25_21_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_25_21_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_25_22 (
    .io_in_r_data         (pe_mat_25_21_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_25_21_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_25_21_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_25_22_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_25_22_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_25_22_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_24_22_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_24_22_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_25_22_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_25_22_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_25_23 (
    .io_in_r_data         (pe_mat_25_22_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_25_22_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_25_22_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_25_23_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_25_23_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_25_23_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_24_23_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_24_23_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_25_23_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_25_23_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_25_24 (
    .io_in_r_data         (pe_mat_25_23_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_25_23_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_25_23_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_25_24_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_25_24_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_25_24_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_24_24_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_24_24_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_25_24_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_25_24_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_25_25 (
    .io_in_r_data         (pe_mat_25_24_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_25_24_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_25_24_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_25_25_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_25_25_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_25_25_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_24_25_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_24_25_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_25_25_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_25_25_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_25_26 (
    .io_in_r_data         (pe_mat_25_25_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_25_25_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_25_25_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_25_26_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_25_26_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_25_26_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_24_26_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_24_26_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_25_26_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_25_26_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_25_27 (
    .io_in_r_data         (pe_mat_25_26_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_25_26_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_25_26_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_25_27_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_25_27_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_25_27_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_24_27_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_24_27_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_25_27_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_25_27_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_25_28 (
    .io_in_r_data         (pe_mat_25_27_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_25_27_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_25_27_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_25_28_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_25_28_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_25_28_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_24_28_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_24_28_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_25_28_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_25_28_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_25_29 (
    .io_in_r_data         (pe_mat_25_28_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_25_28_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_25_28_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_25_29_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_25_29_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_25_29_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_24_29_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_24_29_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_25_29_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_25_29_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_25_30 (
    .io_in_r_data         (pe_mat_25_29_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_25_29_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_25_29_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_25_30_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_25_30_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_25_30_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_24_30_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_24_30_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_25_30_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_25_30_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_25_31 (
    .io_in_r_data         (pe_mat_25_30_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_25_30_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_25_30_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_25_31_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_25_31_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_25_31_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_24_31_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_24_31_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_25_31_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_25_31_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_26_0 (
    .io_in_r_data         (io_in_r_26_data[15:0]           ), //i
    .io_in_r_stop_weight  (io_in_r_26_stop_weight          ), //i
    .io_in_r_stall        (io_in_r_26_stall                ), //i
    .io_out_r_data        (pe_mat_26_0_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_26_0_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_26_0_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_25_0_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_25_0_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_26_0_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_26_0_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_26_1 (
    .io_in_r_data         (pe_mat_26_0_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_26_0_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_26_0_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_26_1_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_26_1_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_26_1_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_25_1_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_25_1_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_26_1_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_26_1_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_26_2 (
    .io_in_r_data         (pe_mat_26_1_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_26_1_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_26_1_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_26_2_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_26_2_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_26_2_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_25_2_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_25_2_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_26_2_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_26_2_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_26_3 (
    .io_in_r_data         (pe_mat_26_2_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_26_2_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_26_2_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_26_3_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_26_3_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_26_3_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_25_3_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_25_3_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_26_3_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_26_3_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_26_4 (
    .io_in_r_data         (pe_mat_26_3_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_26_3_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_26_3_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_26_4_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_26_4_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_26_4_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_25_4_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_25_4_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_26_4_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_26_4_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_26_5 (
    .io_in_r_data         (pe_mat_26_4_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_26_4_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_26_4_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_26_5_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_26_5_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_26_5_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_25_5_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_25_5_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_26_5_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_26_5_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_26_6 (
    .io_in_r_data         (pe_mat_26_5_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_26_5_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_26_5_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_26_6_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_26_6_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_26_6_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_25_6_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_25_6_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_26_6_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_26_6_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_26_7 (
    .io_in_r_data         (pe_mat_26_6_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_26_6_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_26_6_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_26_7_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_26_7_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_26_7_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_25_7_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_25_7_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_26_7_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_26_7_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_26_8 (
    .io_in_r_data         (pe_mat_26_7_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_26_7_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_26_7_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_26_8_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_26_8_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_26_8_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_25_8_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_25_8_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_26_8_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_26_8_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_26_9 (
    .io_in_r_data         (pe_mat_26_8_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_26_8_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_26_8_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_26_9_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_26_9_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_26_9_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_25_9_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_25_9_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_26_9_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_26_9_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_26_10 (
    .io_in_r_data         (pe_mat_26_9_io_out_r_data[15:0]  ), //i
    .io_in_r_stop_weight  (pe_mat_26_9_io_out_r_stop_weight ), //i
    .io_in_r_stall        (pe_mat_26_9_io_out_r_stall       ), //i
    .io_out_r_data        (pe_mat_26_10_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_26_10_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_26_10_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_25_10_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_25_10_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_26_10_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_26_10_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_26_11 (
    .io_in_r_data         (pe_mat_26_10_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_26_10_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_26_10_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_26_11_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_26_11_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_26_11_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_25_11_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_25_11_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_26_11_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_26_11_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_26_12 (
    .io_in_r_data         (pe_mat_26_11_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_26_11_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_26_11_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_26_12_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_26_12_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_26_12_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_25_12_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_25_12_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_26_12_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_26_12_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_26_13 (
    .io_in_r_data         (pe_mat_26_12_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_26_12_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_26_12_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_26_13_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_26_13_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_26_13_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_25_13_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_25_13_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_26_13_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_26_13_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_26_14 (
    .io_in_r_data         (pe_mat_26_13_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_26_13_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_26_13_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_26_14_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_26_14_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_26_14_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_25_14_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_25_14_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_26_14_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_26_14_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_26_15 (
    .io_in_r_data         (pe_mat_26_14_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_26_14_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_26_14_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_26_15_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_26_15_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_26_15_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_25_15_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_25_15_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_26_15_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_26_15_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_26_16 (
    .io_in_r_data         (pe_mat_26_15_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_26_15_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_26_15_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_26_16_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_26_16_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_26_16_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_25_16_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_25_16_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_26_16_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_26_16_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_26_17 (
    .io_in_r_data         (pe_mat_26_16_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_26_16_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_26_16_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_26_17_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_26_17_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_26_17_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_25_17_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_25_17_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_26_17_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_26_17_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_26_18 (
    .io_in_r_data         (pe_mat_26_17_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_26_17_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_26_17_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_26_18_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_26_18_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_26_18_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_25_18_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_25_18_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_26_18_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_26_18_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_26_19 (
    .io_in_r_data         (pe_mat_26_18_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_26_18_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_26_18_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_26_19_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_26_19_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_26_19_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_25_19_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_25_19_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_26_19_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_26_19_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_26_20 (
    .io_in_r_data         (pe_mat_26_19_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_26_19_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_26_19_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_26_20_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_26_20_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_26_20_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_25_20_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_25_20_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_26_20_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_26_20_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_26_21 (
    .io_in_r_data         (pe_mat_26_20_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_26_20_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_26_20_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_26_21_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_26_21_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_26_21_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_25_21_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_25_21_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_26_21_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_26_21_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_26_22 (
    .io_in_r_data         (pe_mat_26_21_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_26_21_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_26_21_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_26_22_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_26_22_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_26_22_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_25_22_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_25_22_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_26_22_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_26_22_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_26_23 (
    .io_in_r_data         (pe_mat_26_22_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_26_22_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_26_22_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_26_23_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_26_23_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_26_23_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_25_23_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_25_23_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_26_23_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_26_23_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_26_24 (
    .io_in_r_data         (pe_mat_26_23_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_26_23_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_26_23_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_26_24_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_26_24_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_26_24_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_25_24_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_25_24_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_26_24_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_26_24_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_26_25 (
    .io_in_r_data         (pe_mat_26_24_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_26_24_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_26_24_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_26_25_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_26_25_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_26_25_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_25_25_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_25_25_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_26_25_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_26_25_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_26_26 (
    .io_in_r_data         (pe_mat_26_25_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_26_25_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_26_25_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_26_26_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_26_26_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_26_26_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_25_26_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_25_26_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_26_26_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_26_26_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_26_27 (
    .io_in_r_data         (pe_mat_26_26_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_26_26_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_26_26_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_26_27_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_26_27_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_26_27_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_25_27_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_25_27_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_26_27_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_26_27_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_26_28 (
    .io_in_r_data         (pe_mat_26_27_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_26_27_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_26_27_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_26_28_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_26_28_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_26_28_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_25_28_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_25_28_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_26_28_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_26_28_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_26_29 (
    .io_in_r_data         (pe_mat_26_28_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_26_28_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_26_28_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_26_29_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_26_29_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_26_29_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_25_29_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_25_29_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_26_29_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_26_29_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_26_30 (
    .io_in_r_data         (pe_mat_26_29_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_26_29_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_26_29_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_26_30_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_26_30_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_26_30_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_25_30_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_25_30_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_26_30_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_26_30_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_26_31 (
    .io_in_r_data         (pe_mat_26_30_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_26_30_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_26_30_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_26_31_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_26_31_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_26_31_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_25_31_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_25_31_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_26_31_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_26_31_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_27_0 (
    .io_in_r_data         (io_in_r_27_data[15:0]           ), //i
    .io_in_r_stop_weight  (io_in_r_27_stop_weight          ), //i
    .io_in_r_stall        (io_in_r_27_stall                ), //i
    .io_out_r_data        (pe_mat_27_0_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_27_0_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_27_0_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_26_0_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_26_0_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_27_0_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_27_0_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_27_1 (
    .io_in_r_data         (pe_mat_27_0_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_27_0_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_27_0_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_27_1_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_27_1_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_27_1_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_26_1_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_26_1_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_27_1_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_27_1_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_27_2 (
    .io_in_r_data         (pe_mat_27_1_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_27_1_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_27_1_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_27_2_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_27_2_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_27_2_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_26_2_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_26_2_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_27_2_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_27_2_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_27_3 (
    .io_in_r_data         (pe_mat_27_2_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_27_2_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_27_2_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_27_3_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_27_3_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_27_3_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_26_3_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_26_3_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_27_3_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_27_3_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_27_4 (
    .io_in_r_data         (pe_mat_27_3_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_27_3_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_27_3_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_27_4_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_27_4_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_27_4_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_26_4_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_26_4_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_27_4_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_27_4_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_27_5 (
    .io_in_r_data         (pe_mat_27_4_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_27_4_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_27_4_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_27_5_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_27_5_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_27_5_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_26_5_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_26_5_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_27_5_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_27_5_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_27_6 (
    .io_in_r_data         (pe_mat_27_5_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_27_5_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_27_5_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_27_6_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_27_6_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_27_6_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_26_6_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_26_6_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_27_6_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_27_6_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_27_7 (
    .io_in_r_data         (pe_mat_27_6_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_27_6_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_27_6_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_27_7_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_27_7_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_27_7_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_26_7_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_26_7_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_27_7_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_27_7_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_27_8 (
    .io_in_r_data         (pe_mat_27_7_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_27_7_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_27_7_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_27_8_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_27_8_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_27_8_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_26_8_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_26_8_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_27_8_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_27_8_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_27_9 (
    .io_in_r_data         (pe_mat_27_8_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_27_8_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_27_8_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_27_9_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_27_9_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_27_9_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_26_9_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_26_9_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_27_9_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_27_9_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_27_10 (
    .io_in_r_data         (pe_mat_27_9_io_out_r_data[15:0]  ), //i
    .io_in_r_stop_weight  (pe_mat_27_9_io_out_r_stop_weight ), //i
    .io_in_r_stall        (pe_mat_27_9_io_out_r_stall       ), //i
    .io_out_r_data        (pe_mat_27_10_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_27_10_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_27_10_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_26_10_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_26_10_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_27_10_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_27_10_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_27_11 (
    .io_in_r_data         (pe_mat_27_10_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_27_10_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_27_10_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_27_11_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_27_11_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_27_11_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_26_11_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_26_11_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_27_11_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_27_11_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_27_12 (
    .io_in_r_data         (pe_mat_27_11_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_27_11_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_27_11_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_27_12_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_27_12_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_27_12_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_26_12_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_26_12_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_27_12_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_27_12_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_27_13 (
    .io_in_r_data         (pe_mat_27_12_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_27_12_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_27_12_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_27_13_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_27_13_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_27_13_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_26_13_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_26_13_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_27_13_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_27_13_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_27_14 (
    .io_in_r_data         (pe_mat_27_13_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_27_13_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_27_13_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_27_14_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_27_14_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_27_14_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_26_14_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_26_14_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_27_14_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_27_14_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_27_15 (
    .io_in_r_data         (pe_mat_27_14_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_27_14_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_27_14_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_27_15_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_27_15_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_27_15_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_26_15_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_26_15_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_27_15_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_27_15_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_27_16 (
    .io_in_r_data         (pe_mat_27_15_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_27_15_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_27_15_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_27_16_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_27_16_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_27_16_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_26_16_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_26_16_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_27_16_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_27_16_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_27_17 (
    .io_in_r_data         (pe_mat_27_16_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_27_16_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_27_16_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_27_17_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_27_17_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_27_17_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_26_17_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_26_17_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_27_17_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_27_17_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_27_18 (
    .io_in_r_data         (pe_mat_27_17_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_27_17_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_27_17_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_27_18_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_27_18_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_27_18_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_26_18_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_26_18_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_27_18_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_27_18_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_27_19 (
    .io_in_r_data         (pe_mat_27_18_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_27_18_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_27_18_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_27_19_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_27_19_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_27_19_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_26_19_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_26_19_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_27_19_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_27_19_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_27_20 (
    .io_in_r_data         (pe_mat_27_19_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_27_19_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_27_19_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_27_20_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_27_20_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_27_20_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_26_20_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_26_20_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_27_20_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_27_20_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_27_21 (
    .io_in_r_data         (pe_mat_27_20_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_27_20_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_27_20_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_27_21_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_27_21_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_27_21_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_26_21_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_26_21_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_27_21_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_27_21_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_27_22 (
    .io_in_r_data         (pe_mat_27_21_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_27_21_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_27_21_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_27_22_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_27_22_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_27_22_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_26_22_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_26_22_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_27_22_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_27_22_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_27_23 (
    .io_in_r_data         (pe_mat_27_22_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_27_22_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_27_22_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_27_23_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_27_23_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_27_23_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_26_23_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_26_23_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_27_23_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_27_23_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_27_24 (
    .io_in_r_data         (pe_mat_27_23_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_27_23_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_27_23_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_27_24_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_27_24_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_27_24_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_26_24_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_26_24_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_27_24_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_27_24_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_27_25 (
    .io_in_r_data         (pe_mat_27_24_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_27_24_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_27_24_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_27_25_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_27_25_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_27_25_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_26_25_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_26_25_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_27_25_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_27_25_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_27_26 (
    .io_in_r_data         (pe_mat_27_25_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_27_25_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_27_25_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_27_26_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_27_26_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_27_26_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_26_26_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_26_26_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_27_26_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_27_26_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_27_27 (
    .io_in_r_data         (pe_mat_27_26_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_27_26_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_27_26_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_27_27_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_27_27_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_27_27_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_26_27_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_26_27_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_27_27_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_27_27_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_27_28 (
    .io_in_r_data         (pe_mat_27_27_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_27_27_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_27_27_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_27_28_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_27_28_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_27_28_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_26_28_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_26_28_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_27_28_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_27_28_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_27_29 (
    .io_in_r_data         (pe_mat_27_28_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_27_28_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_27_28_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_27_29_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_27_29_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_27_29_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_26_29_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_26_29_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_27_29_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_27_29_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_27_30 (
    .io_in_r_data         (pe_mat_27_29_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_27_29_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_27_29_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_27_30_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_27_30_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_27_30_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_26_30_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_26_30_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_27_30_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_27_30_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_27_31 (
    .io_in_r_data         (pe_mat_27_30_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_27_30_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_27_30_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_27_31_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_27_31_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_27_31_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_26_31_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_26_31_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_27_31_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_27_31_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_28_0 (
    .io_in_r_data         (io_in_r_28_data[15:0]           ), //i
    .io_in_r_stop_weight  (io_in_r_28_stop_weight          ), //i
    .io_in_r_stall        (io_in_r_28_stall                ), //i
    .io_out_r_data        (pe_mat_28_0_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_28_0_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_28_0_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_27_0_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_27_0_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_28_0_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_28_0_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_28_1 (
    .io_in_r_data         (pe_mat_28_0_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_28_0_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_28_0_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_28_1_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_28_1_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_28_1_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_27_1_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_27_1_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_28_1_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_28_1_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_28_2 (
    .io_in_r_data         (pe_mat_28_1_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_28_1_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_28_1_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_28_2_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_28_2_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_28_2_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_27_2_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_27_2_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_28_2_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_28_2_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_28_3 (
    .io_in_r_data         (pe_mat_28_2_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_28_2_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_28_2_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_28_3_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_28_3_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_28_3_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_27_3_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_27_3_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_28_3_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_28_3_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_28_4 (
    .io_in_r_data         (pe_mat_28_3_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_28_3_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_28_3_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_28_4_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_28_4_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_28_4_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_27_4_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_27_4_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_28_4_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_28_4_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_28_5 (
    .io_in_r_data         (pe_mat_28_4_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_28_4_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_28_4_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_28_5_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_28_5_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_28_5_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_27_5_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_27_5_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_28_5_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_28_5_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_28_6 (
    .io_in_r_data         (pe_mat_28_5_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_28_5_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_28_5_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_28_6_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_28_6_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_28_6_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_27_6_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_27_6_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_28_6_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_28_6_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_28_7 (
    .io_in_r_data         (pe_mat_28_6_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_28_6_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_28_6_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_28_7_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_28_7_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_28_7_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_27_7_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_27_7_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_28_7_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_28_7_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_28_8 (
    .io_in_r_data         (pe_mat_28_7_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_28_7_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_28_7_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_28_8_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_28_8_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_28_8_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_27_8_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_27_8_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_28_8_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_28_8_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_28_9 (
    .io_in_r_data         (pe_mat_28_8_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_28_8_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_28_8_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_28_9_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_28_9_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_28_9_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_27_9_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_27_9_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_28_9_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_28_9_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_28_10 (
    .io_in_r_data         (pe_mat_28_9_io_out_r_data[15:0]  ), //i
    .io_in_r_stop_weight  (pe_mat_28_9_io_out_r_stop_weight ), //i
    .io_in_r_stall        (pe_mat_28_9_io_out_r_stall       ), //i
    .io_out_r_data        (pe_mat_28_10_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_28_10_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_28_10_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_27_10_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_27_10_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_28_10_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_28_10_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_28_11 (
    .io_in_r_data         (pe_mat_28_10_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_28_10_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_28_10_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_28_11_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_28_11_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_28_11_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_27_11_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_27_11_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_28_11_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_28_11_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_28_12 (
    .io_in_r_data         (pe_mat_28_11_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_28_11_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_28_11_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_28_12_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_28_12_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_28_12_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_27_12_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_27_12_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_28_12_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_28_12_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_28_13 (
    .io_in_r_data         (pe_mat_28_12_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_28_12_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_28_12_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_28_13_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_28_13_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_28_13_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_27_13_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_27_13_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_28_13_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_28_13_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_28_14 (
    .io_in_r_data         (pe_mat_28_13_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_28_13_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_28_13_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_28_14_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_28_14_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_28_14_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_27_14_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_27_14_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_28_14_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_28_14_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_28_15 (
    .io_in_r_data         (pe_mat_28_14_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_28_14_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_28_14_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_28_15_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_28_15_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_28_15_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_27_15_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_27_15_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_28_15_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_28_15_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_28_16 (
    .io_in_r_data         (pe_mat_28_15_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_28_15_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_28_15_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_28_16_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_28_16_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_28_16_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_27_16_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_27_16_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_28_16_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_28_16_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_28_17 (
    .io_in_r_data         (pe_mat_28_16_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_28_16_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_28_16_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_28_17_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_28_17_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_28_17_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_27_17_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_27_17_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_28_17_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_28_17_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_28_18 (
    .io_in_r_data         (pe_mat_28_17_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_28_17_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_28_17_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_28_18_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_28_18_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_28_18_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_27_18_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_27_18_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_28_18_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_28_18_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_28_19 (
    .io_in_r_data         (pe_mat_28_18_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_28_18_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_28_18_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_28_19_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_28_19_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_28_19_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_27_19_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_27_19_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_28_19_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_28_19_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_28_20 (
    .io_in_r_data         (pe_mat_28_19_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_28_19_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_28_19_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_28_20_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_28_20_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_28_20_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_27_20_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_27_20_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_28_20_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_28_20_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_28_21 (
    .io_in_r_data         (pe_mat_28_20_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_28_20_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_28_20_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_28_21_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_28_21_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_28_21_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_27_21_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_27_21_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_28_21_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_28_21_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_28_22 (
    .io_in_r_data         (pe_mat_28_21_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_28_21_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_28_21_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_28_22_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_28_22_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_28_22_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_27_22_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_27_22_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_28_22_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_28_22_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_28_23 (
    .io_in_r_data         (pe_mat_28_22_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_28_22_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_28_22_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_28_23_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_28_23_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_28_23_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_27_23_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_27_23_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_28_23_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_28_23_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_28_24 (
    .io_in_r_data         (pe_mat_28_23_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_28_23_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_28_23_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_28_24_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_28_24_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_28_24_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_27_24_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_27_24_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_28_24_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_28_24_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_28_25 (
    .io_in_r_data         (pe_mat_28_24_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_28_24_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_28_24_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_28_25_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_28_25_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_28_25_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_27_25_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_27_25_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_28_25_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_28_25_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_28_26 (
    .io_in_r_data         (pe_mat_28_25_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_28_25_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_28_25_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_28_26_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_28_26_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_28_26_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_27_26_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_27_26_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_28_26_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_28_26_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_28_27 (
    .io_in_r_data         (pe_mat_28_26_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_28_26_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_28_26_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_28_27_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_28_27_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_28_27_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_27_27_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_27_27_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_28_27_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_28_27_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_28_28 (
    .io_in_r_data         (pe_mat_28_27_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_28_27_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_28_27_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_28_28_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_28_28_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_28_28_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_27_28_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_27_28_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_28_28_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_28_28_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_28_29 (
    .io_in_r_data         (pe_mat_28_28_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_28_28_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_28_28_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_28_29_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_28_29_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_28_29_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_27_29_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_27_29_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_28_29_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_28_29_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_28_30 (
    .io_in_r_data         (pe_mat_28_29_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_28_29_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_28_29_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_28_30_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_28_30_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_28_30_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_27_30_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_27_30_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_28_30_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_28_30_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_28_31 (
    .io_in_r_data         (pe_mat_28_30_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_28_30_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_28_30_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_28_31_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_28_31_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_28_31_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_27_31_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_27_31_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_28_31_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_28_31_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_29_0 (
    .io_in_r_data         (io_in_r_29_data[15:0]           ), //i
    .io_in_r_stop_weight  (io_in_r_29_stop_weight          ), //i
    .io_in_r_stall        (io_in_r_29_stall                ), //i
    .io_out_r_data        (pe_mat_29_0_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_29_0_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_29_0_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_28_0_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_28_0_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_29_0_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_29_0_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_29_1 (
    .io_in_r_data         (pe_mat_29_0_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_29_0_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_29_0_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_29_1_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_29_1_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_29_1_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_28_1_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_28_1_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_29_1_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_29_1_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_29_2 (
    .io_in_r_data         (pe_mat_29_1_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_29_1_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_29_1_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_29_2_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_29_2_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_29_2_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_28_2_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_28_2_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_29_2_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_29_2_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_29_3 (
    .io_in_r_data         (pe_mat_29_2_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_29_2_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_29_2_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_29_3_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_29_3_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_29_3_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_28_3_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_28_3_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_29_3_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_29_3_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_29_4 (
    .io_in_r_data         (pe_mat_29_3_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_29_3_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_29_3_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_29_4_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_29_4_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_29_4_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_28_4_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_28_4_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_29_4_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_29_4_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_29_5 (
    .io_in_r_data         (pe_mat_29_4_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_29_4_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_29_4_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_29_5_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_29_5_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_29_5_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_28_5_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_28_5_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_29_5_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_29_5_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_29_6 (
    .io_in_r_data         (pe_mat_29_5_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_29_5_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_29_5_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_29_6_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_29_6_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_29_6_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_28_6_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_28_6_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_29_6_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_29_6_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_29_7 (
    .io_in_r_data         (pe_mat_29_6_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_29_6_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_29_6_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_29_7_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_29_7_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_29_7_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_28_7_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_28_7_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_29_7_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_29_7_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_29_8 (
    .io_in_r_data         (pe_mat_29_7_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_29_7_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_29_7_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_29_8_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_29_8_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_29_8_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_28_8_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_28_8_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_29_8_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_29_8_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_29_9 (
    .io_in_r_data         (pe_mat_29_8_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_29_8_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_29_8_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_29_9_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_29_9_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_29_9_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_28_9_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_28_9_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_29_9_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_29_9_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_29_10 (
    .io_in_r_data         (pe_mat_29_9_io_out_r_data[15:0]  ), //i
    .io_in_r_stop_weight  (pe_mat_29_9_io_out_r_stop_weight ), //i
    .io_in_r_stall        (pe_mat_29_9_io_out_r_stall       ), //i
    .io_out_r_data        (pe_mat_29_10_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_29_10_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_29_10_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_28_10_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_28_10_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_29_10_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_29_10_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_29_11 (
    .io_in_r_data         (pe_mat_29_10_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_29_10_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_29_10_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_29_11_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_29_11_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_29_11_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_28_11_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_28_11_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_29_11_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_29_11_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_29_12 (
    .io_in_r_data         (pe_mat_29_11_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_29_11_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_29_11_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_29_12_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_29_12_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_29_12_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_28_12_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_28_12_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_29_12_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_29_12_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_29_13 (
    .io_in_r_data         (pe_mat_29_12_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_29_12_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_29_12_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_29_13_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_29_13_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_29_13_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_28_13_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_28_13_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_29_13_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_29_13_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_29_14 (
    .io_in_r_data         (pe_mat_29_13_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_29_13_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_29_13_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_29_14_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_29_14_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_29_14_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_28_14_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_28_14_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_29_14_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_29_14_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_29_15 (
    .io_in_r_data         (pe_mat_29_14_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_29_14_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_29_14_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_29_15_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_29_15_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_29_15_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_28_15_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_28_15_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_29_15_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_29_15_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_29_16 (
    .io_in_r_data         (pe_mat_29_15_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_29_15_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_29_15_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_29_16_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_29_16_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_29_16_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_28_16_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_28_16_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_29_16_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_29_16_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_29_17 (
    .io_in_r_data         (pe_mat_29_16_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_29_16_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_29_16_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_29_17_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_29_17_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_29_17_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_28_17_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_28_17_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_29_17_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_29_17_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_29_18 (
    .io_in_r_data         (pe_mat_29_17_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_29_17_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_29_17_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_29_18_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_29_18_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_29_18_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_28_18_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_28_18_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_29_18_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_29_18_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_29_19 (
    .io_in_r_data         (pe_mat_29_18_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_29_18_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_29_18_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_29_19_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_29_19_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_29_19_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_28_19_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_28_19_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_29_19_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_29_19_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_29_20 (
    .io_in_r_data         (pe_mat_29_19_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_29_19_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_29_19_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_29_20_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_29_20_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_29_20_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_28_20_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_28_20_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_29_20_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_29_20_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_29_21 (
    .io_in_r_data         (pe_mat_29_20_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_29_20_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_29_20_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_29_21_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_29_21_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_29_21_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_28_21_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_28_21_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_29_21_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_29_21_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_29_22 (
    .io_in_r_data         (pe_mat_29_21_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_29_21_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_29_21_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_29_22_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_29_22_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_29_22_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_28_22_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_28_22_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_29_22_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_29_22_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_29_23 (
    .io_in_r_data         (pe_mat_29_22_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_29_22_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_29_22_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_29_23_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_29_23_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_29_23_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_28_23_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_28_23_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_29_23_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_29_23_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_29_24 (
    .io_in_r_data         (pe_mat_29_23_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_29_23_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_29_23_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_29_24_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_29_24_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_29_24_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_28_24_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_28_24_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_29_24_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_29_24_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_29_25 (
    .io_in_r_data         (pe_mat_29_24_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_29_24_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_29_24_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_29_25_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_29_25_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_29_25_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_28_25_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_28_25_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_29_25_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_29_25_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_29_26 (
    .io_in_r_data         (pe_mat_29_25_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_29_25_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_29_25_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_29_26_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_29_26_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_29_26_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_28_26_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_28_26_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_29_26_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_29_26_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_29_27 (
    .io_in_r_data         (pe_mat_29_26_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_29_26_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_29_26_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_29_27_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_29_27_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_29_27_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_28_27_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_28_27_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_29_27_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_29_27_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_29_28 (
    .io_in_r_data         (pe_mat_29_27_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_29_27_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_29_27_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_29_28_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_29_28_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_29_28_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_28_28_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_28_28_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_29_28_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_29_28_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_29_29 (
    .io_in_r_data         (pe_mat_29_28_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_29_28_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_29_28_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_29_29_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_29_29_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_29_29_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_28_29_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_28_29_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_29_29_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_29_29_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_29_30 (
    .io_in_r_data         (pe_mat_29_29_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_29_29_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_29_29_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_29_30_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_29_30_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_29_30_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_28_30_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_28_30_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_29_30_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_29_30_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_29_31 (
    .io_in_r_data         (pe_mat_29_30_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_29_30_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_29_30_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_29_31_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_29_31_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_29_31_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_28_31_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_28_31_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_29_31_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_29_31_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_30_0 (
    .io_in_r_data         (io_in_r_30_data[15:0]           ), //i
    .io_in_r_stop_weight  (io_in_r_30_stop_weight          ), //i
    .io_in_r_stall        (io_in_r_30_stall                ), //i
    .io_out_r_data        (pe_mat_30_0_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_30_0_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_30_0_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_29_0_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_29_0_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_30_0_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_30_0_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_30_1 (
    .io_in_r_data         (pe_mat_30_0_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_30_0_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_30_0_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_30_1_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_30_1_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_30_1_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_29_1_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_29_1_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_30_1_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_30_1_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_30_2 (
    .io_in_r_data         (pe_mat_30_1_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_30_1_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_30_1_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_30_2_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_30_2_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_30_2_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_29_2_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_29_2_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_30_2_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_30_2_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_30_3 (
    .io_in_r_data         (pe_mat_30_2_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_30_2_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_30_2_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_30_3_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_30_3_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_30_3_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_29_3_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_29_3_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_30_3_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_30_3_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_30_4 (
    .io_in_r_data         (pe_mat_30_3_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_30_3_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_30_3_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_30_4_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_30_4_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_30_4_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_29_4_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_29_4_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_30_4_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_30_4_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_30_5 (
    .io_in_r_data         (pe_mat_30_4_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_30_4_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_30_4_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_30_5_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_30_5_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_30_5_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_29_5_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_29_5_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_30_5_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_30_5_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_30_6 (
    .io_in_r_data         (pe_mat_30_5_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_30_5_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_30_5_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_30_6_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_30_6_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_30_6_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_29_6_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_29_6_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_30_6_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_30_6_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_30_7 (
    .io_in_r_data         (pe_mat_30_6_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_30_6_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_30_6_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_30_7_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_30_7_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_30_7_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_29_7_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_29_7_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_30_7_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_30_7_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_30_8 (
    .io_in_r_data         (pe_mat_30_7_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_30_7_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_30_7_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_30_8_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_30_8_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_30_8_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_29_8_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_29_8_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_30_8_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_30_8_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_30_9 (
    .io_in_r_data         (pe_mat_30_8_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_30_8_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_30_8_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_30_9_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_30_9_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_30_9_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_29_9_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_29_9_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_30_9_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_30_9_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_30_10 (
    .io_in_r_data         (pe_mat_30_9_io_out_r_data[15:0]  ), //i
    .io_in_r_stop_weight  (pe_mat_30_9_io_out_r_stop_weight ), //i
    .io_in_r_stall        (pe_mat_30_9_io_out_r_stall       ), //i
    .io_out_r_data        (pe_mat_30_10_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_30_10_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_30_10_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_29_10_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_29_10_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_30_10_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_30_10_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_30_11 (
    .io_in_r_data         (pe_mat_30_10_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_30_10_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_30_10_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_30_11_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_30_11_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_30_11_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_29_11_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_29_11_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_30_11_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_30_11_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_30_12 (
    .io_in_r_data         (pe_mat_30_11_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_30_11_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_30_11_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_30_12_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_30_12_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_30_12_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_29_12_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_29_12_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_30_12_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_30_12_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_30_13 (
    .io_in_r_data         (pe_mat_30_12_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_30_12_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_30_12_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_30_13_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_30_13_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_30_13_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_29_13_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_29_13_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_30_13_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_30_13_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_30_14 (
    .io_in_r_data         (pe_mat_30_13_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_30_13_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_30_13_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_30_14_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_30_14_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_30_14_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_29_14_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_29_14_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_30_14_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_30_14_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_30_15 (
    .io_in_r_data         (pe_mat_30_14_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_30_14_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_30_14_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_30_15_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_30_15_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_30_15_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_29_15_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_29_15_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_30_15_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_30_15_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_30_16 (
    .io_in_r_data         (pe_mat_30_15_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_30_15_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_30_15_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_30_16_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_30_16_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_30_16_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_29_16_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_29_16_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_30_16_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_30_16_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_30_17 (
    .io_in_r_data         (pe_mat_30_16_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_30_16_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_30_16_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_30_17_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_30_17_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_30_17_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_29_17_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_29_17_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_30_17_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_30_17_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_30_18 (
    .io_in_r_data         (pe_mat_30_17_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_30_17_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_30_17_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_30_18_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_30_18_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_30_18_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_29_18_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_29_18_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_30_18_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_30_18_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_30_19 (
    .io_in_r_data         (pe_mat_30_18_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_30_18_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_30_18_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_30_19_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_30_19_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_30_19_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_29_19_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_29_19_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_30_19_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_30_19_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_30_20 (
    .io_in_r_data         (pe_mat_30_19_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_30_19_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_30_19_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_30_20_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_30_20_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_30_20_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_29_20_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_29_20_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_30_20_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_30_20_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_30_21 (
    .io_in_r_data         (pe_mat_30_20_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_30_20_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_30_20_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_30_21_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_30_21_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_30_21_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_29_21_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_29_21_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_30_21_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_30_21_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_30_22 (
    .io_in_r_data         (pe_mat_30_21_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_30_21_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_30_21_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_30_22_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_30_22_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_30_22_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_29_22_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_29_22_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_30_22_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_30_22_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_30_23 (
    .io_in_r_data         (pe_mat_30_22_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_30_22_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_30_22_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_30_23_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_30_23_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_30_23_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_29_23_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_29_23_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_30_23_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_30_23_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_30_24 (
    .io_in_r_data         (pe_mat_30_23_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_30_23_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_30_23_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_30_24_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_30_24_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_30_24_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_29_24_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_29_24_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_30_24_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_30_24_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_30_25 (
    .io_in_r_data         (pe_mat_30_24_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_30_24_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_30_24_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_30_25_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_30_25_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_30_25_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_29_25_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_29_25_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_30_25_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_30_25_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_30_26 (
    .io_in_r_data         (pe_mat_30_25_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_30_25_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_30_25_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_30_26_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_30_26_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_30_26_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_29_26_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_29_26_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_30_26_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_30_26_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_30_27 (
    .io_in_r_data         (pe_mat_30_26_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_30_26_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_30_26_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_30_27_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_30_27_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_30_27_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_29_27_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_29_27_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_30_27_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_30_27_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_30_28 (
    .io_in_r_data         (pe_mat_30_27_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_30_27_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_30_27_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_30_28_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_30_28_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_30_28_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_29_28_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_29_28_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_30_28_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_30_28_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_30_29 (
    .io_in_r_data         (pe_mat_30_28_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_30_28_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_30_28_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_30_29_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_30_29_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_30_29_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_29_29_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_29_29_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_30_29_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_30_29_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_30_30 (
    .io_in_r_data         (pe_mat_30_29_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_30_29_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_30_29_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_30_30_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_30_30_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_30_30_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_29_30_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_29_30_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_30_30_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_30_30_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_30_31 (
    .io_in_r_data         (pe_mat_30_30_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_30_30_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_30_30_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_30_31_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_30_31_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_30_31_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_29_31_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_29_31_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_30_31_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_30_31_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_31_0 (
    .io_in_r_data         (io_in_r_31_data[15:0]           ), //i
    .io_in_r_stop_weight  (io_in_r_31_stop_weight          ), //i
    .io_in_r_stall        (io_in_r_31_stall                ), //i
    .io_out_r_data        (pe_mat_31_0_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_31_0_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_31_0_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_30_0_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_30_0_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_31_0_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_31_0_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_31_1 (
    .io_in_r_data         (pe_mat_31_0_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_31_0_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_31_0_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_31_1_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_31_1_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_31_1_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_30_1_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_30_1_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_31_1_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_31_1_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_31_2 (
    .io_in_r_data         (pe_mat_31_1_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_31_1_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_31_1_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_31_2_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_31_2_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_31_2_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_30_2_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_30_2_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_31_2_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_31_2_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_31_3 (
    .io_in_r_data         (pe_mat_31_2_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_31_2_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_31_2_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_31_3_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_31_3_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_31_3_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_30_3_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_30_3_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_31_3_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_31_3_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_31_4 (
    .io_in_r_data         (pe_mat_31_3_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_31_3_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_31_3_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_31_4_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_31_4_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_31_4_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_30_4_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_30_4_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_31_4_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_31_4_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_31_5 (
    .io_in_r_data         (pe_mat_31_4_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_31_4_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_31_4_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_31_5_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_31_5_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_31_5_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_30_5_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_30_5_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_31_5_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_31_5_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_31_6 (
    .io_in_r_data         (pe_mat_31_5_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_31_5_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_31_5_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_31_6_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_31_6_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_31_6_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_30_6_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_30_6_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_31_6_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_31_6_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_31_7 (
    .io_in_r_data         (pe_mat_31_6_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_31_6_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_31_6_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_31_7_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_31_7_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_31_7_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_30_7_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_30_7_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_31_7_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_31_7_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_31_8 (
    .io_in_r_data         (pe_mat_31_7_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_31_7_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_31_7_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_31_8_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_31_8_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_31_8_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_30_8_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_30_8_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_31_8_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_31_8_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_31_9 (
    .io_in_r_data         (pe_mat_31_8_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_31_8_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_31_8_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_31_9_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_31_9_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_31_9_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_30_9_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_30_9_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_31_9_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_31_9_io_out_c_is_weight  ), //o
    .clk                  (clk                             ), //i
    .reset                (reset                           )  //i
  );
  PEWS_1023 pe_mat_31_10 (
    .io_in_r_data         (pe_mat_31_9_io_out_r_data[15:0]  ), //i
    .io_in_r_stop_weight  (pe_mat_31_9_io_out_r_stop_weight ), //i
    .io_in_r_stall        (pe_mat_31_9_io_out_r_stall       ), //i
    .io_out_r_data        (pe_mat_31_10_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_31_10_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_31_10_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_30_10_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_30_10_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_31_10_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_31_10_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_31_11 (
    .io_in_r_data         (pe_mat_31_10_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_31_10_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_31_10_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_31_11_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_31_11_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_31_11_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_30_11_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_30_11_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_31_11_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_31_11_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_31_12 (
    .io_in_r_data         (pe_mat_31_11_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_31_11_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_31_11_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_31_12_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_31_12_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_31_12_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_30_12_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_30_12_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_31_12_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_31_12_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_31_13 (
    .io_in_r_data         (pe_mat_31_12_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_31_12_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_31_12_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_31_13_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_31_13_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_31_13_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_30_13_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_30_13_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_31_13_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_31_13_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_31_14 (
    .io_in_r_data         (pe_mat_31_13_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_31_13_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_31_13_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_31_14_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_31_14_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_31_14_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_30_14_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_30_14_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_31_14_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_31_14_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_31_15 (
    .io_in_r_data         (pe_mat_31_14_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_31_14_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_31_14_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_31_15_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_31_15_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_31_15_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_30_15_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_30_15_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_31_15_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_31_15_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_31_16 (
    .io_in_r_data         (pe_mat_31_15_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_31_15_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_31_15_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_31_16_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_31_16_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_31_16_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_30_16_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_30_16_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_31_16_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_31_16_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_31_17 (
    .io_in_r_data         (pe_mat_31_16_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_31_16_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_31_16_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_31_17_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_31_17_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_31_17_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_30_17_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_30_17_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_31_17_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_31_17_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_31_18 (
    .io_in_r_data         (pe_mat_31_17_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_31_17_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_31_17_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_31_18_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_31_18_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_31_18_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_30_18_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_30_18_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_31_18_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_31_18_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_31_19 (
    .io_in_r_data         (pe_mat_31_18_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_31_18_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_31_18_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_31_19_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_31_19_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_31_19_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_30_19_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_30_19_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_31_19_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_31_19_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_31_20 (
    .io_in_r_data         (pe_mat_31_19_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_31_19_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_31_19_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_31_20_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_31_20_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_31_20_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_30_20_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_30_20_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_31_20_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_31_20_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_31_21 (
    .io_in_r_data         (pe_mat_31_20_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_31_20_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_31_20_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_31_21_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_31_21_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_31_21_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_30_21_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_30_21_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_31_21_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_31_21_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_31_22 (
    .io_in_r_data         (pe_mat_31_21_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_31_21_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_31_21_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_31_22_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_31_22_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_31_22_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_30_22_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_30_22_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_31_22_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_31_22_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_31_23 (
    .io_in_r_data         (pe_mat_31_22_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_31_22_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_31_22_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_31_23_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_31_23_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_31_23_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_30_23_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_30_23_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_31_23_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_31_23_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_31_24 (
    .io_in_r_data         (pe_mat_31_23_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_31_23_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_31_23_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_31_24_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_31_24_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_31_24_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_30_24_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_30_24_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_31_24_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_31_24_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_31_25 (
    .io_in_r_data         (pe_mat_31_24_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_31_24_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_31_24_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_31_25_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_31_25_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_31_25_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_30_25_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_30_25_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_31_25_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_31_25_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_31_26 (
    .io_in_r_data         (pe_mat_31_25_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_31_25_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_31_25_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_31_26_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_31_26_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_31_26_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_30_26_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_30_26_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_31_26_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_31_26_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_31_27 (
    .io_in_r_data         (pe_mat_31_26_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_31_26_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_31_26_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_31_27_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_31_27_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_31_27_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_30_27_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_30_27_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_31_27_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_31_27_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_31_28 (
    .io_in_r_data         (pe_mat_31_27_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_31_27_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_31_27_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_31_28_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_31_28_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_31_28_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_30_28_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_30_28_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_31_28_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_31_28_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_31_29 (
    .io_in_r_data         (pe_mat_31_28_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_31_28_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_31_28_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_31_29_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_31_29_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_31_29_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_30_29_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_30_29_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_31_29_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_31_29_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_31_30 (
    .io_in_r_data         (pe_mat_31_29_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_31_29_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_31_29_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_31_30_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_31_30_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_31_30_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_30_30_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_30_30_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_31_30_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_31_30_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  PEWS_1023 pe_mat_31_31 (
    .io_in_r_data         (pe_mat_31_30_io_out_r_data[15:0] ), //i
    .io_in_r_stop_weight  (pe_mat_31_30_io_out_r_stop_weight), //i
    .io_in_r_stall        (pe_mat_31_30_io_out_r_stall      ), //i
    .io_out_r_data        (pe_mat_31_31_io_out_r_data[15:0] ), //o
    .io_out_r_stop_weight (pe_mat_31_31_io_out_r_stop_weight), //o
    .io_out_r_stall       (pe_mat_31_31_io_out_r_stall      ), //o
    .io_in_c_data         (pe_mat_30_31_io_out_c_data[15:0] ), //i
    .io_in_c_is_weight    (pe_mat_30_31_io_out_c_is_weight  ), //i
    .io_out_c_data        (pe_mat_31_31_io_out_c_data[15:0] ), //o
    .io_out_c_is_weight   (pe_mat_31_31_io_out_c_is_weight  ), //o
    .clk                  (clk                              ), //i
    .reset                (reset                            )  //i
  );
  assign io_out_r_0_data = pe_mat_0_31_io_out_r_data; // @[SystolicConnect.scala 50:16]
  assign io_out_r_0_stop_weight = pe_mat_0_31_io_out_r_stop_weight; // @[SystolicConnect.scala 50:16]
  assign io_out_r_0_stall = pe_mat_0_31_io_out_r_stall; // @[SystolicConnect.scala 50:16]
  assign io_out_r_1_data = pe_mat_1_31_io_out_r_data; // @[SystolicConnect.scala 50:16]
  assign io_out_r_1_stop_weight = pe_mat_1_31_io_out_r_stop_weight; // @[SystolicConnect.scala 50:16]
  assign io_out_r_1_stall = pe_mat_1_31_io_out_r_stall; // @[SystolicConnect.scala 50:16]
  assign io_out_r_2_data = pe_mat_2_31_io_out_r_data; // @[SystolicConnect.scala 50:16]
  assign io_out_r_2_stop_weight = pe_mat_2_31_io_out_r_stop_weight; // @[SystolicConnect.scala 50:16]
  assign io_out_r_2_stall = pe_mat_2_31_io_out_r_stall; // @[SystolicConnect.scala 50:16]
  assign io_out_r_3_data = pe_mat_3_31_io_out_r_data; // @[SystolicConnect.scala 50:16]
  assign io_out_r_3_stop_weight = pe_mat_3_31_io_out_r_stop_weight; // @[SystolicConnect.scala 50:16]
  assign io_out_r_3_stall = pe_mat_3_31_io_out_r_stall; // @[SystolicConnect.scala 50:16]
  assign io_out_r_4_data = pe_mat_4_31_io_out_r_data; // @[SystolicConnect.scala 50:16]
  assign io_out_r_4_stop_weight = pe_mat_4_31_io_out_r_stop_weight; // @[SystolicConnect.scala 50:16]
  assign io_out_r_4_stall = pe_mat_4_31_io_out_r_stall; // @[SystolicConnect.scala 50:16]
  assign io_out_r_5_data = pe_mat_5_31_io_out_r_data; // @[SystolicConnect.scala 50:16]
  assign io_out_r_5_stop_weight = pe_mat_5_31_io_out_r_stop_weight; // @[SystolicConnect.scala 50:16]
  assign io_out_r_5_stall = pe_mat_5_31_io_out_r_stall; // @[SystolicConnect.scala 50:16]
  assign io_out_r_6_data = pe_mat_6_31_io_out_r_data; // @[SystolicConnect.scala 50:16]
  assign io_out_r_6_stop_weight = pe_mat_6_31_io_out_r_stop_weight; // @[SystolicConnect.scala 50:16]
  assign io_out_r_6_stall = pe_mat_6_31_io_out_r_stall; // @[SystolicConnect.scala 50:16]
  assign io_out_r_7_data = pe_mat_7_31_io_out_r_data; // @[SystolicConnect.scala 50:16]
  assign io_out_r_7_stop_weight = pe_mat_7_31_io_out_r_stop_weight; // @[SystolicConnect.scala 50:16]
  assign io_out_r_7_stall = pe_mat_7_31_io_out_r_stall; // @[SystolicConnect.scala 50:16]
  assign io_out_r_8_data = pe_mat_8_31_io_out_r_data; // @[SystolicConnect.scala 50:16]
  assign io_out_r_8_stop_weight = pe_mat_8_31_io_out_r_stop_weight; // @[SystolicConnect.scala 50:16]
  assign io_out_r_8_stall = pe_mat_8_31_io_out_r_stall; // @[SystolicConnect.scala 50:16]
  assign io_out_r_9_data = pe_mat_9_31_io_out_r_data; // @[SystolicConnect.scala 50:16]
  assign io_out_r_9_stop_weight = pe_mat_9_31_io_out_r_stop_weight; // @[SystolicConnect.scala 50:16]
  assign io_out_r_9_stall = pe_mat_9_31_io_out_r_stall; // @[SystolicConnect.scala 50:16]
  assign io_out_r_10_data = pe_mat_10_31_io_out_r_data; // @[SystolicConnect.scala 50:16]
  assign io_out_r_10_stop_weight = pe_mat_10_31_io_out_r_stop_weight; // @[SystolicConnect.scala 50:16]
  assign io_out_r_10_stall = pe_mat_10_31_io_out_r_stall; // @[SystolicConnect.scala 50:16]
  assign io_out_r_11_data = pe_mat_11_31_io_out_r_data; // @[SystolicConnect.scala 50:16]
  assign io_out_r_11_stop_weight = pe_mat_11_31_io_out_r_stop_weight; // @[SystolicConnect.scala 50:16]
  assign io_out_r_11_stall = pe_mat_11_31_io_out_r_stall; // @[SystolicConnect.scala 50:16]
  assign io_out_r_12_data = pe_mat_12_31_io_out_r_data; // @[SystolicConnect.scala 50:16]
  assign io_out_r_12_stop_weight = pe_mat_12_31_io_out_r_stop_weight; // @[SystolicConnect.scala 50:16]
  assign io_out_r_12_stall = pe_mat_12_31_io_out_r_stall; // @[SystolicConnect.scala 50:16]
  assign io_out_r_13_data = pe_mat_13_31_io_out_r_data; // @[SystolicConnect.scala 50:16]
  assign io_out_r_13_stop_weight = pe_mat_13_31_io_out_r_stop_weight; // @[SystolicConnect.scala 50:16]
  assign io_out_r_13_stall = pe_mat_13_31_io_out_r_stall; // @[SystolicConnect.scala 50:16]
  assign io_out_r_14_data = pe_mat_14_31_io_out_r_data; // @[SystolicConnect.scala 50:16]
  assign io_out_r_14_stop_weight = pe_mat_14_31_io_out_r_stop_weight; // @[SystolicConnect.scala 50:16]
  assign io_out_r_14_stall = pe_mat_14_31_io_out_r_stall; // @[SystolicConnect.scala 50:16]
  assign io_out_r_15_data = pe_mat_15_31_io_out_r_data; // @[SystolicConnect.scala 50:16]
  assign io_out_r_15_stop_weight = pe_mat_15_31_io_out_r_stop_weight; // @[SystolicConnect.scala 50:16]
  assign io_out_r_15_stall = pe_mat_15_31_io_out_r_stall; // @[SystolicConnect.scala 50:16]
  assign io_out_r_16_data = pe_mat_16_31_io_out_r_data; // @[SystolicConnect.scala 50:16]
  assign io_out_r_16_stop_weight = pe_mat_16_31_io_out_r_stop_weight; // @[SystolicConnect.scala 50:16]
  assign io_out_r_16_stall = pe_mat_16_31_io_out_r_stall; // @[SystolicConnect.scala 50:16]
  assign io_out_r_17_data = pe_mat_17_31_io_out_r_data; // @[SystolicConnect.scala 50:16]
  assign io_out_r_17_stop_weight = pe_mat_17_31_io_out_r_stop_weight; // @[SystolicConnect.scala 50:16]
  assign io_out_r_17_stall = pe_mat_17_31_io_out_r_stall; // @[SystolicConnect.scala 50:16]
  assign io_out_r_18_data = pe_mat_18_31_io_out_r_data; // @[SystolicConnect.scala 50:16]
  assign io_out_r_18_stop_weight = pe_mat_18_31_io_out_r_stop_weight; // @[SystolicConnect.scala 50:16]
  assign io_out_r_18_stall = pe_mat_18_31_io_out_r_stall; // @[SystolicConnect.scala 50:16]
  assign io_out_r_19_data = pe_mat_19_31_io_out_r_data; // @[SystolicConnect.scala 50:16]
  assign io_out_r_19_stop_weight = pe_mat_19_31_io_out_r_stop_weight; // @[SystolicConnect.scala 50:16]
  assign io_out_r_19_stall = pe_mat_19_31_io_out_r_stall; // @[SystolicConnect.scala 50:16]
  assign io_out_r_20_data = pe_mat_20_31_io_out_r_data; // @[SystolicConnect.scala 50:16]
  assign io_out_r_20_stop_weight = pe_mat_20_31_io_out_r_stop_weight; // @[SystolicConnect.scala 50:16]
  assign io_out_r_20_stall = pe_mat_20_31_io_out_r_stall; // @[SystolicConnect.scala 50:16]
  assign io_out_r_21_data = pe_mat_21_31_io_out_r_data; // @[SystolicConnect.scala 50:16]
  assign io_out_r_21_stop_weight = pe_mat_21_31_io_out_r_stop_weight; // @[SystolicConnect.scala 50:16]
  assign io_out_r_21_stall = pe_mat_21_31_io_out_r_stall; // @[SystolicConnect.scala 50:16]
  assign io_out_r_22_data = pe_mat_22_31_io_out_r_data; // @[SystolicConnect.scala 50:16]
  assign io_out_r_22_stop_weight = pe_mat_22_31_io_out_r_stop_weight; // @[SystolicConnect.scala 50:16]
  assign io_out_r_22_stall = pe_mat_22_31_io_out_r_stall; // @[SystolicConnect.scala 50:16]
  assign io_out_r_23_data = pe_mat_23_31_io_out_r_data; // @[SystolicConnect.scala 50:16]
  assign io_out_r_23_stop_weight = pe_mat_23_31_io_out_r_stop_weight; // @[SystolicConnect.scala 50:16]
  assign io_out_r_23_stall = pe_mat_23_31_io_out_r_stall; // @[SystolicConnect.scala 50:16]
  assign io_out_r_24_data = pe_mat_24_31_io_out_r_data; // @[SystolicConnect.scala 50:16]
  assign io_out_r_24_stop_weight = pe_mat_24_31_io_out_r_stop_weight; // @[SystolicConnect.scala 50:16]
  assign io_out_r_24_stall = pe_mat_24_31_io_out_r_stall; // @[SystolicConnect.scala 50:16]
  assign io_out_r_25_data = pe_mat_25_31_io_out_r_data; // @[SystolicConnect.scala 50:16]
  assign io_out_r_25_stop_weight = pe_mat_25_31_io_out_r_stop_weight; // @[SystolicConnect.scala 50:16]
  assign io_out_r_25_stall = pe_mat_25_31_io_out_r_stall; // @[SystolicConnect.scala 50:16]
  assign io_out_r_26_data = pe_mat_26_31_io_out_r_data; // @[SystolicConnect.scala 50:16]
  assign io_out_r_26_stop_weight = pe_mat_26_31_io_out_r_stop_weight; // @[SystolicConnect.scala 50:16]
  assign io_out_r_26_stall = pe_mat_26_31_io_out_r_stall; // @[SystolicConnect.scala 50:16]
  assign io_out_r_27_data = pe_mat_27_31_io_out_r_data; // @[SystolicConnect.scala 50:16]
  assign io_out_r_27_stop_weight = pe_mat_27_31_io_out_r_stop_weight; // @[SystolicConnect.scala 50:16]
  assign io_out_r_27_stall = pe_mat_27_31_io_out_r_stall; // @[SystolicConnect.scala 50:16]
  assign io_out_r_28_data = pe_mat_28_31_io_out_r_data; // @[SystolicConnect.scala 50:16]
  assign io_out_r_28_stop_weight = pe_mat_28_31_io_out_r_stop_weight; // @[SystolicConnect.scala 50:16]
  assign io_out_r_28_stall = pe_mat_28_31_io_out_r_stall; // @[SystolicConnect.scala 50:16]
  assign io_out_r_29_data = pe_mat_29_31_io_out_r_data; // @[SystolicConnect.scala 50:16]
  assign io_out_r_29_stop_weight = pe_mat_29_31_io_out_r_stop_weight; // @[SystolicConnect.scala 50:16]
  assign io_out_r_29_stall = pe_mat_29_31_io_out_r_stall; // @[SystolicConnect.scala 50:16]
  assign io_out_r_30_data = pe_mat_30_31_io_out_r_data; // @[SystolicConnect.scala 50:16]
  assign io_out_r_30_stop_weight = pe_mat_30_31_io_out_r_stop_weight; // @[SystolicConnect.scala 50:16]
  assign io_out_r_30_stall = pe_mat_30_31_io_out_r_stall; // @[SystolicConnect.scala 50:16]
  assign io_out_r_31_data = pe_mat_31_31_io_out_r_data; // @[SystolicConnect.scala 50:16]
  assign io_out_r_31_stop_weight = pe_mat_31_31_io_out_r_stop_weight; // @[SystolicConnect.scala 50:16]
  assign io_out_r_31_stall = pe_mat_31_31_io_out_r_stall; // @[SystolicConnect.scala 50:16]
  assign io_out_c_0_data = pe_mat_31_0_io_out_c_data; // @[SystolicConnect.scala 56:16]
  assign io_out_c_0_is_weight = pe_mat_31_0_io_out_c_is_weight; // @[SystolicConnect.scala 56:16]
  assign io_out_c_1_data = pe_mat_31_1_io_out_c_data; // @[SystolicConnect.scala 56:16]
  assign io_out_c_1_is_weight = pe_mat_31_1_io_out_c_is_weight; // @[SystolicConnect.scala 56:16]
  assign io_out_c_2_data = pe_mat_31_2_io_out_c_data; // @[SystolicConnect.scala 56:16]
  assign io_out_c_2_is_weight = pe_mat_31_2_io_out_c_is_weight; // @[SystolicConnect.scala 56:16]
  assign io_out_c_3_data = pe_mat_31_3_io_out_c_data; // @[SystolicConnect.scala 56:16]
  assign io_out_c_3_is_weight = pe_mat_31_3_io_out_c_is_weight; // @[SystolicConnect.scala 56:16]
  assign io_out_c_4_data = pe_mat_31_4_io_out_c_data; // @[SystolicConnect.scala 56:16]
  assign io_out_c_4_is_weight = pe_mat_31_4_io_out_c_is_weight; // @[SystolicConnect.scala 56:16]
  assign io_out_c_5_data = pe_mat_31_5_io_out_c_data; // @[SystolicConnect.scala 56:16]
  assign io_out_c_5_is_weight = pe_mat_31_5_io_out_c_is_weight; // @[SystolicConnect.scala 56:16]
  assign io_out_c_6_data = pe_mat_31_6_io_out_c_data; // @[SystolicConnect.scala 56:16]
  assign io_out_c_6_is_weight = pe_mat_31_6_io_out_c_is_weight; // @[SystolicConnect.scala 56:16]
  assign io_out_c_7_data = pe_mat_31_7_io_out_c_data; // @[SystolicConnect.scala 56:16]
  assign io_out_c_7_is_weight = pe_mat_31_7_io_out_c_is_weight; // @[SystolicConnect.scala 56:16]
  assign io_out_c_8_data = pe_mat_31_8_io_out_c_data; // @[SystolicConnect.scala 56:16]
  assign io_out_c_8_is_weight = pe_mat_31_8_io_out_c_is_weight; // @[SystolicConnect.scala 56:16]
  assign io_out_c_9_data = pe_mat_31_9_io_out_c_data; // @[SystolicConnect.scala 56:16]
  assign io_out_c_9_is_weight = pe_mat_31_9_io_out_c_is_weight; // @[SystolicConnect.scala 56:16]
  assign io_out_c_10_data = pe_mat_31_10_io_out_c_data; // @[SystolicConnect.scala 56:16]
  assign io_out_c_10_is_weight = pe_mat_31_10_io_out_c_is_weight; // @[SystolicConnect.scala 56:16]
  assign io_out_c_11_data = pe_mat_31_11_io_out_c_data; // @[SystolicConnect.scala 56:16]
  assign io_out_c_11_is_weight = pe_mat_31_11_io_out_c_is_weight; // @[SystolicConnect.scala 56:16]
  assign io_out_c_12_data = pe_mat_31_12_io_out_c_data; // @[SystolicConnect.scala 56:16]
  assign io_out_c_12_is_weight = pe_mat_31_12_io_out_c_is_weight; // @[SystolicConnect.scala 56:16]
  assign io_out_c_13_data = pe_mat_31_13_io_out_c_data; // @[SystolicConnect.scala 56:16]
  assign io_out_c_13_is_weight = pe_mat_31_13_io_out_c_is_weight; // @[SystolicConnect.scala 56:16]
  assign io_out_c_14_data = pe_mat_31_14_io_out_c_data; // @[SystolicConnect.scala 56:16]
  assign io_out_c_14_is_weight = pe_mat_31_14_io_out_c_is_weight; // @[SystolicConnect.scala 56:16]
  assign io_out_c_15_data = pe_mat_31_15_io_out_c_data; // @[SystolicConnect.scala 56:16]
  assign io_out_c_15_is_weight = pe_mat_31_15_io_out_c_is_weight; // @[SystolicConnect.scala 56:16]
  assign io_out_c_16_data = pe_mat_31_16_io_out_c_data; // @[SystolicConnect.scala 56:16]
  assign io_out_c_16_is_weight = pe_mat_31_16_io_out_c_is_weight; // @[SystolicConnect.scala 56:16]
  assign io_out_c_17_data = pe_mat_31_17_io_out_c_data; // @[SystolicConnect.scala 56:16]
  assign io_out_c_17_is_weight = pe_mat_31_17_io_out_c_is_weight; // @[SystolicConnect.scala 56:16]
  assign io_out_c_18_data = pe_mat_31_18_io_out_c_data; // @[SystolicConnect.scala 56:16]
  assign io_out_c_18_is_weight = pe_mat_31_18_io_out_c_is_weight; // @[SystolicConnect.scala 56:16]
  assign io_out_c_19_data = pe_mat_31_19_io_out_c_data; // @[SystolicConnect.scala 56:16]
  assign io_out_c_19_is_weight = pe_mat_31_19_io_out_c_is_weight; // @[SystolicConnect.scala 56:16]
  assign io_out_c_20_data = pe_mat_31_20_io_out_c_data; // @[SystolicConnect.scala 56:16]
  assign io_out_c_20_is_weight = pe_mat_31_20_io_out_c_is_weight; // @[SystolicConnect.scala 56:16]
  assign io_out_c_21_data = pe_mat_31_21_io_out_c_data; // @[SystolicConnect.scala 56:16]
  assign io_out_c_21_is_weight = pe_mat_31_21_io_out_c_is_weight; // @[SystolicConnect.scala 56:16]
  assign io_out_c_22_data = pe_mat_31_22_io_out_c_data; // @[SystolicConnect.scala 56:16]
  assign io_out_c_22_is_weight = pe_mat_31_22_io_out_c_is_weight; // @[SystolicConnect.scala 56:16]
  assign io_out_c_23_data = pe_mat_31_23_io_out_c_data; // @[SystolicConnect.scala 56:16]
  assign io_out_c_23_is_weight = pe_mat_31_23_io_out_c_is_weight; // @[SystolicConnect.scala 56:16]
  assign io_out_c_24_data = pe_mat_31_24_io_out_c_data; // @[SystolicConnect.scala 56:16]
  assign io_out_c_24_is_weight = pe_mat_31_24_io_out_c_is_weight; // @[SystolicConnect.scala 56:16]
  assign io_out_c_25_data = pe_mat_31_25_io_out_c_data; // @[SystolicConnect.scala 56:16]
  assign io_out_c_25_is_weight = pe_mat_31_25_io_out_c_is_weight; // @[SystolicConnect.scala 56:16]
  assign io_out_c_26_data = pe_mat_31_26_io_out_c_data; // @[SystolicConnect.scala 56:16]
  assign io_out_c_26_is_weight = pe_mat_31_26_io_out_c_is_weight; // @[SystolicConnect.scala 56:16]
  assign io_out_c_27_data = pe_mat_31_27_io_out_c_data; // @[SystolicConnect.scala 56:16]
  assign io_out_c_27_is_weight = pe_mat_31_27_io_out_c_is_weight; // @[SystolicConnect.scala 56:16]
  assign io_out_c_28_data = pe_mat_31_28_io_out_c_data; // @[SystolicConnect.scala 56:16]
  assign io_out_c_28_is_weight = pe_mat_31_28_io_out_c_is_weight; // @[SystolicConnect.scala 56:16]
  assign io_out_c_29_data = pe_mat_31_29_io_out_c_data; // @[SystolicConnect.scala 56:16]
  assign io_out_c_29_is_weight = pe_mat_31_29_io_out_c_is_weight; // @[SystolicConnect.scala 56:16]
  assign io_out_c_30_data = pe_mat_31_30_io_out_c_data; // @[SystolicConnect.scala 56:16]
  assign io_out_c_30_is_weight = pe_mat_31_30_io_out_c_is_weight; // @[SystolicConnect.scala 56:16]
  assign io_out_c_31_data = pe_mat_31_31_io_out_c_data; // @[SystolicConnect.scala 56:16]
  assign io_out_c_31_is_weight = pe_mat_31_31_io_out_c_is_weight; // @[SystolicConnect.scala 56:16]

endmodule

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

//PEWS_1023 replaced by PEWS_1023

module PEWS_1023 (
  input      [15:0]   io_in_r_data,
  input               io_in_r_stop_weight,
  input               io_in_r_stall,
  output     [15:0]   io_out_r_data,
  output              io_out_r_stop_weight,
  output              io_out_r_stall,
  input      [15:0]   io_in_c_data,
  input               io_in_c_is_weight,
  output     [15:0]   io_out_c_data,
  output              io_out_c_is_weight,
  input               clk,
  input               reset
);

  wire       [15:0]   mac_1024_io_result;
  wire                ctrl_not_stall;
  wire                when_PEWS_l54;
  reg        [15:0]   weight_reg;
  reg                 io_in_r_stall_regNext;
  reg        [15:0]   io_in_r_data_regNextWhen;
  reg                 io_in_r_stop_weight_regNextWhen;
  reg        [15:0]   _zz_io_out_c_data;
  reg                 io_in_c_is_weight_regNextWhen;

  Mac_1023 mac_1024 (
    .io_psum            (io_in_c_data[15:0]      ), //i
    .io_weight          (weight_reg[15:0]        ), //i
    .io_inputActivation (io_in_r_data[15:0]      ), //i
    .io_result          (mac_1024_io_result[15:0])  //o
  );
  assign ctrl_not_stall = (! io_in_r_stall); // @[BaseType.scala 299:24]
  assign when_PEWS_l54 = (io_in_r_stop_weight && ctrl_not_stall); // @[BaseType.scala 305:24]
  assign io_out_r_stall = io_in_r_stall_regNext; // @[PEWS.scala 64:18]
  assign io_out_r_data = io_in_r_data_regNextWhen; // @[PEWS.scala 65:17]
  assign io_out_r_stop_weight = io_in_r_stop_weight_regNextWhen; // @[PEWS.scala 66:24]
  assign io_out_c_data = _zz_io_out_c_data; // @[PEWS.scala 69:17]
  assign io_out_c_is_weight = io_in_c_is_weight_regNextWhen; // @[PEWS.scala 70:22]
  always @(posedge clk) begin
    if(when_PEWS_l54) begin
      weight_reg <= io_in_c_data; // @[PEWS.scala 54:31]
    end
    io_in_r_stall_regNext <= io_in_r_stall; // @[Reg.scala 39:30]
    if(ctrl_not_stall) begin
      io_in_r_data_regNextWhen <= io_in_r_data; // @[PEWS.scala 65:31]
    end
    if(ctrl_not_stall) begin
      io_in_r_stop_weight_regNextWhen <= io_in_r_stop_weight; // @[PEWS.scala 66:38]
    end
    if(ctrl_not_stall) begin
      _zz_io_out_c_data <= (io_in_c_is_weight ? io_in_c_data : mac_1024_io_result); // @[PEWS.scala 69:31]
    end
    if(ctrl_not_stall) begin
      io_in_c_is_weight_regNextWhen <= io_in_c_is_weight; // @[PEWS.scala 70:36]
    end
  end


endmodule

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

//Mac_1023 replaced by Mac_1023

module Mac_1023 (
  input      [15:0]   io_psum,
  input      [15:0]   io_weight,
  input      [15:0]   io_inputActivation,
  output     [15:0]   io_result
);

  wire       [31:0]   _zz_io_result;
  wire       [31:0]   _zz_io_result_1;
  wire       [31:0]   _zz_io_result_2;

  assign _zz_io_result = ($signed(_zz_io_result_1) + $signed(_zz_io_result_2));
  assign _zz_io_result_1 = ($signed(io_inputActivation) * $signed(io_weight));
  assign _zz_io_result_2 = {{16{io_psum[15]}}, io_psum};
  assign io_result = _zz_io_result[15:0]; // @[Mac.scala 14:31]

endmodule
