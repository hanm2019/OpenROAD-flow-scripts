// Generator : SpinalHDL v1.8.0    git head : 4e3563a282582b41f4eaafc503787757251d23ea
// Component : ArrayGemmini
// Git hash  : 880d730121882c0a9e393151e88289ab6120d150

`timescale 1ns/1ps

module ArrayGemmini (
  input      [15:0]   io_in_r_0_data,
  input               io_in_r_0_load_store,
  input               io_in_r_0_df_is_ws,
  input               io_in_r_0_stall,
  input      [15:0]   io_in_r_1_data,
  input               io_in_r_1_load_store,
  input               io_in_r_1_df_is_ws,
  input               io_in_r_1_stall,
  input      [15:0]   io_in_r_2_data,
  input               io_in_r_2_load_store,
  input               io_in_r_2_df_is_ws,
  input               io_in_r_2_stall,
  input      [15:0]   io_in_r_3_data,
  input               io_in_r_3_load_store,
  input               io_in_r_3_df_is_ws,
  input               io_in_r_3_stall,
  input      [15:0]   io_in_r_4_data,
  input               io_in_r_4_load_store,
  input               io_in_r_4_df_is_ws,
  input               io_in_r_4_stall,
  input      [15:0]   io_in_r_5_data,
  input               io_in_r_5_load_store,
  input               io_in_r_5_df_is_ws,
  input               io_in_r_5_stall,
  input      [15:0]   io_in_r_6_data,
  input               io_in_r_6_load_store,
  input               io_in_r_6_df_is_ws,
  input               io_in_r_6_stall,
  input      [15:0]   io_in_r_7_data,
  input               io_in_r_7_load_store,
  input               io_in_r_7_df_is_ws,
  input               io_in_r_7_stall,
  input      [15:0]   io_in_r_8_data,
  input               io_in_r_8_load_store,
  input               io_in_r_8_df_is_ws,
  input               io_in_r_8_stall,
  input      [15:0]   io_in_r_9_data,
  input               io_in_r_9_load_store,
  input               io_in_r_9_df_is_ws,
  input               io_in_r_9_stall,
  input      [15:0]   io_in_r_10_data,
  input               io_in_r_10_load_store,
  input               io_in_r_10_df_is_ws,
  input               io_in_r_10_stall,
  input      [15:0]   io_in_r_11_data,
  input               io_in_r_11_load_store,
  input               io_in_r_11_df_is_ws,
  input               io_in_r_11_stall,
  input      [15:0]   io_in_r_12_data,
  input               io_in_r_12_load_store,
  input               io_in_r_12_df_is_ws,
  input               io_in_r_12_stall,
  input      [15:0]   io_in_r_13_data,
  input               io_in_r_13_load_store,
  input               io_in_r_13_df_is_ws,
  input               io_in_r_13_stall,
  input      [15:0]   io_in_r_14_data,
  input               io_in_r_14_load_store,
  input               io_in_r_14_df_is_ws,
  input               io_in_r_14_stall,
  input      [15:0]   io_in_r_15_data,
  input               io_in_r_15_load_store,
  input               io_in_r_15_df_is_ws,
  input               io_in_r_15_stall,
  output     [15:0]   io_out_r_0_data,
  output              io_out_r_0_load_store,
  output              io_out_r_0_df_is_ws,
  output              io_out_r_0_stall,
  output     [15:0]   io_out_r_1_data,
  output              io_out_r_1_load_store,
  output              io_out_r_1_df_is_ws,
  output              io_out_r_1_stall,
  output     [15:0]   io_out_r_2_data,
  output              io_out_r_2_load_store,
  output              io_out_r_2_df_is_ws,
  output              io_out_r_2_stall,
  output     [15:0]   io_out_r_3_data,
  output              io_out_r_3_load_store,
  output              io_out_r_3_df_is_ws,
  output              io_out_r_3_stall,
  output     [15:0]   io_out_r_4_data,
  output              io_out_r_4_load_store,
  output              io_out_r_4_df_is_ws,
  output              io_out_r_4_stall,
  output     [15:0]   io_out_r_5_data,
  output              io_out_r_5_load_store,
  output              io_out_r_5_df_is_ws,
  output              io_out_r_5_stall,
  output     [15:0]   io_out_r_6_data,
  output              io_out_r_6_load_store,
  output              io_out_r_6_df_is_ws,
  output              io_out_r_6_stall,
  output     [15:0]   io_out_r_7_data,
  output              io_out_r_7_load_store,
  output              io_out_r_7_df_is_ws,
  output              io_out_r_7_stall,
  output     [15:0]   io_out_r_8_data,
  output              io_out_r_8_load_store,
  output              io_out_r_8_df_is_ws,
  output              io_out_r_8_stall,
  output     [15:0]   io_out_r_9_data,
  output              io_out_r_9_load_store,
  output              io_out_r_9_df_is_ws,
  output              io_out_r_9_stall,
  output     [15:0]   io_out_r_10_data,
  output              io_out_r_10_load_store,
  output              io_out_r_10_df_is_ws,
  output              io_out_r_10_stall,
  output     [15:0]   io_out_r_11_data,
  output              io_out_r_11_load_store,
  output              io_out_r_11_df_is_ws,
  output              io_out_r_11_stall,
  output     [15:0]   io_out_r_12_data,
  output              io_out_r_12_load_store,
  output              io_out_r_12_df_is_ws,
  output              io_out_r_12_stall,
  output     [15:0]   io_out_r_13_data,
  output              io_out_r_13_load_store,
  output              io_out_r_13_df_is_ws,
  output              io_out_r_13_stall,
  output     [15:0]   io_out_r_14_data,
  output              io_out_r_14_load_store,
  output              io_out_r_14_df_is_ws,
  output              io_out_r_14_stall,
  output     [15:0]   io_out_r_15_data,
  output              io_out_r_15_load_store,
  output              io_out_r_15_df_is_ws,
  output              io_out_r_15_stall,
  input      [15:0]   io_in_c_0_data,
  input               io_in_c_0_is_stationary,
  input      [15:0]   io_in_c_1_data,
  input               io_in_c_1_is_stationary,
  input      [15:0]   io_in_c_2_data,
  input               io_in_c_2_is_stationary,
  input      [15:0]   io_in_c_3_data,
  input               io_in_c_3_is_stationary,
  input      [15:0]   io_in_c_4_data,
  input               io_in_c_4_is_stationary,
  input      [15:0]   io_in_c_5_data,
  input               io_in_c_5_is_stationary,
  input      [15:0]   io_in_c_6_data,
  input               io_in_c_6_is_stationary,
  input      [15:0]   io_in_c_7_data,
  input               io_in_c_7_is_stationary,
  input      [15:0]   io_in_c_8_data,
  input               io_in_c_8_is_stationary,
  input      [15:0]   io_in_c_9_data,
  input               io_in_c_9_is_stationary,
  input      [15:0]   io_in_c_10_data,
  input               io_in_c_10_is_stationary,
  input      [15:0]   io_in_c_11_data,
  input               io_in_c_11_is_stationary,
  input      [15:0]   io_in_c_12_data,
  input               io_in_c_12_is_stationary,
  input      [15:0]   io_in_c_13_data,
  input               io_in_c_13_is_stationary,
  input      [15:0]   io_in_c_14_data,
  input               io_in_c_14_is_stationary,
  input      [15:0]   io_in_c_15_data,
  input               io_in_c_15_is_stationary,
  output     [15:0]   io_out_c_0_data,
  output              io_out_c_0_is_stationary,
  output     [15:0]   io_out_c_1_data,
  output              io_out_c_1_is_stationary,
  output     [15:0]   io_out_c_2_data,
  output              io_out_c_2_is_stationary,
  output     [15:0]   io_out_c_3_data,
  output              io_out_c_3_is_stationary,
  output     [15:0]   io_out_c_4_data,
  output              io_out_c_4_is_stationary,
  output     [15:0]   io_out_c_5_data,
  output              io_out_c_5_is_stationary,
  output     [15:0]   io_out_c_6_data,
  output              io_out_c_6_is_stationary,
  output     [15:0]   io_out_c_7_data,
  output              io_out_c_7_is_stationary,
  output     [15:0]   io_out_c_8_data,
  output              io_out_c_8_is_stationary,
  output     [15:0]   io_out_c_9_data,
  output              io_out_c_9_is_stationary,
  output     [15:0]   io_out_c_10_data,
  output              io_out_c_10_is_stationary,
  output     [15:0]   io_out_c_11_data,
  output              io_out_c_11_is_stationary,
  output     [15:0]   io_out_c_12_data,
  output              io_out_c_12_is_stationary,
  output     [15:0]   io_out_c_13_data,
  output              io_out_c_13_is_stationary,
  output     [15:0]   io_out_c_14_data,
  output              io_out_c_14_is_stationary,
  output     [15:0]   io_out_c_15_data,
  output              io_out_c_15_is_stationary,
  input               clk,
  input               reset
);

  wire       [15:0]   pe_mat_0_0_io_out_r_data;
  wire                pe_mat_0_0_io_out_r_load_store;
  wire                pe_mat_0_0_io_out_r_df_is_ws;
  wire                pe_mat_0_0_io_out_r_stall;
  wire       [15:0]   pe_mat_0_0_io_out_c_data;
  wire                pe_mat_0_0_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_0_1_io_out_r_data;
  wire                pe_mat_0_1_io_out_r_load_store;
  wire                pe_mat_0_1_io_out_r_df_is_ws;
  wire                pe_mat_0_1_io_out_r_stall;
  wire       [15:0]   pe_mat_0_1_io_out_c_data;
  wire                pe_mat_0_1_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_0_2_io_out_r_data;
  wire                pe_mat_0_2_io_out_r_load_store;
  wire                pe_mat_0_2_io_out_r_df_is_ws;
  wire                pe_mat_0_2_io_out_r_stall;
  wire       [15:0]   pe_mat_0_2_io_out_c_data;
  wire                pe_mat_0_2_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_0_3_io_out_r_data;
  wire                pe_mat_0_3_io_out_r_load_store;
  wire                pe_mat_0_3_io_out_r_df_is_ws;
  wire                pe_mat_0_3_io_out_r_stall;
  wire       [15:0]   pe_mat_0_3_io_out_c_data;
  wire                pe_mat_0_3_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_0_4_io_out_r_data;
  wire                pe_mat_0_4_io_out_r_load_store;
  wire                pe_mat_0_4_io_out_r_df_is_ws;
  wire                pe_mat_0_4_io_out_r_stall;
  wire       [15:0]   pe_mat_0_4_io_out_c_data;
  wire                pe_mat_0_4_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_0_5_io_out_r_data;
  wire                pe_mat_0_5_io_out_r_load_store;
  wire                pe_mat_0_5_io_out_r_df_is_ws;
  wire                pe_mat_0_5_io_out_r_stall;
  wire       [15:0]   pe_mat_0_5_io_out_c_data;
  wire                pe_mat_0_5_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_0_6_io_out_r_data;
  wire                pe_mat_0_6_io_out_r_load_store;
  wire                pe_mat_0_6_io_out_r_df_is_ws;
  wire                pe_mat_0_6_io_out_r_stall;
  wire       [15:0]   pe_mat_0_6_io_out_c_data;
  wire                pe_mat_0_6_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_0_7_io_out_r_data;
  wire                pe_mat_0_7_io_out_r_load_store;
  wire                pe_mat_0_7_io_out_r_df_is_ws;
  wire                pe_mat_0_7_io_out_r_stall;
  wire       [15:0]   pe_mat_0_7_io_out_c_data;
  wire                pe_mat_0_7_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_0_8_io_out_r_data;
  wire                pe_mat_0_8_io_out_r_load_store;
  wire                pe_mat_0_8_io_out_r_df_is_ws;
  wire                pe_mat_0_8_io_out_r_stall;
  wire       [15:0]   pe_mat_0_8_io_out_c_data;
  wire                pe_mat_0_8_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_0_9_io_out_r_data;
  wire                pe_mat_0_9_io_out_r_load_store;
  wire                pe_mat_0_9_io_out_r_df_is_ws;
  wire                pe_mat_0_9_io_out_r_stall;
  wire       [15:0]   pe_mat_0_9_io_out_c_data;
  wire                pe_mat_0_9_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_0_10_io_out_r_data;
  wire                pe_mat_0_10_io_out_r_load_store;
  wire                pe_mat_0_10_io_out_r_df_is_ws;
  wire                pe_mat_0_10_io_out_r_stall;
  wire       [15:0]   pe_mat_0_10_io_out_c_data;
  wire                pe_mat_0_10_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_0_11_io_out_r_data;
  wire                pe_mat_0_11_io_out_r_load_store;
  wire                pe_mat_0_11_io_out_r_df_is_ws;
  wire                pe_mat_0_11_io_out_r_stall;
  wire       [15:0]   pe_mat_0_11_io_out_c_data;
  wire                pe_mat_0_11_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_0_12_io_out_r_data;
  wire                pe_mat_0_12_io_out_r_load_store;
  wire                pe_mat_0_12_io_out_r_df_is_ws;
  wire                pe_mat_0_12_io_out_r_stall;
  wire       [15:0]   pe_mat_0_12_io_out_c_data;
  wire                pe_mat_0_12_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_0_13_io_out_r_data;
  wire                pe_mat_0_13_io_out_r_load_store;
  wire                pe_mat_0_13_io_out_r_df_is_ws;
  wire                pe_mat_0_13_io_out_r_stall;
  wire       [15:0]   pe_mat_0_13_io_out_c_data;
  wire                pe_mat_0_13_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_0_14_io_out_r_data;
  wire                pe_mat_0_14_io_out_r_load_store;
  wire                pe_mat_0_14_io_out_r_df_is_ws;
  wire                pe_mat_0_14_io_out_r_stall;
  wire       [15:0]   pe_mat_0_14_io_out_c_data;
  wire                pe_mat_0_14_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_0_15_io_out_r_data;
  wire                pe_mat_0_15_io_out_r_load_store;
  wire                pe_mat_0_15_io_out_r_df_is_ws;
  wire                pe_mat_0_15_io_out_r_stall;
  wire       [15:0]   pe_mat_0_15_io_out_c_data;
  wire                pe_mat_0_15_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_1_0_io_out_r_data;
  wire                pe_mat_1_0_io_out_r_load_store;
  wire                pe_mat_1_0_io_out_r_df_is_ws;
  wire                pe_mat_1_0_io_out_r_stall;
  wire       [15:0]   pe_mat_1_0_io_out_c_data;
  wire                pe_mat_1_0_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_1_1_io_out_r_data;
  wire                pe_mat_1_1_io_out_r_load_store;
  wire                pe_mat_1_1_io_out_r_df_is_ws;
  wire                pe_mat_1_1_io_out_r_stall;
  wire       [15:0]   pe_mat_1_1_io_out_c_data;
  wire                pe_mat_1_1_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_1_2_io_out_r_data;
  wire                pe_mat_1_2_io_out_r_load_store;
  wire                pe_mat_1_2_io_out_r_df_is_ws;
  wire                pe_mat_1_2_io_out_r_stall;
  wire       [15:0]   pe_mat_1_2_io_out_c_data;
  wire                pe_mat_1_2_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_1_3_io_out_r_data;
  wire                pe_mat_1_3_io_out_r_load_store;
  wire                pe_mat_1_3_io_out_r_df_is_ws;
  wire                pe_mat_1_3_io_out_r_stall;
  wire       [15:0]   pe_mat_1_3_io_out_c_data;
  wire                pe_mat_1_3_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_1_4_io_out_r_data;
  wire                pe_mat_1_4_io_out_r_load_store;
  wire                pe_mat_1_4_io_out_r_df_is_ws;
  wire                pe_mat_1_4_io_out_r_stall;
  wire       [15:0]   pe_mat_1_4_io_out_c_data;
  wire                pe_mat_1_4_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_1_5_io_out_r_data;
  wire                pe_mat_1_5_io_out_r_load_store;
  wire                pe_mat_1_5_io_out_r_df_is_ws;
  wire                pe_mat_1_5_io_out_r_stall;
  wire       [15:0]   pe_mat_1_5_io_out_c_data;
  wire                pe_mat_1_5_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_1_6_io_out_r_data;
  wire                pe_mat_1_6_io_out_r_load_store;
  wire                pe_mat_1_6_io_out_r_df_is_ws;
  wire                pe_mat_1_6_io_out_r_stall;
  wire       [15:0]   pe_mat_1_6_io_out_c_data;
  wire                pe_mat_1_6_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_1_7_io_out_r_data;
  wire                pe_mat_1_7_io_out_r_load_store;
  wire                pe_mat_1_7_io_out_r_df_is_ws;
  wire                pe_mat_1_7_io_out_r_stall;
  wire       [15:0]   pe_mat_1_7_io_out_c_data;
  wire                pe_mat_1_7_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_1_8_io_out_r_data;
  wire                pe_mat_1_8_io_out_r_load_store;
  wire                pe_mat_1_8_io_out_r_df_is_ws;
  wire                pe_mat_1_8_io_out_r_stall;
  wire       [15:0]   pe_mat_1_8_io_out_c_data;
  wire                pe_mat_1_8_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_1_9_io_out_r_data;
  wire                pe_mat_1_9_io_out_r_load_store;
  wire                pe_mat_1_9_io_out_r_df_is_ws;
  wire                pe_mat_1_9_io_out_r_stall;
  wire       [15:0]   pe_mat_1_9_io_out_c_data;
  wire                pe_mat_1_9_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_1_10_io_out_r_data;
  wire                pe_mat_1_10_io_out_r_load_store;
  wire                pe_mat_1_10_io_out_r_df_is_ws;
  wire                pe_mat_1_10_io_out_r_stall;
  wire       [15:0]   pe_mat_1_10_io_out_c_data;
  wire                pe_mat_1_10_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_1_11_io_out_r_data;
  wire                pe_mat_1_11_io_out_r_load_store;
  wire                pe_mat_1_11_io_out_r_df_is_ws;
  wire                pe_mat_1_11_io_out_r_stall;
  wire       [15:0]   pe_mat_1_11_io_out_c_data;
  wire                pe_mat_1_11_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_1_12_io_out_r_data;
  wire                pe_mat_1_12_io_out_r_load_store;
  wire                pe_mat_1_12_io_out_r_df_is_ws;
  wire                pe_mat_1_12_io_out_r_stall;
  wire       [15:0]   pe_mat_1_12_io_out_c_data;
  wire                pe_mat_1_12_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_1_13_io_out_r_data;
  wire                pe_mat_1_13_io_out_r_load_store;
  wire                pe_mat_1_13_io_out_r_df_is_ws;
  wire                pe_mat_1_13_io_out_r_stall;
  wire       [15:0]   pe_mat_1_13_io_out_c_data;
  wire                pe_mat_1_13_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_1_14_io_out_r_data;
  wire                pe_mat_1_14_io_out_r_load_store;
  wire                pe_mat_1_14_io_out_r_df_is_ws;
  wire                pe_mat_1_14_io_out_r_stall;
  wire       [15:0]   pe_mat_1_14_io_out_c_data;
  wire                pe_mat_1_14_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_1_15_io_out_r_data;
  wire                pe_mat_1_15_io_out_r_load_store;
  wire                pe_mat_1_15_io_out_r_df_is_ws;
  wire                pe_mat_1_15_io_out_r_stall;
  wire       [15:0]   pe_mat_1_15_io_out_c_data;
  wire                pe_mat_1_15_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_2_0_io_out_r_data;
  wire                pe_mat_2_0_io_out_r_load_store;
  wire                pe_mat_2_0_io_out_r_df_is_ws;
  wire                pe_mat_2_0_io_out_r_stall;
  wire       [15:0]   pe_mat_2_0_io_out_c_data;
  wire                pe_mat_2_0_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_2_1_io_out_r_data;
  wire                pe_mat_2_1_io_out_r_load_store;
  wire                pe_mat_2_1_io_out_r_df_is_ws;
  wire                pe_mat_2_1_io_out_r_stall;
  wire       [15:0]   pe_mat_2_1_io_out_c_data;
  wire                pe_mat_2_1_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_2_2_io_out_r_data;
  wire                pe_mat_2_2_io_out_r_load_store;
  wire                pe_mat_2_2_io_out_r_df_is_ws;
  wire                pe_mat_2_2_io_out_r_stall;
  wire       [15:0]   pe_mat_2_2_io_out_c_data;
  wire                pe_mat_2_2_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_2_3_io_out_r_data;
  wire                pe_mat_2_3_io_out_r_load_store;
  wire                pe_mat_2_3_io_out_r_df_is_ws;
  wire                pe_mat_2_3_io_out_r_stall;
  wire       [15:0]   pe_mat_2_3_io_out_c_data;
  wire                pe_mat_2_3_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_2_4_io_out_r_data;
  wire                pe_mat_2_4_io_out_r_load_store;
  wire                pe_mat_2_4_io_out_r_df_is_ws;
  wire                pe_mat_2_4_io_out_r_stall;
  wire       [15:0]   pe_mat_2_4_io_out_c_data;
  wire                pe_mat_2_4_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_2_5_io_out_r_data;
  wire                pe_mat_2_5_io_out_r_load_store;
  wire                pe_mat_2_5_io_out_r_df_is_ws;
  wire                pe_mat_2_5_io_out_r_stall;
  wire       [15:0]   pe_mat_2_5_io_out_c_data;
  wire                pe_mat_2_5_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_2_6_io_out_r_data;
  wire                pe_mat_2_6_io_out_r_load_store;
  wire                pe_mat_2_6_io_out_r_df_is_ws;
  wire                pe_mat_2_6_io_out_r_stall;
  wire       [15:0]   pe_mat_2_6_io_out_c_data;
  wire                pe_mat_2_6_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_2_7_io_out_r_data;
  wire                pe_mat_2_7_io_out_r_load_store;
  wire                pe_mat_2_7_io_out_r_df_is_ws;
  wire                pe_mat_2_7_io_out_r_stall;
  wire       [15:0]   pe_mat_2_7_io_out_c_data;
  wire                pe_mat_2_7_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_2_8_io_out_r_data;
  wire                pe_mat_2_8_io_out_r_load_store;
  wire                pe_mat_2_8_io_out_r_df_is_ws;
  wire                pe_mat_2_8_io_out_r_stall;
  wire       [15:0]   pe_mat_2_8_io_out_c_data;
  wire                pe_mat_2_8_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_2_9_io_out_r_data;
  wire                pe_mat_2_9_io_out_r_load_store;
  wire                pe_mat_2_9_io_out_r_df_is_ws;
  wire                pe_mat_2_9_io_out_r_stall;
  wire       [15:0]   pe_mat_2_9_io_out_c_data;
  wire                pe_mat_2_9_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_2_10_io_out_r_data;
  wire                pe_mat_2_10_io_out_r_load_store;
  wire                pe_mat_2_10_io_out_r_df_is_ws;
  wire                pe_mat_2_10_io_out_r_stall;
  wire       [15:0]   pe_mat_2_10_io_out_c_data;
  wire                pe_mat_2_10_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_2_11_io_out_r_data;
  wire                pe_mat_2_11_io_out_r_load_store;
  wire                pe_mat_2_11_io_out_r_df_is_ws;
  wire                pe_mat_2_11_io_out_r_stall;
  wire       [15:0]   pe_mat_2_11_io_out_c_data;
  wire                pe_mat_2_11_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_2_12_io_out_r_data;
  wire                pe_mat_2_12_io_out_r_load_store;
  wire                pe_mat_2_12_io_out_r_df_is_ws;
  wire                pe_mat_2_12_io_out_r_stall;
  wire       [15:0]   pe_mat_2_12_io_out_c_data;
  wire                pe_mat_2_12_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_2_13_io_out_r_data;
  wire                pe_mat_2_13_io_out_r_load_store;
  wire                pe_mat_2_13_io_out_r_df_is_ws;
  wire                pe_mat_2_13_io_out_r_stall;
  wire       [15:0]   pe_mat_2_13_io_out_c_data;
  wire                pe_mat_2_13_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_2_14_io_out_r_data;
  wire                pe_mat_2_14_io_out_r_load_store;
  wire                pe_mat_2_14_io_out_r_df_is_ws;
  wire                pe_mat_2_14_io_out_r_stall;
  wire       [15:0]   pe_mat_2_14_io_out_c_data;
  wire                pe_mat_2_14_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_2_15_io_out_r_data;
  wire                pe_mat_2_15_io_out_r_load_store;
  wire                pe_mat_2_15_io_out_r_df_is_ws;
  wire                pe_mat_2_15_io_out_r_stall;
  wire       [15:0]   pe_mat_2_15_io_out_c_data;
  wire                pe_mat_2_15_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_3_0_io_out_r_data;
  wire                pe_mat_3_0_io_out_r_load_store;
  wire                pe_mat_3_0_io_out_r_df_is_ws;
  wire                pe_mat_3_0_io_out_r_stall;
  wire       [15:0]   pe_mat_3_0_io_out_c_data;
  wire                pe_mat_3_0_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_3_1_io_out_r_data;
  wire                pe_mat_3_1_io_out_r_load_store;
  wire                pe_mat_3_1_io_out_r_df_is_ws;
  wire                pe_mat_3_1_io_out_r_stall;
  wire       [15:0]   pe_mat_3_1_io_out_c_data;
  wire                pe_mat_3_1_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_3_2_io_out_r_data;
  wire                pe_mat_3_2_io_out_r_load_store;
  wire                pe_mat_3_2_io_out_r_df_is_ws;
  wire                pe_mat_3_2_io_out_r_stall;
  wire       [15:0]   pe_mat_3_2_io_out_c_data;
  wire                pe_mat_3_2_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_3_3_io_out_r_data;
  wire                pe_mat_3_3_io_out_r_load_store;
  wire                pe_mat_3_3_io_out_r_df_is_ws;
  wire                pe_mat_3_3_io_out_r_stall;
  wire       [15:0]   pe_mat_3_3_io_out_c_data;
  wire                pe_mat_3_3_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_3_4_io_out_r_data;
  wire                pe_mat_3_4_io_out_r_load_store;
  wire                pe_mat_3_4_io_out_r_df_is_ws;
  wire                pe_mat_3_4_io_out_r_stall;
  wire       [15:0]   pe_mat_3_4_io_out_c_data;
  wire                pe_mat_3_4_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_3_5_io_out_r_data;
  wire                pe_mat_3_5_io_out_r_load_store;
  wire                pe_mat_3_5_io_out_r_df_is_ws;
  wire                pe_mat_3_5_io_out_r_stall;
  wire       [15:0]   pe_mat_3_5_io_out_c_data;
  wire                pe_mat_3_5_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_3_6_io_out_r_data;
  wire                pe_mat_3_6_io_out_r_load_store;
  wire                pe_mat_3_6_io_out_r_df_is_ws;
  wire                pe_mat_3_6_io_out_r_stall;
  wire       [15:0]   pe_mat_3_6_io_out_c_data;
  wire                pe_mat_3_6_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_3_7_io_out_r_data;
  wire                pe_mat_3_7_io_out_r_load_store;
  wire                pe_mat_3_7_io_out_r_df_is_ws;
  wire                pe_mat_3_7_io_out_r_stall;
  wire       [15:0]   pe_mat_3_7_io_out_c_data;
  wire                pe_mat_3_7_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_3_8_io_out_r_data;
  wire                pe_mat_3_8_io_out_r_load_store;
  wire                pe_mat_3_8_io_out_r_df_is_ws;
  wire                pe_mat_3_8_io_out_r_stall;
  wire       [15:0]   pe_mat_3_8_io_out_c_data;
  wire                pe_mat_3_8_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_3_9_io_out_r_data;
  wire                pe_mat_3_9_io_out_r_load_store;
  wire                pe_mat_3_9_io_out_r_df_is_ws;
  wire                pe_mat_3_9_io_out_r_stall;
  wire       [15:0]   pe_mat_3_9_io_out_c_data;
  wire                pe_mat_3_9_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_3_10_io_out_r_data;
  wire                pe_mat_3_10_io_out_r_load_store;
  wire                pe_mat_3_10_io_out_r_df_is_ws;
  wire                pe_mat_3_10_io_out_r_stall;
  wire       [15:0]   pe_mat_3_10_io_out_c_data;
  wire                pe_mat_3_10_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_3_11_io_out_r_data;
  wire                pe_mat_3_11_io_out_r_load_store;
  wire                pe_mat_3_11_io_out_r_df_is_ws;
  wire                pe_mat_3_11_io_out_r_stall;
  wire       [15:0]   pe_mat_3_11_io_out_c_data;
  wire                pe_mat_3_11_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_3_12_io_out_r_data;
  wire                pe_mat_3_12_io_out_r_load_store;
  wire                pe_mat_3_12_io_out_r_df_is_ws;
  wire                pe_mat_3_12_io_out_r_stall;
  wire       [15:0]   pe_mat_3_12_io_out_c_data;
  wire                pe_mat_3_12_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_3_13_io_out_r_data;
  wire                pe_mat_3_13_io_out_r_load_store;
  wire                pe_mat_3_13_io_out_r_df_is_ws;
  wire                pe_mat_3_13_io_out_r_stall;
  wire       [15:0]   pe_mat_3_13_io_out_c_data;
  wire                pe_mat_3_13_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_3_14_io_out_r_data;
  wire                pe_mat_3_14_io_out_r_load_store;
  wire                pe_mat_3_14_io_out_r_df_is_ws;
  wire                pe_mat_3_14_io_out_r_stall;
  wire       [15:0]   pe_mat_3_14_io_out_c_data;
  wire                pe_mat_3_14_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_3_15_io_out_r_data;
  wire                pe_mat_3_15_io_out_r_load_store;
  wire                pe_mat_3_15_io_out_r_df_is_ws;
  wire                pe_mat_3_15_io_out_r_stall;
  wire       [15:0]   pe_mat_3_15_io_out_c_data;
  wire                pe_mat_3_15_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_4_0_io_out_r_data;
  wire                pe_mat_4_0_io_out_r_load_store;
  wire                pe_mat_4_0_io_out_r_df_is_ws;
  wire                pe_mat_4_0_io_out_r_stall;
  wire       [15:0]   pe_mat_4_0_io_out_c_data;
  wire                pe_mat_4_0_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_4_1_io_out_r_data;
  wire                pe_mat_4_1_io_out_r_load_store;
  wire                pe_mat_4_1_io_out_r_df_is_ws;
  wire                pe_mat_4_1_io_out_r_stall;
  wire       [15:0]   pe_mat_4_1_io_out_c_data;
  wire                pe_mat_4_1_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_4_2_io_out_r_data;
  wire                pe_mat_4_2_io_out_r_load_store;
  wire                pe_mat_4_2_io_out_r_df_is_ws;
  wire                pe_mat_4_2_io_out_r_stall;
  wire       [15:0]   pe_mat_4_2_io_out_c_data;
  wire                pe_mat_4_2_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_4_3_io_out_r_data;
  wire                pe_mat_4_3_io_out_r_load_store;
  wire                pe_mat_4_3_io_out_r_df_is_ws;
  wire                pe_mat_4_3_io_out_r_stall;
  wire       [15:0]   pe_mat_4_3_io_out_c_data;
  wire                pe_mat_4_3_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_4_4_io_out_r_data;
  wire                pe_mat_4_4_io_out_r_load_store;
  wire                pe_mat_4_4_io_out_r_df_is_ws;
  wire                pe_mat_4_4_io_out_r_stall;
  wire       [15:0]   pe_mat_4_4_io_out_c_data;
  wire                pe_mat_4_4_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_4_5_io_out_r_data;
  wire                pe_mat_4_5_io_out_r_load_store;
  wire                pe_mat_4_5_io_out_r_df_is_ws;
  wire                pe_mat_4_5_io_out_r_stall;
  wire       [15:0]   pe_mat_4_5_io_out_c_data;
  wire                pe_mat_4_5_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_4_6_io_out_r_data;
  wire                pe_mat_4_6_io_out_r_load_store;
  wire                pe_mat_4_6_io_out_r_df_is_ws;
  wire                pe_mat_4_6_io_out_r_stall;
  wire       [15:0]   pe_mat_4_6_io_out_c_data;
  wire                pe_mat_4_6_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_4_7_io_out_r_data;
  wire                pe_mat_4_7_io_out_r_load_store;
  wire                pe_mat_4_7_io_out_r_df_is_ws;
  wire                pe_mat_4_7_io_out_r_stall;
  wire       [15:0]   pe_mat_4_7_io_out_c_data;
  wire                pe_mat_4_7_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_4_8_io_out_r_data;
  wire                pe_mat_4_8_io_out_r_load_store;
  wire                pe_mat_4_8_io_out_r_df_is_ws;
  wire                pe_mat_4_8_io_out_r_stall;
  wire       [15:0]   pe_mat_4_8_io_out_c_data;
  wire                pe_mat_4_8_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_4_9_io_out_r_data;
  wire                pe_mat_4_9_io_out_r_load_store;
  wire                pe_mat_4_9_io_out_r_df_is_ws;
  wire                pe_mat_4_9_io_out_r_stall;
  wire       [15:0]   pe_mat_4_9_io_out_c_data;
  wire                pe_mat_4_9_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_4_10_io_out_r_data;
  wire                pe_mat_4_10_io_out_r_load_store;
  wire                pe_mat_4_10_io_out_r_df_is_ws;
  wire                pe_mat_4_10_io_out_r_stall;
  wire       [15:0]   pe_mat_4_10_io_out_c_data;
  wire                pe_mat_4_10_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_4_11_io_out_r_data;
  wire                pe_mat_4_11_io_out_r_load_store;
  wire                pe_mat_4_11_io_out_r_df_is_ws;
  wire                pe_mat_4_11_io_out_r_stall;
  wire       [15:0]   pe_mat_4_11_io_out_c_data;
  wire                pe_mat_4_11_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_4_12_io_out_r_data;
  wire                pe_mat_4_12_io_out_r_load_store;
  wire                pe_mat_4_12_io_out_r_df_is_ws;
  wire                pe_mat_4_12_io_out_r_stall;
  wire       [15:0]   pe_mat_4_12_io_out_c_data;
  wire                pe_mat_4_12_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_4_13_io_out_r_data;
  wire                pe_mat_4_13_io_out_r_load_store;
  wire                pe_mat_4_13_io_out_r_df_is_ws;
  wire                pe_mat_4_13_io_out_r_stall;
  wire       [15:0]   pe_mat_4_13_io_out_c_data;
  wire                pe_mat_4_13_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_4_14_io_out_r_data;
  wire                pe_mat_4_14_io_out_r_load_store;
  wire                pe_mat_4_14_io_out_r_df_is_ws;
  wire                pe_mat_4_14_io_out_r_stall;
  wire       [15:0]   pe_mat_4_14_io_out_c_data;
  wire                pe_mat_4_14_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_4_15_io_out_r_data;
  wire                pe_mat_4_15_io_out_r_load_store;
  wire                pe_mat_4_15_io_out_r_df_is_ws;
  wire                pe_mat_4_15_io_out_r_stall;
  wire       [15:0]   pe_mat_4_15_io_out_c_data;
  wire                pe_mat_4_15_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_5_0_io_out_r_data;
  wire                pe_mat_5_0_io_out_r_load_store;
  wire                pe_mat_5_0_io_out_r_df_is_ws;
  wire                pe_mat_5_0_io_out_r_stall;
  wire       [15:0]   pe_mat_5_0_io_out_c_data;
  wire                pe_mat_5_0_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_5_1_io_out_r_data;
  wire                pe_mat_5_1_io_out_r_load_store;
  wire                pe_mat_5_1_io_out_r_df_is_ws;
  wire                pe_mat_5_1_io_out_r_stall;
  wire       [15:0]   pe_mat_5_1_io_out_c_data;
  wire                pe_mat_5_1_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_5_2_io_out_r_data;
  wire                pe_mat_5_2_io_out_r_load_store;
  wire                pe_mat_5_2_io_out_r_df_is_ws;
  wire                pe_mat_5_2_io_out_r_stall;
  wire       [15:0]   pe_mat_5_2_io_out_c_data;
  wire                pe_mat_5_2_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_5_3_io_out_r_data;
  wire                pe_mat_5_3_io_out_r_load_store;
  wire                pe_mat_5_3_io_out_r_df_is_ws;
  wire                pe_mat_5_3_io_out_r_stall;
  wire       [15:0]   pe_mat_5_3_io_out_c_data;
  wire                pe_mat_5_3_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_5_4_io_out_r_data;
  wire                pe_mat_5_4_io_out_r_load_store;
  wire                pe_mat_5_4_io_out_r_df_is_ws;
  wire                pe_mat_5_4_io_out_r_stall;
  wire       [15:0]   pe_mat_5_4_io_out_c_data;
  wire                pe_mat_5_4_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_5_5_io_out_r_data;
  wire                pe_mat_5_5_io_out_r_load_store;
  wire                pe_mat_5_5_io_out_r_df_is_ws;
  wire                pe_mat_5_5_io_out_r_stall;
  wire       [15:0]   pe_mat_5_5_io_out_c_data;
  wire                pe_mat_5_5_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_5_6_io_out_r_data;
  wire                pe_mat_5_6_io_out_r_load_store;
  wire                pe_mat_5_6_io_out_r_df_is_ws;
  wire                pe_mat_5_6_io_out_r_stall;
  wire       [15:0]   pe_mat_5_6_io_out_c_data;
  wire                pe_mat_5_6_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_5_7_io_out_r_data;
  wire                pe_mat_5_7_io_out_r_load_store;
  wire                pe_mat_5_7_io_out_r_df_is_ws;
  wire                pe_mat_5_7_io_out_r_stall;
  wire       [15:0]   pe_mat_5_7_io_out_c_data;
  wire                pe_mat_5_7_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_5_8_io_out_r_data;
  wire                pe_mat_5_8_io_out_r_load_store;
  wire                pe_mat_5_8_io_out_r_df_is_ws;
  wire                pe_mat_5_8_io_out_r_stall;
  wire       [15:0]   pe_mat_5_8_io_out_c_data;
  wire                pe_mat_5_8_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_5_9_io_out_r_data;
  wire                pe_mat_5_9_io_out_r_load_store;
  wire                pe_mat_5_9_io_out_r_df_is_ws;
  wire                pe_mat_5_9_io_out_r_stall;
  wire       [15:0]   pe_mat_5_9_io_out_c_data;
  wire                pe_mat_5_9_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_5_10_io_out_r_data;
  wire                pe_mat_5_10_io_out_r_load_store;
  wire                pe_mat_5_10_io_out_r_df_is_ws;
  wire                pe_mat_5_10_io_out_r_stall;
  wire       [15:0]   pe_mat_5_10_io_out_c_data;
  wire                pe_mat_5_10_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_5_11_io_out_r_data;
  wire                pe_mat_5_11_io_out_r_load_store;
  wire                pe_mat_5_11_io_out_r_df_is_ws;
  wire                pe_mat_5_11_io_out_r_stall;
  wire       [15:0]   pe_mat_5_11_io_out_c_data;
  wire                pe_mat_5_11_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_5_12_io_out_r_data;
  wire                pe_mat_5_12_io_out_r_load_store;
  wire                pe_mat_5_12_io_out_r_df_is_ws;
  wire                pe_mat_5_12_io_out_r_stall;
  wire       [15:0]   pe_mat_5_12_io_out_c_data;
  wire                pe_mat_5_12_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_5_13_io_out_r_data;
  wire                pe_mat_5_13_io_out_r_load_store;
  wire                pe_mat_5_13_io_out_r_df_is_ws;
  wire                pe_mat_5_13_io_out_r_stall;
  wire       [15:0]   pe_mat_5_13_io_out_c_data;
  wire                pe_mat_5_13_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_5_14_io_out_r_data;
  wire                pe_mat_5_14_io_out_r_load_store;
  wire                pe_mat_5_14_io_out_r_df_is_ws;
  wire                pe_mat_5_14_io_out_r_stall;
  wire       [15:0]   pe_mat_5_14_io_out_c_data;
  wire                pe_mat_5_14_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_5_15_io_out_r_data;
  wire                pe_mat_5_15_io_out_r_load_store;
  wire                pe_mat_5_15_io_out_r_df_is_ws;
  wire                pe_mat_5_15_io_out_r_stall;
  wire       [15:0]   pe_mat_5_15_io_out_c_data;
  wire                pe_mat_5_15_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_6_0_io_out_r_data;
  wire                pe_mat_6_0_io_out_r_load_store;
  wire                pe_mat_6_0_io_out_r_df_is_ws;
  wire                pe_mat_6_0_io_out_r_stall;
  wire       [15:0]   pe_mat_6_0_io_out_c_data;
  wire                pe_mat_6_0_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_6_1_io_out_r_data;
  wire                pe_mat_6_1_io_out_r_load_store;
  wire                pe_mat_6_1_io_out_r_df_is_ws;
  wire                pe_mat_6_1_io_out_r_stall;
  wire       [15:0]   pe_mat_6_1_io_out_c_data;
  wire                pe_mat_6_1_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_6_2_io_out_r_data;
  wire                pe_mat_6_2_io_out_r_load_store;
  wire                pe_mat_6_2_io_out_r_df_is_ws;
  wire                pe_mat_6_2_io_out_r_stall;
  wire       [15:0]   pe_mat_6_2_io_out_c_data;
  wire                pe_mat_6_2_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_6_3_io_out_r_data;
  wire                pe_mat_6_3_io_out_r_load_store;
  wire                pe_mat_6_3_io_out_r_df_is_ws;
  wire                pe_mat_6_3_io_out_r_stall;
  wire       [15:0]   pe_mat_6_3_io_out_c_data;
  wire                pe_mat_6_3_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_6_4_io_out_r_data;
  wire                pe_mat_6_4_io_out_r_load_store;
  wire                pe_mat_6_4_io_out_r_df_is_ws;
  wire                pe_mat_6_4_io_out_r_stall;
  wire       [15:0]   pe_mat_6_4_io_out_c_data;
  wire                pe_mat_6_4_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_6_5_io_out_r_data;
  wire                pe_mat_6_5_io_out_r_load_store;
  wire                pe_mat_6_5_io_out_r_df_is_ws;
  wire                pe_mat_6_5_io_out_r_stall;
  wire       [15:0]   pe_mat_6_5_io_out_c_data;
  wire                pe_mat_6_5_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_6_6_io_out_r_data;
  wire                pe_mat_6_6_io_out_r_load_store;
  wire                pe_mat_6_6_io_out_r_df_is_ws;
  wire                pe_mat_6_6_io_out_r_stall;
  wire       [15:0]   pe_mat_6_6_io_out_c_data;
  wire                pe_mat_6_6_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_6_7_io_out_r_data;
  wire                pe_mat_6_7_io_out_r_load_store;
  wire                pe_mat_6_7_io_out_r_df_is_ws;
  wire                pe_mat_6_7_io_out_r_stall;
  wire       [15:0]   pe_mat_6_7_io_out_c_data;
  wire                pe_mat_6_7_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_6_8_io_out_r_data;
  wire                pe_mat_6_8_io_out_r_load_store;
  wire                pe_mat_6_8_io_out_r_df_is_ws;
  wire                pe_mat_6_8_io_out_r_stall;
  wire       [15:0]   pe_mat_6_8_io_out_c_data;
  wire                pe_mat_6_8_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_6_9_io_out_r_data;
  wire                pe_mat_6_9_io_out_r_load_store;
  wire                pe_mat_6_9_io_out_r_df_is_ws;
  wire                pe_mat_6_9_io_out_r_stall;
  wire       [15:0]   pe_mat_6_9_io_out_c_data;
  wire                pe_mat_6_9_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_6_10_io_out_r_data;
  wire                pe_mat_6_10_io_out_r_load_store;
  wire                pe_mat_6_10_io_out_r_df_is_ws;
  wire                pe_mat_6_10_io_out_r_stall;
  wire       [15:0]   pe_mat_6_10_io_out_c_data;
  wire                pe_mat_6_10_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_6_11_io_out_r_data;
  wire                pe_mat_6_11_io_out_r_load_store;
  wire                pe_mat_6_11_io_out_r_df_is_ws;
  wire                pe_mat_6_11_io_out_r_stall;
  wire       [15:0]   pe_mat_6_11_io_out_c_data;
  wire                pe_mat_6_11_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_6_12_io_out_r_data;
  wire                pe_mat_6_12_io_out_r_load_store;
  wire                pe_mat_6_12_io_out_r_df_is_ws;
  wire                pe_mat_6_12_io_out_r_stall;
  wire       [15:0]   pe_mat_6_12_io_out_c_data;
  wire                pe_mat_6_12_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_6_13_io_out_r_data;
  wire                pe_mat_6_13_io_out_r_load_store;
  wire                pe_mat_6_13_io_out_r_df_is_ws;
  wire                pe_mat_6_13_io_out_r_stall;
  wire       [15:0]   pe_mat_6_13_io_out_c_data;
  wire                pe_mat_6_13_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_6_14_io_out_r_data;
  wire                pe_mat_6_14_io_out_r_load_store;
  wire                pe_mat_6_14_io_out_r_df_is_ws;
  wire                pe_mat_6_14_io_out_r_stall;
  wire       [15:0]   pe_mat_6_14_io_out_c_data;
  wire                pe_mat_6_14_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_6_15_io_out_r_data;
  wire                pe_mat_6_15_io_out_r_load_store;
  wire                pe_mat_6_15_io_out_r_df_is_ws;
  wire                pe_mat_6_15_io_out_r_stall;
  wire       [15:0]   pe_mat_6_15_io_out_c_data;
  wire                pe_mat_6_15_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_7_0_io_out_r_data;
  wire                pe_mat_7_0_io_out_r_load_store;
  wire                pe_mat_7_0_io_out_r_df_is_ws;
  wire                pe_mat_7_0_io_out_r_stall;
  wire       [15:0]   pe_mat_7_0_io_out_c_data;
  wire                pe_mat_7_0_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_7_1_io_out_r_data;
  wire                pe_mat_7_1_io_out_r_load_store;
  wire                pe_mat_7_1_io_out_r_df_is_ws;
  wire                pe_mat_7_1_io_out_r_stall;
  wire       [15:0]   pe_mat_7_1_io_out_c_data;
  wire                pe_mat_7_1_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_7_2_io_out_r_data;
  wire                pe_mat_7_2_io_out_r_load_store;
  wire                pe_mat_7_2_io_out_r_df_is_ws;
  wire                pe_mat_7_2_io_out_r_stall;
  wire       [15:0]   pe_mat_7_2_io_out_c_data;
  wire                pe_mat_7_2_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_7_3_io_out_r_data;
  wire                pe_mat_7_3_io_out_r_load_store;
  wire                pe_mat_7_3_io_out_r_df_is_ws;
  wire                pe_mat_7_3_io_out_r_stall;
  wire       [15:0]   pe_mat_7_3_io_out_c_data;
  wire                pe_mat_7_3_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_7_4_io_out_r_data;
  wire                pe_mat_7_4_io_out_r_load_store;
  wire                pe_mat_7_4_io_out_r_df_is_ws;
  wire                pe_mat_7_4_io_out_r_stall;
  wire       [15:0]   pe_mat_7_4_io_out_c_data;
  wire                pe_mat_7_4_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_7_5_io_out_r_data;
  wire                pe_mat_7_5_io_out_r_load_store;
  wire                pe_mat_7_5_io_out_r_df_is_ws;
  wire                pe_mat_7_5_io_out_r_stall;
  wire       [15:0]   pe_mat_7_5_io_out_c_data;
  wire                pe_mat_7_5_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_7_6_io_out_r_data;
  wire                pe_mat_7_6_io_out_r_load_store;
  wire                pe_mat_7_6_io_out_r_df_is_ws;
  wire                pe_mat_7_6_io_out_r_stall;
  wire       [15:0]   pe_mat_7_6_io_out_c_data;
  wire                pe_mat_7_6_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_7_7_io_out_r_data;
  wire                pe_mat_7_7_io_out_r_load_store;
  wire                pe_mat_7_7_io_out_r_df_is_ws;
  wire                pe_mat_7_7_io_out_r_stall;
  wire       [15:0]   pe_mat_7_7_io_out_c_data;
  wire                pe_mat_7_7_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_7_8_io_out_r_data;
  wire                pe_mat_7_8_io_out_r_load_store;
  wire                pe_mat_7_8_io_out_r_df_is_ws;
  wire                pe_mat_7_8_io_out_r_stall;
  wire       [15:0]   pe_mat_7_8_io_out_c_data;
  wire                pe_mat_7_8_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_7_9_io_out_r_data;
  wire                pe_mat_7_9_io_out_r_load_store;
  wire                pe_mat_7_9_io_out_r_df_is_ws;
  wire                pe_mat_7_9_io_out_r_stall;
  wire       [15:0]   pe_mat_7_9_io_out_c_data;
  wire                pe_mat_7_9_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_7_10_io_out_r_data;
  wire                pe_mat_7_10_io_out_r_load_store;
  wire                pe_mat_7_10_io_out_r_df_is_ws;
  wire                pe_mat_7_10_io_out_r_stall;
  wire       [15:0]   pe_mat_7_10_io_out_c_data;
  wire                pe_mat_7_10_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_7_11_io_out_r_data;
  wire                pe_mat_7_11_io_out_r_load_store;
  wire                pe_mat_7_11_io_out_r_df_is_ws;
  wire                pe_mat_7_11_io_out_r_stall;
  wire       [15:0]   pe_mat_7_11_io_out_c_data;
  wire                pe_mat_7_11_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_7_12_io_out_r_data;
  wire                pe_mat_7_12_io_out_r_load_store;
  wire                pe_mat_7_12_io_out_r_df_is_ws;
  wire                pe_mat_7_12_io_out_r_stall;
  wire       [15:0]   pe_mat_7_12_io_out_c_data;
  wire                pe_mat_7_12_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_7_13_io_out_r_data;
  wire                pe_mat_7_13_io_out_r_load_store;
  wire                pe_mat_7_13_io_out_r_df_is_ws;
  wire                pe_mat_7_13_io_out_r_stall;
  wire       [15:0]   pe_mat_7_13_io_out_c_data;
  wire                pe_mat_7_13_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_7_14_io_out_r_data;
  wire                pe_mat_7_14_io_out_r_load_store;
  wire                pe_mat_7_14_io_out_r_df_is_ws;
  wire                pe_mat_7_14_io_out_r_stall;
  wire       [15:0]   pe_mat_7_14_io_out_c_data;
  wire                pe_mat_7_14_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_7_15_io_out_r_data;
  wire                pe_mat_7_15_io_out_r_load_store;
  wire                pe_mat_7_15_io_out_r_df_is_ws;
  wire                pe_mat_7_15_io_out_r_stall;
  wire       [15:0]   pe_mat_7_15_io_out_c_data;
  wire                pe_mat_7_15_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_8_0_io_out_r_data;
  wire                pe_mat_8_0_io_out_r_load_store;
  wire                pe_mat_8_0_io_out_r_df_is_ws;
  wire                pe_mat_8_0_io_out_r_stall;
  wire       [15:0]   pe_mat_8_0_io_out_c_data;
  wire                pe_mat_8_0_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_8_1_io_out_r_data;
  wire                pe_mat_8_1_io_out_r_load_store;
  wire                pe_mat_8_1_io_out_r_df_is_ws;
  wire                pe_mat_8_1_io_out_r_stall;
  wire       [15:0]   pe_mat_8_1_io_out_c_data;
  wire                pe_mat_8_1_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_8_2_io_out_r_data;
  wire                pe_mat_8_2_io_out_r_load_store;
  wire                pe_mat_8_2_io_out_r_df_is_ws;
  wire                pe_mat_8_2_io_out_r_stall;
  wire       [15:0]   pe_mat_8_2_io_out_c_data;
  wire                pe_mat_8_2_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_8_3_io_out_r_data;
  wire                pe_mat_8_3_io_out_r_load_store;
  wire                pe_mat_8_3_io_out_r_df_is_ws;
  wire                pe_mat_8_3_io_out_r_stall;
  wire       [15:0]   pe_mat_8_3_io_out_c_data;
  wire                pe_mat_8_3_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_8_4_io_out_r_data;
  wire                pe_mat_8_4_io_out_r_load_store;
  wire                pe_mat_8_4_io_out_r_df_is_ws;
  wire                pe_mat_8_4_io_out_r_stall;
  wire       [15:0]   pe_mat_8_4_io_out_c_data;
  wire                pe_mat_8_4_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_8_5_io_out_r_data;
  wire                pe_mat_8_5_io_out_r_load_store;
  wire                pe_mat_8_5_io_out_r_df_is_ws;
  wire                pe_mat_8_5_io_out_r_stall;
  wire       [15:0]   pe_mat_8_5_io_out_c_data;
  wire                pe_mat_8_5_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_8_6_io_out_r_data;
  wire                pe_mat_8_6_io_out_r_load_store;
  wire                pe_mat_8_6_io_out_r_df_is_ws;
  wire                pe_mat_8_6_io_out_r_stall;
  wire       [15:0]   pe_mat_8_6_io_out_c_data;
  wire                pe_mat_8_6_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_8_7_io_out_r_data;
  wire                pe_mat_8_7_io_out_r_load_store;
  wire                pe_mat_8_7_io_out_r_df_is_ws;
  wire                pe_mat_8_7_io_out_r_stall;
  wire       [15:0]   pe_mat_8_7_io_out_c_data;
  wire                pe_mat_8_7_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_8_8_io_out_r_data;
  wire                pe_mat_8_8_io_out_r_load_store;
  wire                pe_mat_8_8_io_out_r_df_is_ws;
  wire                pe_mat_8_8_io_out_r_stall;
  wire       [15:0]   pe_mat_8_8_io_out_c_data;
  wire                pe_mat_8_8_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_8_9_io_out_r_data;
  wire                pe_mat_8_9_io_out_r_load_store;
  wire                pe_mat_8_9_io_out_r_df_is_ws;
  wire                pe_mat_8_9_io_out_r_stall;
  wire       [15:0]   pe_mat_8_9_io_out_c_data;
  wire                pe_mat_8_9_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_8_10_io_out_r_data;
  wire                pe_mat_8_10_io_out_r_load_store;
  wire                pe_mat_8_10_io_out_r_df_is_ws;
  wire                pe_mat_8_10_io_out_r_stall;
  wire       [15:0]   pe_mat_8_10_io_out_c_data;
  wire                pe_mat_8_10_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_8_11_io_out_r_data;
  wire                pe_mat_8_11_io_out_r_load_store;
  wire                pe_mat_8_11_io_out_r_df_is_ws;
  wire                pe_mat_8_11_io_out_r_stall;
  wire       [15:0]   pe_mat_8_11_io_out_c_data;
  wire                pe_mat_8_11_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_8_12_io_out_r_data;
  wire                pe_mat_8_12_io_out_r_load_store;
  wire                pe_mat_8_12_io_out_r_df_is_ws;
  wire                pe_mat_8_12_io_out_r_stall;
  wire       [15:0]   pe_mat_8_12_io_out_c_data;
  wire                pe_mat_8_12_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_8_13_io_out_r_data;
  wire                pe_mat_8_13_io_out_r_load_store;
  wire                pe_mat_8_13_io_out_r_df_is_ws;
  wire                pe_mat_8_13_io_out_r_stall;
  wire       [15:0]   pe_mat_8_13_io_out_c_data;
  wire                pe_mat_8_13_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_8_14_io_out_r_data;
  wire                pe_mat_8_14_io_out_r_load_store;
  wire                pe_mat_8_14_io_out_r_df_is_ws;
  wire                pe_mat_8_14_io_out_r_stall;
  wire       [15:0]   pe_mat_8_14_io_out_c_data;
  wire                pe_mat_8_14_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_8_15_io_out_r_data;
  wire                pe_mat_8_15_io_out_r_load_store;
  wire                pe_mat_8_15_io_out_r_df_is_ws;
  wire                pe_mat_8_15_io_out_r_stall;
  wire       [15:0]   pe_mat_8_15_io_out_c_data;
  wire                pe_mat_8_15_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_9_0_io_out_r_data;
  wire                pe_mat_9_0_io_out_r_load_store;
  wire                pe_mat_9_0_io_out_r_df_is_ws;
  wire                pe_mat_9_0_io_out_r_stall;
  wire       [15:0]   pe_mat_9_0_io_out_c_data;
  wire                pe_mat_9_0_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_9_1_io_out_r_data;
  wire                pe_mat_9_1_io_out_r_load_store;
  wire                pe_mat_9_1_io_out_r_df_is_ws;
  wire                pe_mat_9_1_io_out_r_stall;
  wire       [15:0]   pe_mat_9_1_io_out_c_data;
  wire                pe_mat_9_1_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_9_2_io_out_r_data;
  wire                pe_mat_9_2_io_out_r_load_store;
  wire                pe_mat_9_2_io_out_r_df_is_ws;
  wire                pe_mat_9_2_io_out_r_stall;
  wire       [15:0]   pe_mat_9_2_io_out_c_data;
  wire                pe_mat_9_2_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_9_3_io_out_r_data;
  wire                pe_mat_9_3_io_out_r_load_store;
  wire                pe_mat_9_3_io_out_r_df_is_ws;
  wire                pe_mat_9_3_io_out_r_stall;
  wire       [15:0]   pe_mat_9_3_io_out_c_data;
  wire                pe_mat_9_3_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_9_4_io_out_r_data;
  wire                pe_mat_9_4_io_out_r_load_store;
  wire                pe_mat_9_4_io_out_r_df_is_ws;
  wire                pe_mat_9_4_io_out_r_stall;
  wire       [15:0]   pe_mat_9_4_io_out_c_data;
  wire                pe_mat_9_4_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_9_5_io_out_r_data;
  wire                pe_mat_9_5_io_out_r_load_store;
  wire                pe_mat_9_5_io_out_r_df_is_ws;
  wire                pe_mat_9_5_io_out_r_stall;
  wire       [15:0]   pe_mat_9_5_io_out_c_data;
  wire                pe_mat_9_5_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_9_6_io_out_r_data;
  wire                pe_mat_9_6_io_out_r_load_store;
  wire                pe_mat_9_6_io_out_r_df_is_ws;
  wire                pe_mat_9_6_io_out_r_stall;
  wire       [15:0]   pe_mat_9_6_io_out_c_data;
  wire                pe_mat_9_6_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_9_7_io_out_r_data;
  wire                pe_mat_9_7_io_out_r_load_store;
  wire                pe_mat_9_7_io_out_r_df_is_ws;
  wire                pe_mat_9_7_io_out_r_stall;
  wire       [15:0]   pe_mat_9_7_io_out_c_data;
  wire                pe_mat_9_7_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_9_8_io_out_r_data;
  wire                pe_mat_9_8_io_out_r_load_store;
  wire                pe_mat_9_8_io_out_r_df_is_ws;
  wire                pe_mat_9_8_io_out_r_stall;
  wire       [15:0]   pe_mat_9_8_io_out_c_data;
  wire                pe_mat_9_8_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_9_9_io_out_r_data;
  wire                pe_mat_9_9_io_out_r_load_store;
  wire                pe_mat_9_9_io_out_r_df_is_ws;
  wire                pe_mat_9_9_io_out_r_stall;
  wire       [15:0]   pe_mat_9_9_io_out_c_data;
  wire                pe_mat_9_9_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_9_10_io_out_r_data;
  wire                pe_mat_9_10_io_out_r_load_store;
  wire                pe_mat_9_10_io_out_r_df_is_ws;
  wire                pe_mat_9_10_io_out_r_stall;
  wire       [15:0]   pe_mat_9_10_io_out_c_data;
  wire                pe_mat_9_10_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_9_11_io_out_r_data;
  wire                pe_mat_9_11_io_out_r_load_store;
  wire                pe_mat_9_11_io_out_r_df_is_ws;
  wire                pe_mat_9_11_io_out_r_stall;
  wire       [15:0]   pe_mat_9_11_io_out_c_data;
  wire                pe_mat_9_11_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_9_12_io_out_r_data;
  wire                pe_mat_9_12_io_out_r_load_store;
  wire                pe_mat_9_12_io_out_r_df_is_ws;
  wire                pe_mat_9_12_io_out_r_stall;
  wire       [15:0]   pe_mat_9_12_io_out_c_data;
  wire                pe_mat_9_12_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_9_13_io_out_r_data;
  wire                pe_mat_9_13_io_out_r_load_store;
  wire                pe_mat_9_13_io_out_r_df_is_ws;
  wire                pe_mat_9_13_io_out_r_stall;
  wire       [15:0]   pe_mat_9_13_io_out_c_data;
  wire                pe_mat_9_13_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_9_14_io_out_r_data;
  wire                pe_mat_9_14_io_out_r_load_store;
  wire                pe_mat_9_14_io_out_r_df_is_ws;
  wire                pe_mat_9_14_io_out_r_stall;
  wire       [15:0]   pe_mat_9_14_io_out_c_data;
  wire                pe_mat_9_14_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_9_15_io_out_r_data;
  wire                pe_mat_9_15_io_out_r_load_store;
  wire                pe_mat_9_15_io_out_r_df_is_ws;
  wire                pe_mat_9_15_io_out_r_stall;
  wire       [15:0]   pe_mat_9_15_io_out_c_data;
  wire                pe_mat_9_15_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_10_0_io_out_r_data;
  wire                pe_mat_10_0_io_out_r_load_store;
  wire                pe_mat_10_0_io_out_r_df_is_ws;
  wire                pe_mat_10_0_io_out_r_stall;
  wire       [15:0]   pe_mat_10_0_io_out_c_data;
  wire                pe_mat_10_0_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_10_1_io_out_r_data;
  wire                pe_mat_10_1_io_out_r_load_store;
  wire                pe_mat_10_1_io_out_r_df_is_ws;
  wire                pe_mat_10_1_io_out_r_stall;
  wire       [15:0]   pe_mat_10_1_io_out_c_data;
  wire                pe_mat_10_1_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_10_2_io_out_r_data;
  wire                pe_mat_10_2_io_out_r_load_store;
  wire                pe_mat_10_2_io_out_r_df_is_ws;
  wire                pe_mat_10_2_io_out_r_stall;
  wire       [15:0]   pe_mat_10_2_io_out_c_data;
  wire                pe_mat_10_2_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_10_3_io_out_r_data;
  wire                pe_mat_10_3_io_out_r_load_store;
  wire                pe_mat_10_3_io_out_r_df_is_ws;
  wire                pe_mat_10_3_io_out_r_stall;
  wire       [15:0]   pe_mat_10_3_io_out_c_data;
  wire                pe_mat_10_3_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_10_4_io_out_r_data;
  wire                pe_mat_10_4_io_out_r_load_store;
  wire                pe_mat_10_4_io_out_r_df_is_ws;
  wire                pe_mat_10_4_io_out_r_stall;
  wire       [15:0]   pe_mat_10_4_io_out_c_data;
  wire                pe_mat_10_4_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_10_5_io_out_r_data;
  wire                pe_mat_10_5_io_out_r_load_store;
  wire                pe_mat_10_5_io_out_r_df_is_ws;
  wire                pe_mat_10_5_io_out_r_stall;
  wire       [15:0]   pe_mat_10_5_io_out_c_data;
  wire                pe_mat_10_5_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_10_6_io_out_r_data;
  wire                pe_mat_10_6_io_out_r_load_store;
  wire                pe_mat_10_6_io_out_r_df_is_ws;
  wire                pe_mat_10_6_io_out_r_stall;
  wire       [15:0]   pe_mat_10_6_io_out_c_data;
  wire                pe_mat_10_6_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_10_7_io_out_r_data;
  wire                pe_mat_10_7_io_out_r_load_store;
  wire                pe_mat_10_7_io_out_r_df_is_ws;
  wire                pe_mat_10_7_io_out_r_stall;
  wire       [15:0]   pe_mat_10_7_io_out_c_data;
  wire                pe_mat_10_7_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_10_8_io_out_r_data;
  wire                pe_mat_10_8_io_out_r_load_store;
  wire                pe_mat_10_8_io_out_r_df_is_ws;
  wire                pe_mat_10_8_io_out_r_stall;
  wire       [15:0]   pe_mat_10_8_io_out_c_data;
  wire                pe_mat_10_8_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_10_9_io_out_r_data;
  wire                pe_mat_10_9_io_out_r_load_store;
  wire                pe_mat_10_9_io_out_r_df_is_ws;
  wire                pe_mat_10_9_io_out_r_stall;
  wire       [15:0]   pe_mat_10_9_io_out_c_data;
  wire                pe_mat_10_9_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_10_10_io_out_r_data;
  wire                pe_mat_10_10_io_out_r_load_store;
  wire                pe_mat_10_10_io_out_r_df_is_ws;
  wire                pe_mat_10_10_io_out_r_stall;
  wire       [15:0]   pe_mat_10_10_io_out_c_data;
  wire                pe_mat_10_10_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_10_11_io_out_r_data;
  wire                pe_mat_10_11_io_out_r_load_store;
  wire                pe_mat_10_11_io_out_r_df_is_ws;
  wire                pe_mat_10_11_io_out_r_stall;
  wire       [15:0]   pe_mat_10_11_io_out_c_data;
  wire                pe_mat_10_11_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_10_12_io_out_r_data;
  wire                pe_mat_10_12_io_out_r_load_store;
  wire                pe_mat_10_12_io_out_r_df_is_ws;
  wire                pe_mat_10_12_io_out_r_stall;
  wire       [15:0]   pe_mat_10_12_io_out_c_data;
  wire                pe_mat_10_12_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_10_13_io_out_r_data;
  wire                pe_mat_10_13_io_out_r_load_store;
  wire                pe_mat_10_13_io_out_r_df_is_ws;
  wire                pe_mat_10_13_io_out_r_stall;
  wire       [15:0]   pe_mat_10_13_io_out_c_data;
  wire                pe_mat_10_13_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_10_14_io_out_r_data;
  wire                pe_mat_10_14_io_out_r_load_store;
  wire                pe_mat_10_14_io_out_r_df_is_ws;
  wire                pe_mat_10_14_io_out_r_stall;
  wire       [15:0]   pe_mat_10_14_io_out_c_data;
  wire                pe_mat_10_14_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_10_15_io_out_r_data;
  wire                pe_mat_10_15_io_out_r_load_store;
  wire                pe_mat_10_15_io_out_r_df_is_ws;
  wire                pe_mat_10_15_io_out_r_stall;
  wire       [15:0]   pe_mat_10_15_io_out_c_data;
  wire                pe_mat_10_15_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_11_0_io_out_r_data;
  wire                pe_mat_11_0_io_out_r_load_store;
  wire                pe_mat_11_0_io_out_r_df_is_ws;
  wire                pe_mat_11_0_io_out_r_stall;
  wire       [15:0]   pe_mat_11_0_io_out_c_data;
  wire                pe_mat_11_0_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_11_1_io_out_r_data;
  wire                pe_mat_11_1_io_out_r_load_store;
  wire                pe_mat_11_1_io_out_r_df_is_ws;
  wire                pe_mat_11_1_io_out_r_stall;
  wire       [15:0]   pe_mat_11_1_io_out_c_data;
  wire                pe_mat_11_1_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_11_2_io_out_r_data;
  wire                pe_mat_11_2_io_out_r_load_store;
  wire                pe_mat_11_2_io_out_r_df_is_ws;
  wire                pe_mat_11_2_io_out_r_stall;
  wire       [15:0]   pe_mat_11_2_io_out_c_data;
  wire                pe_mat_11_2_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_11_3_io_out_r_data;
  wire                pe_mat_11_3_io_out_r_load_store;
  wire                pe_mat_11_3_io_out_r_df_is_ws;
  wire                pe_mat_11_3_io_out_r_stall;
  wire       [15:0]   pe_mat_11_3_io_out_c_data;
  wire                pe_mat_11_3_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_11_4_io_out_r_data;
  wire                pe_mat_11_4_io_out_r_load_store;
  wire                pe_mat_11_4_io_out_r_df_is_ws;
  wire                pe_mat_11_4_io_out_r_stall;
  wire       [15:0]   pe_mat_11_4_io_out_c_data;
  wire                pe_mat_11_4_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_11_5_io_out_r_data;
  wire                pe_mat_11_5_io_out_r_load_store;
  wire                pe_mat_11_5_io_out_r_df_is_ws;
  wire                pe_mat_11_5_io_out_r_stall;
  wire       [15:0]   pe_mat_11_5_io_out_c_data;
  wire                pe_mat_11_5_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_11_6_io_out_r_data;
  wire                pe_mat_11_6_io_out_r_load_store;
  wire                pe_mat_11_6_io_out_r_df_is_ws;
  wire                pe_mat_11_6_io_out_r_stall;
  wire       [15:0]   pe_mat_11_6_io_out_c_data;
  wire                pe_mat_11_6_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_11_7_io_out_r_data;
  wire                pe_mat_11_7_io_out_r_load_store;
  wire                pe_mat_11_7_io_out_r_df_is_ws;
  wire                pe_mat_11_7_io_out_r_stall;
  wire       [15:0]   pe_mat_11_7_io_out_c_data;
  wire                pe_mat_11_7_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_11_8_io_out_r_data;
  wire                pe_mat_11_8_io_out_r_load_store;
  wire                pe_mat_11_8_io_out_r_df_is_ws;
  wire                pe_mat_11_8_io_out_r_stall;
  wire       [15:0]   pe_mat_11_8_io_out_c_data;
  wire                pe_mat_11_8_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_11_9_io_out_r_data;
  wire                pe_mat_11_9_io_out_r_load_store;
  wire                pe_mat_11_9_io_out_r_df_is_ws;
  wire                pe_mat_11_9_io_out_r_stall;
  wire       [15:0]   pe_mat_11_9_io_out_c_data;
  wire                pe_mat_11_9_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_11_10_io_out_r_data;
  wire                pe_mat_11_10_io_out_r_load_store;
  wire                pe_mat_11_10_io_out_r_df_is_ws;
  wire                pe_mat_11_10_io_out_r_stall;
  wire       [15:0]   pe_mat_11_10_io_out_c_data;
  wire                pe_mat_11_10_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_11_11_io_out_r_data;
  wire                pe_mat_11_11_io_out_r_load_store;
  wire                pe_mat_11_11_io_out_r_df_is_ws;
  wire                pe_mat_11_11_io_out_r_stall;
  wire       [15:0]   pe_mat_11_11_io_out_c_data;
  wire                pe_mat_11_11_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_11_12_io_out_r_data;
  wire                pe_mat_11_12_io_out_r_load_store;
  wire                pe_mat_11_12_io_out_r_df_is_ws;
  wire                pe_mat_11_12_io_out_r_stall;
  wire       [15:0]   pe_mat_11_12_io_out_c_data;
  wire                pe_mat_11_12_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_11_13_io_out_r_data;
  wire                pe_mat_11_13_io_out_r_load_store;
  wire                pe_mat_11_13_io_out_r_df_is_ws;
  wire                pe_mat_11_13_io_out_r_stall;
  wire       [15:0]   pe_mat_11_13_io_out_c_data;
  wire                pe_mat_11_13_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_11_14_io_out_r_data;
  wire                pe_mat_11_14_io_out_r_load_store;
  wire                pe_mat_11_14_io_out_r_df_is_ws;
  wire                pe_mat_11_14_io_out_r_stall;
  wire       [15:0]   pe_mat_11_14_io_out_c_data;
  wire                pe_mat_11_14_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_11_15_io_out_r_data;
  wire                pe_mat_11_15_io_out_r_load_store;
  wire                pe_mat_11_15_io_out_r_df_is_ws;
  wire                pe_mat_11_15_io_out_r_stall;
  wire       [15:0]   pe_mat_11_15_io_out_c_data;
  wire                pe_mat_11_15_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_12_0_io_out_r_data;
  wire                pe_mat_12_0_io_out_r_load_store;
  wire                pe_mat_12_0_io_out_r_df_is_ws;
  wire                pe_mat_12_0_io_out_r_stall;
  wire       [15:0]   pe_mat_12_0_io_out_c_data;
  wire                pe_mat_12_0_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_12_1_io_out_r_data;
  wire                pe_mat_12_1_io_out_r_load_store;
  wire                pe_mat_12_1_io_out_r_df_is_ws;
  wire                pe_mat_12_1_io_out_r_stall;
  wire       [15:0]   pe_mat_12_1_io_out_c_data;
  wire                pe_mat_12_1_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_12_2_io_out_r_data;
  wire                pe_mat_12_2_io_out_r_load_store;
  wire                pe_mat_12_2_io_out_r_df_is_ws;
  wire                pe_mat_12_2_io_out_r_stall;
  wire       [15:0]   pe_mat_12_2_io_out_c_data;
  wire                pe_mat_12_2_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_12_3_io_out_r_data;
  wire                pe_mat_12_3_io_out_r_load_store;
  wire                pe_mat_12_3_io_out_r_df_is_ws;
  wire                pe_mat_12_3_io_out_r_stall;
  wire       [15:0]   pe_mat_12_3_io_out_c_data;
  wire                pe_mat_12_3_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_12_4_io_out_r_data;
  wire                pe_mat_12_4_io_out_r_load_store;
  wire                pe_mat_12_4_io_out_r_df_is_ws;
  wire                pe_mat_12_4_io_out_r_stall;
  wire       [15:0]   pe_mat_12_4_io_out_c_data;
  wire                pe_mat_12_4_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_12_5_io_out_r_data;
  wire                pe_mat_12_5_io_out_r_load_store;
  wire                pe_mat_12_5_io_out_r_df_is_ws;
  wire                pe_mat_12_5_io_out_r_stall;
  wire       [15:0]   pe_mat_12_5_io_out_c_data;
  wire                pe_mat_12_5_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_12_6_io_out_r_data;
  wire                pe_mat_12_6_io_out_r_load_store;
  wire                pe_mat_12_6_io_out_r_df_is_ws;
  wire                pe_mat_12_6_io_out_r_stall;
  wire       [15:0]   pe_mat_12_6_io_out_c_data;
  wire                pe_mat_12_6_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_12_7_io_out_r_data;
  wire                pe_mat_12_7_io_out_r_load_store;
  wire                pe_mat_12_7_io_out_r_df_is_ws;
  wire                pe_mat_12_7_io_out_r_stall;
  wire       [15:0]   pe_mat_12_7_io_out_c_data;
  wire                pe_mat_12_7_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_12_8_io_out_r_data;
  wire                pe_mat_12_8_io_out_r_load_store;
  wire                pe_mat_12_8_io_out_r_df_is_ws;
  wire                pe_mat_12_8_io_out_r_stall;
  wire       [15:0]   pe_mat_12_8_io_out_c_data;
  wire                pe_mat_12_8_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_12_9_io_out_r_data;
  wire                pe_mat_12_9_io_out_r_load_store;
  wire                pe_mat_12_9_io_out_r_df_is_ws;
  wire                pe_mat_12_9_io_out_r_stall;
  wire       [15:0]   pe_mat_12_9_io_out_c_data;
  wire                pe_mat_12_9_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_12_10_io_out_r_data;
  wire                pe_mat_12_10_io_out_r_load_store;
  wire                pe_mat_12_10_io_out_r_df_is_ws;
  wire                pe_mat_12_10_io_out_r_stall;
  wire       [15:0]   pe_mat_12_10_io_out_c_data;
  wire                pe_mat_12_10_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_12_11_io_out_r_data;
  wire                pe_mat_12_11_io_out_r_load_store;
  wire                pe_mat_12_11_io_out_r_df_is_ws;
  wire                pe_mat_12_11_io_out_r_stall;
  wire       [15:0]   pe_mat_12_11_io_out_c_data;
  wire                pe_mat_12_11_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_12_12_io_out_r_data;
  wire                pe_mat_12_12_io_out_r_load_store;
  wire                pe_mat_12_12_io_out_r_df_is_ws;
  wire                pe_mat_12_12_io_out_r_stall;
  wire       [15:0]   pe_mat_12_12_io_out_c_data;
  wire                pe_mat_12_12_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_12_13_io_out_r_data;
  wire                pe_mat_12_13_io_out_r_load_store;
  wire                pe_mat_12_13_io_out_r_df_is_ws;
  wire                pe_mat_12_13_io_out_r_stall;
  wire       [15:0]   pe_mat_12_13_io_out_c_data;
  wire                pe_mat_12_13_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_12_14_io_out_r_data;
  wire                pe_mat_12_14_io_out_r_load_store;
  wire                pe_mat_12_14_io_out_r_df_is_ws;
  wire                pe_mat_12_14_io_out_r_stall;
  wire       [15:0]   pe_mat_12_14_io_out_c_data;
  wire                pe_mat_12_14_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_12_15_io_out_r_data;
  wire                pe_mat_12_15_io_out_r_load_store;
  wire                pe_mat_12_15_io_out_r_df_is_ws;
  wire                pe_mat_12_15_io_out_r_stall;
  wire       [15:0]   pe_mat_12_15_io_out_c_data;
  wire                pe_mat_12_15_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_13_0_io_out_r_data;
  wire                pe_mat_13_0_io_out_r_load_store;
  wire                pe_mat_13_0_io_out_r_df_is_ws;
  wire                pe_mat_13_0_io_out_r_stall;
  wire       [15:0]   pe_mat_13_0_io_out_c_data;
  wire                pe_mat_13_0_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_13_1_io_out_r_data;
  wire                pe_mat_13_1_io_out_r_load_store;
  wire                pe_mat_13_1_io_out_r_df_is_ws;
  wire                pe_mat_13_1_io_out_r_stall;
  wire       [15:0]   pe_mat_13_1_io_out_c_data;
  wire                pe_mat_13_1_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_13_2_io_out_r_data;
  wire                pe_mat_13_2_io_out_r_load_store;
  wire                pe_mat_13_2_io_out_r_df_is_ws;
  wire                pe_mat_13_2_io_out_r_stall;
  wire       [15:0]   pe_mat_13_2_io_out_c_data;
  wire                pe_mat_13_2_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_13_3_io_out_r_data;
  wire                pe_mat_13_3_io_out_r_load_store;
  wire                pe_mat_13_3_io_out_r_df_is_ws;
  wire                pe_mat_13_3_io_out_r_stall;
  wire       [15:0]   pe_mat_13_3_io_out_c_data;
  wire                pe_mat_13_3_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_13_4_io_out_r_data;
  wire                pe_mat_13_4_io_out_r_load_store;
  wire                pe_mat_13_4_io_out_r_df_is_ws;
  wire                pe_mat_13_4_io_out_r_stall;
  wire       [15:0]   pe_mat_13_4_io_out_c_data;
  wire                pe_mat_13_4_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_13_5_io_out_r_data;
  wire                pe_mat_13_5_io_out_r_load_store;
  wire                pe_mat_13_5_io_out_r_df_is_ws;
  wire                pe_mat_13_5_io_out_r_stall;
  wire       [15:0]   pe_mat_13_5_io_out_c_data;
  wire                pe_mat_13_5_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_13_6_io_out_r_data;
  wire                pe_mat_13_6_io_out_r_load_store;
  wire                pe_mat_13_6_io_out_r_df_is_ws;
  wire                pe_mat_13_6_io_out_r_stall;
  wire       [15:0]   pe_mat_13_6_io_out_c_data;
  wire                pe_mat_13_6_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_13_7_io_out_r_data;
  wire                pe_mat_13_7_io_out_r_load_store;
  wire                pe_mat_13_7_io_out_r_df_is_ws;
  wire                pe_mat_13_7_io_out_r_stall;
  wire       [15:0]   pe_mat_13_7_io_out_c_data;
  wire                pe_mat_13_7_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_13_8_io_out_r_data;
  wire                pe_mat_13_8_io_out_r_load_store;
  wire                pe_mat_13_8_io_out_r_df_is_ws;
  wire                pe_mat_13_8_io_out_r_stall;
  wire       [15:0]   pe_mat_13_8_io_out_c_data;
  wire                pe_mat_13_8_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_13_9_io_out_r_data;
  wire                pe_mat_13_9_io_out_r_load_store;
  wire                pe_mat_13_9_io_out_r_df_is_ws;
  wire                pe_mat_13_9_io_out_r_stall;
  wire       [15:0]   pe_mat_13_9_io_out_c_data;
  wire                pe_mat_13_9_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_13_10_io_out_r_data;
  wire                pe_mat_13_10_io_out_r_load_store;
  wire                pe_mat_13_10_io_out_r_df_is_ws;
  wire                pe_mat_13_10_io_out_r_stall;
  wire       [15:0]   pe_mat_13_10_io_out_c_data;
  wire                pe_mat_13_10_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_13_11_io_out_r_data;
  wire                pe_mat_13_11_io_out_r_load_store;
  wire                pe_mat_13_11_io_out_r_df_is_ws;
  wire                pe_mat_13_11_io_out_r_stall;
  wire       [15:0]   pe_mat_13_11_io_out_c_data;
  wire                pe_mat_13_11_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_13_12_io_out_r_data;
  wire                pe_mat_13_12_io_out_r_load_store;
  wire                pe_mat_13_12_io_out_r_df_is_ws;
  wire                pe_mat_13_12_io_out_r_stall;
  wire       [15:0]   pe_mat_13_12_io_out_c_data;
  wire                pe_mat_13_12_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_13_13_io_out_r_data;
  wire                pe_mat_13_13_io_out_r_load_store;
  wire                pe_mat_13_13_io_out_r_df_is_ws;
  wire                pe_mat_13_13_io_out_r_stall;
  wire       [15:0]   pe_mat_13_13_io_out_c_data;
  wire                pe_mat_13_13_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_13_14_io_out_r_data;
  wire                pe_mat_13_14_io_out_r_load_store;
  wire                pe_mat_13_14_io_out_r_df_is_ws;
  wire                pe_mat_13_14_io_out_r_stall;
  wire       [15:0]   pe_mat_13_14_io_out_c_data;
  wire                pe_mat_13_14_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_13_15_io_out_r_data;
  wire                pe_mat_13_15_io_out_r_load_store;
  wire                pe_mat_13_15_io_out_r_df_is_ws;
  wire                pe_mat_13_15_io_out_r_stall;
  wire       [15:0]   pe_mat_13_15_io_out_c_data;
  wire                pe_mat_13_15_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_14_0_io_out_r_data;
  wire                pe_mat_14_0_io_out_r_load_store;
  wire                pe_mat_14_0_io_out_r_df_is_ws;
  wire                pe_mat_14_0_io_out_r_stall;
  wire       [15:0]   pe_mat_14_0_io_out_c_data;
  wire                pe_mat_14_0_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_14_1_io_out_r_data;
  wire                pe_mat_14_1_io_out_r_load_store;
  wire                pe_mat_14_1_io_out_r_df_is_ws;
  wire                pe_mat_14_1_io_out_r_stall;
  wire       [15:0]   pe_mat_14_1_io_out_c_data;
  wire                pe_mat_14_1_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_14_2_io_out_r_data;
  wire                pe_mat_14_2_io_out_r_load_store;
  wire                pe_mat_14_2_io_out_r_df_is_ws;
  wire                pe_mat_14_2_io_out_r_stall;
  wire       [15:0]   pe_mat_14_2_io_out_c_data;
  wire                pe_mat_14_2_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_14_3_io_out_r_data;
  wire                pe_mat_14_3_io_out_r_load_store;
  wire                pe_mat_14_3_io_out_r_df_is_ws;
  wire                pe_mat_14_3_io_out_r_stall;
  wire       [15:0]   pe_mat_14_3_io_out_c_data;
  wire                pe_mat_14_3_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_14_4_io_out_r_data;
  wire                pe_mat_14_4_io_out_r_load_store;
  wire                pe_mat_14_4_io_out_r_df_is_ws;
  wire                pe_mat_14_4_io_out_r_stall;
  wire       [15:0]   pe_mat_14_4_io_out_c_data;
  wire                pe_mat_14_4_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_14_5_io_out_r_data;
  wire                pe_mat_14_5_io_out_r_load_store;
  wire                pe_mat_14_5_io_out_r_df_is_ws;
  wire                pe_mat_14_5_io_out_r_stall;
  wire       [15:0]   pe_mat_14_5_io_out_c_data;
  wire                pe_mat_14_5_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_14_6_io_out_r_data;
  wire                pe_mat_14_6_io_out_r_load_store;
  wire                pe_mat_14_6_io_out_r_df_is_ws;
  wire                pe_mat_14_6_io_out_r_stall;
  wire       [15:0]   pe_mat_14_6_io_out_c_data;
  wire                pe_mat_14_6_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_14_7_io_out_r_data;
  wire                pe_mat_14_7_io_out_r_load_store;
  wire                pe_mat_14_7_io_out_r_df_is_ws;
  wire                pe_mat_14_7_io_out_r_stall;
  wire       [15:0]   pe_mat_14_7_io_out_c_data;
  wire                pe_mat_14_7_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_14_8_io_out_r_data;
  wire                pe_mat_14_8_io_out_r_load_store;
  wire                pe_mat_14_8_io_out_r_df_is_ws;
  wire                pe_mat_14_8_io_out_r_stall;
  wire       [15:0]   pe_mat_14_8_io_out_c_data;
  wire                pe_mat_14_8_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_14_9_io_out_r_data;
  wire                pe_mat_14_9_io_out_r_load_store;
  wire                pe_mat_14_9_io_out_r_df_is_ws;
  wire                pe_mat_14_9_io_out_r_stall;
  wire       [15:0]   pe_mat_14_9_io_out_c_data;
  wire                pe_mat_14_9_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_14_10_io_out_r_data;
  wire                pe_mat_14_10_io_out_r_load_store;
  wire                pe_mat_14_10_io_out_r_df_is_ws;
  wire                pe_mat_14_10_io_out_r_stall;
  wire       [15:0]   pe_mat_14_10_io_out_c_data;
  wire                pe_mat_14_10_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_14_11_io_out_r_data;
  wire                pe_mat_14_11_io_out_r_load_store;
  wire                pe_mat_14_11_io_out_r_df_is_ws;
  wire                pe_mat_14_11_io_out_r_stall;
  wire       [15:0]   pe_mat_14_11_io_out_c_data;
  wire                pe_mat_14_11_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_14_12_io_out_r_data;
  wire                pe_mat_14_12_io_out_r_load_store;
  wire                pe_mat_14_12_io_out_r_df_is_ws;
  wire                pe_mat_14_12_io_out_r_stall;
  wire       [15:0]   pe_mat_14_12_io_out_c_data;
  wire                pe_mat_14_12_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_14_13_io_out_r_data;
  wire                pe_mat_14_13_io_out_r_load_store;
  wire                pe_mat_14_13_io_out_r_df_is_ws;
  wire                pe_mat_14_13_io_out_r_stall;
  wire       [15:0]   pe_mat_14_13_io_out_c_data;
  wire                pe_mat_14_13_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_14_14_io_out_r_data;
  wire                pe_mat_14_14_io_out_r_load_store;
  wire                pe_mat_14_14_io_out_r_df_is_ws;
  wire                pe_mat_14_14_io_out_r_stall;
  wire       [15:0]   pe_mat_14_14_io_out_c_data;
  wire                pe_mat_14_14_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_14_15_io_out_r_data;
  wire                pe_mat_14_15_io_out_r_load_store;
  wire                pe_mat_14_15_io_out_r_df_is_ws;
  wire                pe_mat_14_15_io_out_r_stall;
  wire       [15:0]   pe_mat_14_15_io_out_c_data;
  wire                pe_mat_14_15_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_15_0_io_out_r_data;
  wire                pe_mat_15_0_io_out_r_load_store;
  wire                pe_mat_15_0_io_out_r_df_is_ws;
  wire                pe_mat_15_0_io_out_r_stall;
  wire       [15:0]   pe_mat_15_0_io_out_c_data;
  wire                pe_mat_15_0_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_15_1_io_out_r_data;
  wire                pe_mat_15_1_io_out_r_load_store;
  wire                pe_mat_15_1_io_out_r_df_is_ws;
  wire                pe_mat_15_1_io_out_r_stall;
  wire       [15:0]   pe_mat_15_1_io_out_c_data;
  wire                pe_mat_15_1_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_15_2_io_out_r_data;
  wire                pe_mat_15_2_io_out_r_load_store;
  wire                pe_mat_15_2_io_out_r_df_is_ws;
  wire                pe_mat_15_2_io_out_r_stall;
  wire       [15:0]   pe_mat_15_2_io_out_c_data;
  wire                pe_mat_15_2_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_15_3_io_out_r_data;
  wire                pe_mat_15_3_io_out_r_load_store;
  wire                pe_mat_15_3_io_out_r_df_is_ws;
  wire                pe_mat_15_3_io_out_r_stall;
  wire       [15:0]   pe_mat_15_3_io_out_c_data;
  wire                pe_mat_15_3_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_15_4_io_out_r_data;
  wire                pe_mat_15_4_io_out_r_load_store;
  wire                pe_mat_15_4_io_out_r_df_is_ws;
  wire                pe_mat_15_4_io_out_r_stall;
  wire       [15:0]   pe_mat_15_4_io_out_c_data;
  wire                pe_mat_15_4_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_15_5_io_out_r_data;
  wire                pe_mat_15_5_io_out_r_load_store;
  wire                pe_mat_15_5_io_out_r_df_is_ws;
  wire                pe_mat_15_5_io_out_r_stall;
  wire       [15:0]   pe_mat_15_5_io_out_c_data;
  wire                pe_mat_15_5_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_15_6_io_out_r_data;
  wire                pe_mat_15_6_io_out_r_load_store;
  wire                pe_mat_15_6_io_out_r_df_is_ws;
  wire                pe_mat_15_6_io_out_r_stall;
  wire       [15:0]   pe_mat_15_6_io_out_c_data;
  wire                pe_mat_15_6_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_15_7_io_out_r_data;
  wire                pe_mat_15_7_io_out_r_load_store;
  wire                pe_mat_15_7_io_out_r_df_is_ws;
  wire                pe_mat_15_7_io_out_r_stall;
  wire       [15:0]   pe_mat_15_7_io_out_c_data;
  wire                pe_mat_15_7_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_15_8_io_out_r_data;
  wire                pe_mat_15_8_io_out_r_load_store;
  wire                pe_mat_15_8_io_out_r_df_is_ws;
  wire                pe_mat_15_8_io_out_r_stall;
  wire       [15:0]   pe_mat_15_8_io_out_c_data;
  wire                pe_mat_15_8_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_15_9_io_out_r_data;
  wire                pe_mat_15_9_io_out_r_load_store;
  wire                pe_mat_15_9_io_out_r_df_is_ws;
  wire                pe_mat_15_9_io_out_r_stall;
  wire       [15:0]   pe_mat_15_9_io_out_c_data;
  wire                pe_mat_15_9_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_15_10_io_out_r_data;
  wire                pe_mat_15_10_io_out_r_load_store;
  wire                pe_mat_15_10_io_out_r_df_is_ws;
  wire                pe_mat_15_10_io_out_r_stall;
  wire       [15:0]   pe_mat_15_10_io_out_c_data;
  wire                pe_mat_15_10_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_15_11_io_out_r_data;
  wire                pe_mat_15_11_io_out_r_load_store;
  wire                pe_mat_15_11_io_out_r_df_is_ws;
  wire                pe_mat_15_11_io_out_r_stall;
  wire       [15:0]   pe_mat_15_11_io_out_c_data;
  wire                pe_mat_15_11_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_15_12_io_out_r_data;
  wire                pe_mat_15_12_io_out_r_load_store;
  wire                pe_mat_15_12_io_out_r_df_is_ws;
  wire                pe_mat_15_12_io_out_r_stall;
  wire       [15:0]   pe_mat_15_12_io_out_c_data;
  wire                pe_mat_15_12_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_15_13_io_out_r_data;
  wire                pe_mat_15_13_io_out_r_load_store;
  wire                pe_mat_15_13_io_out_r_df_is_ws;
  wire                pe_mat_15_13_io_out_r_stall;
  wire       [15:0]   pe_mat_15_13_io_out_c_data;
  wire                pe_mat_15_13_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_15_14_io_out_r_data;
  wire                pe_mat_15_14_io_out_r_load_store;
  wire                pe_mat_15_14_io_out_r_df_is_ws;
  wire                pe_mat_15_14_io_out_r_stall;
  wire       [15:0]   pe_mat_15_14_io_out_c_data;
  wire                pe_mat_15_14_io_out_c_is_stationary;
  wire       [15:0]   pe_mat_15_15_io_out_r_data;
  wire                pe_mat_15_15_io_out_r_load_store;
  wire                pe_mat_15_15_io_out_r_df_is_ws;
  wire                pe_mat_15_15_io_out_r_stall;
  wire       [15:0]   pe_mat_15_15_io_out_c_data;
  wire                pe_mat_15_15_io_out_c_is_stationary;

  PEWSOS_255 pe_mat_0_0 (
    .io_in_r_data           (io_in_r_0_data[15:0]             ), //i
    .io_in_r_load_store     (io_in_r_0_load_store             ), //i
    .io_in_r_df_is_ws       (io_in_r_0_df_is_ws               ), //i
    .io_in_r_stall          (io_in_r_0_stall                  ), //i
    .io_out_r_data          (pe_mat_0_0_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_0_0_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_0_0_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_0_0_io_out_r_stall        ), //o
    .io_in_c_data           (io_in_c_0_data[15:0]             ), //i
    .io_in_c_is_stationary  (io_in_c_0_is_stationary          ), //i
    .io_out_c_data          (pe_mat_0_0_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_0_0_io_out_c_is_stationary), //o
    .clk                    (clk                              ), //i
    .reset                  (reset                            )  //i
  );
  PEWSOS_255 pe_mat_0_1 (
    .io_in_r_data           (pe_mat_0_0_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pe_mat_0_0_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pe_mat_0_0_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pe_mat_0_0_io_out_r_stall        ), //i
    .io_out_r_data          (pe_mat_0_1_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_0_1_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_0_1_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_0_1_io_out_r_stall        ), //o
    .io_in_c_data           (io_in_c_1_data[15:0]             ), //i
    .io_in_c_is_stationary  (io_in_c_1_is_stationary          ), //i
    .io_out_c_data          (pe_mat_0_1_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_0_1_io_out_c_is_stationary), //o
    .clk                    (clk                              ), //i
    .reset                  (reset                            )  //i
  );
  PEWSOS_255 pe_mat_0_2 (
    .io_in_r_data           (pe_mat_0_1_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pe_mat_0_1_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pe_mat_0_1_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pe_mat_0_1_io_out_r_stall        ), //i
    .io_out_r_data          (pe_mat_0_2_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_0_2_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_0_2_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_0_2_io_out_r_stall        ), //o
    .io_in_c_data           (io_in_c_2_data[15:0]             ), //i
    .io_in_c_is_stationary  (io_in_c_2_is_stationary          ), //i
    .io_out_c_data          (pe_mat_0_2_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_0_2_io_out_c_is_stationary), //o
    .clk                    (clk                              ), //i
    .reset                  (reset                            )  //i
  );
  PEWSOS_255 pe_mat_0_3 (
    .io_in_r_data           (pe_mat_0_2_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pe_mat_0_2_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pe_mat_0_2_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pe_mat_0_2_io_out_r_stall        ), //i
    .io_out_r_data          (pe_mat_0_3_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_0_3_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_0_3_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_0_3_io_out_r_stall        ), //o
    .io_in_c_data           (io_in_c_3_data[15:0]             ), //i
    .io_in_c_is_stationary  (io_in_c_3_is_stationary          ), //i
    .io_out_c_data          (pe_mat_0_3_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_0_3_io_out_c_is_stationary), //o
    .clk                    (clk                              ), //i
    .reset                  (reset                            )  //i
  );
  PEWSOS_255 pe_mat_0_4 (
    .io_in_r_data           (pe_mat_0_3_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pe_mat_0_3_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pe_mat_0_3_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pe_mat_0_3_io_out_r_stall        ), //i
    .io_out_r_data          (pe_mat_0_4_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_0_4_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_0_4_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_0_4_io_out_r_stall        ), //o
    .io_in_c_data           (io_in_c_4_data[15:0]             ), //i
    .io_in_c_is_stationary  (io_in_c_4_is_stationary          ), //i
    .io_out_c_data          (pe_mat_0_4_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_0_4_io_out_c_is_stationary), //o
    .clk                    (clk                              ), //i
    .reset                  (reset                            )  //i
  );
  PEWSOS_255 pe_mat_0_5 (
    .io_in_r_data           (pe_mat_0_4_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pe_mat_0_4_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pe_mat_0_4_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pe_mat_0_4_io_out_r_stall        ), //i
    .io_out_r_data          (pe_mat_0_5_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_0_5_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_0_5_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_0_5_io_out_r_stall        ), //o
    .io_in_c_data           (io_in_c_5_data[15:0]             ), //i
    .io_in_c_is_stationary  (io_in_c_5_is_stationary          ), //i
    .io_out_c_data          (pe_mat_0_5_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_0_5_io_out_c_is_stationary), //o
    .clk                    (clk                              ), //i
    .reset                  (reset                            )  //i
  );
  PEWSOS_255 pe_mat_0_6 (
    .io_in_r_data           (pe_mat_0_5_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pe_mat_0_5_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pe_mat_0_5_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pe_mat_0_5_io_out_r_stall        ), //i
    .io_out_r_data          (pe_mat_0_6_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_0_6_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_0_6_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_0_6_io_out_r_stall        ), //o
    .io_in_c_data           (io_in_c_6_data[15:0]             ), //i
    .io_in_c_is_stationary  (io_in_c_6_is_stationary          ), //i
    .io_out_c_data          (pe_mat_0_6_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_0_6_io_out_c_is_stationary), //o
    .clk                    (clk                              ), //i
    .reset                  (reset                            )  //i
  );
  PEWSOS_255 pe_mat_0_7 (
    .io_in_r_data           (pe_mat_0_6_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pe_mat_0_6_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pe_mat_0_6_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pe_mat_0_6_io_out_r_stall        ), //i
    .io_out_r_data          (pe_mat_0_7_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_0_7_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_0_7_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_0_7_io_out_r_stall        ), //o
    .io_in_c_data           (io_in_c_7_data[15:0]             ), //i
    .io_in_c_is_stationary  (io_in_c_7_is_stationary          ), //i
    .io_out_c_data          (pe_mat_0_7_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_0_7_io_out_c_is_stationary), //o
    .clk                    (clk                              ), //i
    .reset                  (reset                            )  //i
  );
  PEWSOS_255 pe_mat_0_8 (
    .io_in_r_data           (pe_mat_0_7_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pe_mat_0_7_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pe_mat_0_7_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pe_mat_0_7_io_out_r_stall        ), //i
    .io_out_r_data          (pe_mat_0_8_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_0_8_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_0_8_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_0_8_io_out_r_stall        ), //o
    .io_in_c_data           (io_in_c_8_data[15:0]             ), //i
    .io_in_c_is_stationary  (io_in_c_8_is_stationary          ), //i
    .io_out_c_data          (pe_mat_0_8_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_0_8_io_out_c_is_stationary), //o
    .clk                    (clk                              ), //i
    .reset                  (reset                            )  //i
  );
  PEWSOS_255 pe_mat_0_9 (
    .io_in_r_data           (pe_mat_0_8_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pe_mat_0_8_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pe_mat_0_8_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pe_mat_0_8_io_out_r_stall        ), //i
    .io_out_r_data          (pe_mat_0_9_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_0_9_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_0_9_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_0_9_io_out_r_stall        ), //o
    .io_in_c_data           (io_in_c_9_data[15:0]             ), //i
    .io_in_c_is_stationary  (io_in_c_9_is_stationary          ), //i
    .io_out_c_data          (pe_mat_0_9_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_0_9_io_out_c_is_stationary), //o
    .clk                    (clk                              ), //i
    .reset                  (reset                            )  //i
  );
  PEWSOS_255 pe_mat_0_10 (
    .io_in_r_data           (pe_mat_0_9_io_out_r_data[15:0]    ), //i
    .io_in_r_load_store     (pe_mat_0_9_io_out_r_load_store    ), //i
    .io_in_r_df_is_ws       (pe_mat_0_9_io_out_r_df_is_ws      ), //i
    .io_in_r_stall          (pe_mat_0_9_io_out_r_stall         ), //i
    .io_out_r_data          (pe_mat_0_10_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_0_10_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_0_10_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_0_10_io_out_r_stall        ), //o
    .io_in_c_data           (io_in_c_10_data[15:0]             ), //i
    .io_in_c_is_stationary  (io_in_c_10_is_stationary          ), //i
    .io_out_c_data          (pe_mat_0_10_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_0_10_io_out_c_is_stationary), //o
    .clk                    (clk                               ), //i
    .reset                  (reset                             )  //i
  );
  PEWSOS_255 pe_mat_0_11 (
    .io_in_r_data           (pe_mat_0_10_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pe_mat_0_10_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pe_mat_0_10_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pe_mat_0_10_io_out_r_stall        ), //i
    .io_out_r_data          (pe_mat_0_11_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_0_11_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_0_11_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_0_11_io_out_r_stall        ), //o
    .io_in_c_data           (io_in_c_11_data[15:0]             ), //i
    .io_in_c_is_stationary  (io_in_c_11_is_stationary          ), //i
    .io_out_c_data          (pe_mat_0_11_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_0_11_io_out_c_is_stationary), //o
    .clk                    (clk                               ), //i
    .reset                  (reset                             )  //i
  );
  PEWSOS_255 pe_mat_0_12 (
    .io_in_r_data           (pe_mat_0_11_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pe_mat_0_11_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pe_mat_0_11_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pe_mat_0_11_io_out_r_stall        ), //i
    .io_out_r_data          (pe_mat_0_12_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_0_12_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_0_12_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_0_12_io_out_r_stall        ), //o
    .io_in_c_data           (io_in_c_12_data[15:0]             ), //i
    .io_in_c_is_stationary  (io_in_c_12_is_stationary          ), //i
    .io_out_c_data          (pe_mat_0_12_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_0_12_io_out_c_is_stationary), //o
    .clk                    (clk                               ), //i
    .reset                  (reset                             )  //i
  );
  PEWSOS_255 pe_mat_0_13 (
    .io_in_r_data           (pe_mat_0_12_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pe_mat_0_12_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pe_mat_0_12_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pe_mat_0_12_io_out_r_stall        ), //i
    .io_out_r_data          (pe_mat_0_13_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_0_13_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_0_13_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_0_13_io_out_r_stall        ), //o
    .io_in_c_data           (io_in_c_13_data[15:0]             ), //i
    .io_in_c_is_stationary  (io_in_c_13_is_stationary          ), //i
    .io_out_c_data          (pe_mat_0_13_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_0_13_io_out_c_is_stationary), //o
    .clk                    (clk                               ), //i
    .reset                  (reset                             )  //i
  );
  PEWSOS_255 pe_mat_0_14 (
    .io_in_r_data           (pe_mat_0_13_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pe_mat_0_13_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pe_mat_0_13_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pe_mat_0_13_io_out_r_stall        ), //i
    .io_out_r_data          (pe_mat_0_14_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_0_14_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_0_14_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_0_14_io_out_r_stall        ), //o
    .io_in_c_data           (io_in_c_14_data[15:0]             ), //i
    .io_in_c_is_stationary  (io_in_c_14_is_stationary          ), //i
    .io_out_c_data          (pe_mat_0_14_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_0_14_io_out_c_is_stationary), //o
    .clk                    (clk                               ), //i
    .reset                  (reset                             )  //i
  );
  PEWSOS_255 pe_mat_0_15 (
    .io_in_r_data           (pe_mat_0_14_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pe_mat_0_14_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pe_mat_0_14_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pe_mat_0_14_io_out_r_stall        ), //i
    .io_out_r_data          (pe_mat_0_15_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_0_15_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_0_15_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_0_15_io_out_r_stall        ), //o
    .io_in_c_data           (io_in_c_15_data[15:0]             ), //i
    .io_in_c_is_stationary  (io_in_c_15_is_stationary          ), //i
    .io_out_c_data          (pe_mat_0_15_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_0_15_io_out_c_is_stationary), //o
    .clk                    (clk                               ), //i
    .reset                  (reset                             )  //i
  );
  PEWSOS_255 pe_mat_1_0 (
    .io_in_r_data           (io_in_r_1_data[15:0]             ), //i
    .io_in_r_load_store     (io_in_r_1_load_store             ), //i
    .io_in_r_df_is_ws       (io_in_r_1_df_is_ws               ), //i
    .io_in_r_stall          (io_in_r_1_stall                  ), //i
    .io_out_r_data          (pe_mat_1_0_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_1_0_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_1_0_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_1_0_io_out_r_stall        ), //o
    .io_in_c_data           (pe_mat_0_0_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pe_mat_0_0_io_out_c_is_stationary), //i
    .io_out_c_data          (pe_mat_1_0_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_1_0_io_out_c_is_stationary), //o
    .clk                    (clk                              ), //i
    .reset                  (reset                            )  //i
  );
  PEWSOS_255 pe_mat_1_1 (
    .io_in_r_data           (pe_mat_1_0_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pe_mat_1_0_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pe_mat_1_0_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pe_mat_1_0_io_out_r_stall        ), //i
    .io_out_r_data          (pe_mat_1_1_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_1_1_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_1_1_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_1_1_io_out_r_stall        ), //o
    .io_in_c_data           (pe_mat_0_1_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pe_mat_0_1_io_out_c_is_stationary), //i
    .io_out_c_data          (pe_mat_1_1_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_1_1_io_out_c_is_stationary), //o
    .clk                    (clk                              ), //i
    .reset                  (reset                            )  //i
  );
  PEWSOS_255 pe_mat_1_2 (
    .io_in_r_data           (pe_mat_1_1_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pe_mat_1_1_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pe_mat_1_1_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pe_mat_1_1_io_out_r_stall        ), //i
    .io_out_r_data          (pe_mat_1_2_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_1_2_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_1_2_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_1_2_io_out_r_stall        ), //o
    .io_in_c_data           (pe_mat_0_2_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pe_mat_0_2_io_out_c_is_stationary), //i
    .io_out_c_data          (pe_mat_1_2_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_1_2_io_out_c_is_stationary), //o
    .clk                    (clk                              ), //i
    .reset                  (reset                            )  //i
  );
  PEWSOS_255 pe_mat_1_3 (
    .io_in_r_data           (pe_mat_1_2_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pe_mat_1_2_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pe_mat_1_2_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pe_mat_1_2_io_out_r_stall        ), //i
    .io_out_r_data          (pe_mat_1_3_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_1_3_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_1_3_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_1_3_io_out_r_stall        ), //o
    .io_in_c_data           (pe_mat_0_3_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pe_mat_0_3_io_out_c_is_stationary), //i
    .io_out_c_data          (pe_mat_1_3_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_1_3_io_out_c_is_stationary), //o
    .clk                    (clk                              ), //i
    .reset                  (reset                            )  //i
  );
  PEWSOS_255 pe_mat_1_4 (
    .io_in_r_data           (pe_mat_1_3_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pe_mat_1_3_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pe_mat_1_3_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pe_mat_1_3_io_out_r_stall        ), //i
    .io_out_r_data          (pe_mat_1_4_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_1_4_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_1_4_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_1_4_io_out_r_stall        ), //o
    .io_in_c_data           (pe_mat_0_4_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pe_mat_0_4_io_out_c_is_stationary), //i
    .io_out_c_data          (pe_mat_1_4_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_1_4_io_out_c_is_stationary), //o
    .clk                    (clk                              ), //i
    .reset                  (reset                            )  //i
  );
  PEWSOS_255 pe_mat_1_5 (
    .io_in_r_data           (pe_mat_1_4_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pe_mat_1_4_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pe_mat_1_4_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pe_mat_1_4_io_out_r_stall        ), //i
    .io_out_r_data          (pe_mat_1_5_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_1_5_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_1_5_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_1_5_io_out_r_stall        ), //o
    .io_in_c_data           (pe_mat_0_5_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pe_mat_0_5_io_out_c_is_stationary), //i
    .io_out_c_data          (pe_mat_1_5_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_1_5_io_out_c_is_stationary), //o
    .clk                    (clk                              ), //i
    .reset                  (reset                            )  //i
  );
  PEWSOS_255 pe_mat_1_6 (
    .io_in_r_data           (pe_mat_1_5_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pe_mat_1_5_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pe_mat_1_5_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pe_mat_1_5_io_out_r_stall        ), //i
    .io_out_r_data          (pe_mat_1_6_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_1_6_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_1_6_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_1_6_io_out_r_stall        ), //o
    .io_in_c_data           (pe_mat_0_6_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pe_mat_0_6_io_out_c_is_stationary), //i
    .io_out_c_data          (pe_mat_1_6_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_1_6_io_out_c_is_stationary), //o
    .clk                    (clk                              ), //i
    .reset                  (reset                            )  //i
  );
  PEWSOS_255 pe_mat_1_7 (
    .io_in_r_data           (pe_mat_1_6_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pe_mat_1_6_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pe_mat_1_6_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pe_mat_1_6_io_out_r_stall        ), //i
    .io_out_r_data          (pe_mat_1_7_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_1_7_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_1_7_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_1_7_io_out_r_stall        ), //o
    .io_in_c_data           (pe_mat_0_7_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pe_mat_0_7_io_out_c_is_stationary), //i
    .io_out_c_data          (pe_mat_1_7_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_1_7_io_out_c_is_stationary), //o
    .clk                    (clk                              ), //i
    .reset                  (reset                            )  //i
  );
  PEWSOS_255 pe_mat_1_8 (
    .io_in_r_data           (pe_mat_1_7_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pe_mat_1_7_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pe_mat_1_7_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pe_mat_1_7_io_out_r_stall        ), //i
    .io_out_r_data          (pe_mat_1_8_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_1_8_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_1_8_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_1_8_io_out_r_stall        ), //o
    .io_in_c_data           (pe_mat_0_8_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pe_mat_0_8_io_out_c_is_stationary), //i
    .io_out_c_data          (pe_mat_1_8_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_1_8_io_out_c_is_stationary), //o
    .clk                    (clk                              ), //i
    .reset                  (reset                            )  //i
  );
  PEWSOS_255 pe_mat_1_9 (
    .io_in_r_data           (pe_mat_1_8_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pe_mat_1_8_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pe_mat_1_8_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pe_mat_1_8_io_out_r_stall        ), //i
    .io_out_r_data          (pe_mat_1_9_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_1_9_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_1_9_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_1_9_io_out_r_stall        ), //o
    .io_in_c_data           (pe_mat_0_9_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pe_mat_0_9_io_out_c_is_stationary), //i
    .io_out_c_data          (pe_mat_1_9_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_1_9_io_out_c_is_stationary), //o
    .clk                    (clk                              ), //i
    .reset                  (reset                            )  //i
  );
  PEWSOS_255 pe_mat_1_10 (
    .io_in_r_data           (pe_mat_1_9_io_out_r_data[15:0]    ), //i
    .io_in_r_load_store     (pe_mat_1_9_io_out_r_load_store    ), //i
    .io_in_r_df_is_ws       (pe_mat_1_9_io_out_r_df_is_ws      ), //i
    .io_in_r_stall          (pe_mat_1_9_io_out_r_stall         ), //i
    .io_out_r_data          (pe_mat_1_10_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_1_10_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_1_10_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_1_10_io_out_r_stall        ), //o
    .io_in_c_data           (pe_mat_0_10_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pe_mat_0_10_io_out_c_is_stationary), //i
    .io_out_c_data          (pe_mat_1_10_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_1_10_io_out_c_is_stationary), //o
    .clk                    (clk                               ), //i
    .reset                  (reset                             )  //i
  );
  PEWSOS_255 pe_mat_1_11 (
    .io_in_r_data           (pe_mat_1_10_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pe_mat_1_10_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pe_mat_1_10_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pe_mat_1_10_io_out_r_stall        ), //i
    .io_out_r_data          (pe_mat_1_11_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_1_11_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_1_11_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_1_11_io_out_r_stall        ), //o
    .io_in_c_data           (pe_mat_0_11_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pe_mat_0_11_io_out_c_is_stationary), //i
    .io_out_c_data          (pe_mat_1_11_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_1_11_io_out_c_is_stationary), //o
    .clk                    (clk                               ), //i
    .reset                  (reset                             )  //i
  );
  PEWSOS_255 pe_mat_1_12 (
    .io_in_r_data           (pe_mat_1_11_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pe_mat_1_11_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pe_mat_1_11_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pe_mat_1_11_io_out_r_stall        ), //i
    .io_out_r_data          (pe_mat_1_12_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_1_12_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_1_12_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_1_12_io_out_r_stall        ), //o
    .io_in_c_data           (pe_mat_0_12_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pe_mat_0_12_io_out_c_is_stationary), //i
    .io_out_c_data          (pe_mat_1_12_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_1_12_io_out_c_is_stationary), //o
    .clk                    (clk                               ), //i
    .reset                  (reset                             )  //i
  );
  PEWSOS_255 pe_mat_1_13 (
    .io_in_r_data           (pe_mat_1_12_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pe_mat_1_12_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pe_mat_1_12_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pe_mat_1_12_io_out_r_stall        ), //i
    .io_out_r_data          (pe_mat_1_13_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_1_13_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_1_13_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_1_13_io_out_r_stall        ), //o
    .io_in_c_data           (pe_mat_0_13_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pe_mat_0_13_io_out_c_is_stationary), //i
    .io_out_c_data          (pe_mat_1_13_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_1_13_io_out_c_is_stationary), //o
    .clk                    (clk                               ), //i
    .reset                  (reset                             )  //i
  );
  PEWSOS_255 pe_mat_1_14 (
    .io_in_r_data           (pe_mat_1_13_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pe_mat_1_13_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pe_mat_1_13_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pe_mat_1_13_io_out_r_stall        ), //i
    .io_out_r_data          (pe_mat_1_14_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_1_14_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_1_14_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_1_14_io_out_r_stall        ), //o
    .io_in_c_data           (pe_mat_0_14_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pe_mat_0_14_io_out_c_is_stationary), //i
    .io_out_c_data          (pe_mat_1_14_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_1_14_io_out_c_is_stationary), //o
    .clk                    (clk                               ), //i
    .reset                  (reset                             )  //i
  );
  PEWSOS_255 pe_mat_1_15 (
    .io_in_r_data           (pe_mat_1_14_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pe_mat_1_14_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pe_mat_1_14_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pe_mat_1_14_io_out_r_stall        ), //i
    .io_out_r_data          (pe_mat_1_15_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_1_15_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_1_15_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_1_15_io_out_r_stall        ), //o
    .io_in_c_data           (pe_mat_0_15_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pe_mat_0_15_io_out_c_is_stationary), //i
    .io_out_c_data          (pe_mat_1_15_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_1_15_io_out_c_is_stationary), //o
    .clk                    (clk                               ), //i
    .reset                  (reset                             )  //i
  );
  PEWSOS_255 pe_mat_2_0 (
    .io_in_r_data           (io_in_r_2_data[15:0]             ), //i
    .io_in_r_load_store     (io_in_r_2_load_store             ), //i
    .io_in_r_df_is_ws       (io_in_r_2_df_is_ws               ), //i
    .io_in_r_stall          (io_in_r_2_stall                  ), //i
    .io_out_r_data          (pe_mat_2_0_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_2_0_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_2_0_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_2_0_io_out_r_stall        ), //o
    .io_in_c_data           (pe_mat_1_0_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pe_mat_1_0_io_out_c_is_stationary), //i
    .io_out_c_data          (pe_mat_2_0_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_2_0_io_out_c_is_stationary), //o
    .clk                    (clk                              ), //i
    .reset                  (reset                            )  //i
  );
  PEWSOS_255 pe_mat_2_1 (
    .io_in_r_data           (pe_mat_2_0_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pe_mat_2_0_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pe_mat_2_0_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pe_mat_2_0_io_out_r_stall        ), //i
    .io_out_r_data          (pe_mat_2_1_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_2_1_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_2_1_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_2_1_io_out_r_stall        ), //o
    .io_in_c_data           (pe_mat_1_1_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pe_mat_1_1_io_out_c_is_stationary), //i
    .io_out_c_data          (pe_mat_2_1_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_2_1_io_out_c_is_stationary), //o
    .clk                    (clk                              ), //i
    .reset                  (reset                            )  //i
  );
  PEWSOS_255 pe_mat_2_2 (
    .io_in_r_data           (pe_mat_2_1_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pe_mat_2_1_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pe_mat_2_1_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pe_mat_2_1_io_out_r_stall        ), //i
    .io_out_r_data          (pe_mat_2_2_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_2_2_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_2_2_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_2_2_io_out_r_stall        ), //o
    .io_in_c_data           (pe_mat_1_2_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pe_mat_1_2_io_out_c_is_stationary), //i
    .io_out_c_data          (pe_mat_2_2_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_2_2_io_out_c_is_stationary), //o
    .clk                    (clk                              ), //i
    .reset                  (reset                            )  //i
  );
  PEWSOS_255 pe_mat_2_3 (
    .io_in_r_data           (pe_mat_2_2_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pe_mat_2_2_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pe_mat_2_2_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pe_mat_2_2_io_out_r_stall        ), //i
    .io_out_r_data          (pe_mat_2_3_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_2_3_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_2_3_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_2_3_io_out_r_stall        ), //o
    .io_in_c_data           (pe_mat_1_3_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pe_mat_1_3_io_out_c_is_stationary), //i
    .io_out_c_data          (pe_mat_2_3_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_2_3_io_out_c_is_stationary), //o
    .clk                    (clk                              ), //i
    .reset                  (reset                            )  //i
  );
  PEWSOS_255 pe_mat_2_4 (
    .io_in_r_data           (pe_mat_2_3_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pe_mat_2_3_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pe_mat_2_3_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pe_mat_2_3_io_out_r_stall        ), //i
    .io_out_r_data          (pe_mat_2_4_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_2_4_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_2_4_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_2_4_io_out_r_stall        ), //o
    .io_in_c_data           (pe_mat_1_4_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pe_mat_1_4_io_out_c_is_stationary), //i
    .io_out_c_data          (pe_mat_2_4_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_2_4_io_out_c_is_stationary), //o
    .clk                    (clk                              ), //i
    .reset                  (reset                            )  //i
  );
  PEWSOS_255 pe_mat_2_5 (
    .io_in_r_data           (pe_mat_2_4_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pe_mat_2_4_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pe_mat_2_4_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pe_mat_2_4_io_out_r_stall        ), //i
    .io_out_r_data          (pe_mat_2_5_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_2_5_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_2_5_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_2_5_io_out_r_stall        ), //o
    .io_in_c_data           (pe_mat_1_5_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pe_mat_1_5_io_out_c_is_stationary), //i
    .io_out_c_data          (pe_mat_2_5_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_2_5_io_out_c_is_stationary), //o
    .clk                    (clk                              ), //i
    .reset                  (reset                            )  //i
  );
  PEWSOS_255 pe_mat_2_6 (
    .io_in_r_data           (pe_mat_2_5_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pe_mat_2_5_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pe_mat_2_5_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pe_mat_2_5_io_out_r_stall        ), //i
    .io_out_r_data          (pe_mat_2_6_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_2_6_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_2_6_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_2_6_io_out_r_stall        ), //o
    .io_in_c_data           (pe_mat_1_6_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pe_mat_1_6_io_out_c_is_stationary), //i
    .io_out_c_data          (pe_mat_2_6_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_2_6_io_out_c_is_stationary), //o
    .clk                    (clk                              ), //i
    .reset                  (reset                            )  //i
  );
  PEWSOS_255 pe_mat_2_7 (
    .io_in_r_data           (pe_mat_2_6_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pe_mat_2_6_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pe_mat_2_6_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pe_mat_2_6_io_out_r_stall        ), //i
    .io_out_r_data          (pe_mat_2_7_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_2_7_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_2_7_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_2_7_io_out_r_stall        ), //o
    .io_in_c_data           (pe_mat_1_7_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pe_mat_1_7_io_out_c_is_stationary), //i
    .io_out_c_data          (pe_mat_2_7_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_2_7_io_out_c_is_stationary), //o
    .clk                    (clk                              ), //i
    .reset                  (reset                            )  //i
  );
  PEWSOS_255 pe_mat_2_8 (
    .io_in_r_data           (pe_mat_2_7_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pe_mat_2_7_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pe_mat_2_7_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pe_mat_2_7_io_out_r_stall        ), //i
    .io_out_r_data          (pe_mat_2_8_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_2_8_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_2_8_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_2_8_io_out_r_stall        ), //o
    .io_in_c_data           (pe_mat_1_8_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pe_mat_1_8_io_out_c_is_stationary), //i
    .io_out_c_data          (pe_mat_2_8_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_2_8_io_out_c_is_stationary), //o
    .clk                    (clk                              ), //i
    .reset                  (reset                            )  //i
  );
  PEWSOS_255 pe_mat_2_9 (
    .io_in_r_data           (pe_mat_2_8_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pe_mat_2_8_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pe_mat_2_8_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pe_mat_2_8_io_out_r_stall        ), //i
    .io_out_r_data          (pe_mat_2_9_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_2_9_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_2_9_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_2_9_io_out_r_stall        ), //o
    .io_in_c_data           (pe_mat_1_9_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pe_mat_1_9_io_out_c_is_stationary), //i
    .io_out_c_data          (pe_mat_2_9_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_2_9_io_out_c_is_stationary), //o
    .clk                    (clk                              ), //i
    .reset                  (reset                            )  //i
  );
  PEWSOS_255 pe_mat_2_10 (
    .io_in_r_data           (pe_mat_2_9_io_out_r_data[15:0]    ), //i
    .io_in_r_load_store     (pe_mat_2_9_io_out_r_load_store    ), //i
    .io_in_r_df_is_ws       (pe_mat_2_9_io_out_r_df_is_ws      ), //i
    .io_in_r_stall          (pe_mat_2_9_io_out_r_stall         ), //i
    .io_out_r_data          (pe_mat_2_10_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_2_10_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_2_10_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_2_10_io_out_r_stall        ), //o
    .io_in_c_data           (pe_mat_1_10_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pe_mat_1_10_io_out_c_is_stationary), //i
    .io_out_c_data          (pe_mat_2_10_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_2_10_io_out_c_is_stationary), //o
    .clk                    (clk                               ), //i
    .reset                  (reset                             )  //i
  );
  PEWSOS_255 pe_mat_2_11 (
    .io_in_r_data           (pe_mat_2_10_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pe_mat_2_10_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pe_mat_2_10_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pe_mat_2_10_io_out_r_stall        ), //i
    .io_out_r_data          (pe_mat_2_11_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_2_11_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_2_11_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_2_11_io_out_r_stall        ), //o
    .io_in_c_data           (pe_mat_1_11_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pe_mat_1_11_io_out_c_is_stationary), //i
    .io_out_c_data          (pe_mat_2_11_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_2_11_io_out_c_is_stationary), //o
    .clk                    (clk                               ), //i
    .reset                  (reset                             )  //i
  );
  PEWSOS_255 pe_mat_2_12 (
    .io_in_r_data           (pe_mat_2_11_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pe_mat_2_11_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pe_mat_2_11_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pe_mat_2_11_io_out_r_stall        ), //i
    .io_out_r_data          (pe_mat_2_12_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_2_12_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_2_12_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_2_12_io_out_r_stall        ), //o
    .io_in_c_data           (pe_mat_1_12_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pe_mat_1_12_io_out_c_is_stationary), //i
    .io_out_c_data          (pe_mat_2_12_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_2_12_io_out_c_is_stationary), //o
    .clk                    (clk                               ), //i
    .reset                  (reset                             )  //i
  );
  PEWSOS_255 pe_mat_2_13 (
    .io_in_r_data           (pe_mat_2_12_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pe_mat_2_12_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pe_mat_2_12_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pe_mat_2_12_io_out_r_stall        ), //i
    .io_out_r_data          (pe_mat_2_13_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_2_13_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_2_13_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_2_13_io_out_r_stall        ), //o
    .io_in_c_data           (pe_mat_1_13_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pe_mat_1_13_io_out_c_is_stationary), //i
    .io_out_c_data          (pe_mat_2_13_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_2_13_io_out_c_is_stationary), //o
    .clk                    (clk                               ), //i
    .reset                  (reset                             )  //i
  );
  PEWSOS_255 pe_mat_2_14 (
    .io_in_r_data           (pe_mat_2_13_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pe_mat_2_13_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pe_mat_2_13_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pe_mat_2_13_io_out_r_stall        ), //i
    .io_out_r_data          (pe_mat_2_14_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_2_14_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_2_14_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_2_14_io_out_r_stall        ), //o
    .io_in_c_data           (pe_mat_1_14_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pe_mat_1_14_io_out_c_is_stationary), //i
    .io_out_c_data          (pe_mat_2_14_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_2_14_io_out_c_is_stationary), //o
    .clk                    (clk                               ), //i
    .reset                  (reset                             )  //i
  );
  PEWSOS_255 pe_mat_2_15 (
    .io_in_r_data           (pe_mat_2_14_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pe_mat_2_14_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pe_mat_2_14_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pe_mat_2_14_io_out_r_stall        ), //i
    .io_out_r_data          (pe_mat_2_15_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_2_15_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_2_15_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_2_15_io_out_r_stall        ), //o
    .io_in_c_data           (pe_mat_1_15_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pe_mat_1_15_io_out_c_is_stationary), //i
    .io_out_c_data          (pe_mat_2_15_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_2_15_io_out_c_is_stationary), //o
    .clk                    (clk                               ), //i
    .reset                  (reset                             )  //i
  );
  PEWSOS_255 pe_mat_3_0 (
    .io_in_r_data           (io_in_r_3_data[15:0]             ), //i
    .io_in_r_load_store     (io_in_r_3_load_store             ), //i
    .io_in_r_df_is_ws       (io_in_r_3_df_is_ws               ), //i
    .io_in_r_stall          (io_in_r_3_stall                  ), //i
    .io_out_r_data          (pe_mat_3_0_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_3_0_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_3_0_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_3_0_io_out_r_stall        ), //o
    .io_in_c_data           (pe_mat_2_0_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pe_mat_2_0_io_out_c_is_stationary), //i
    .io_out_c_data          (pe_mat_3_0_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_3_0_io_out_c_is_stationary), //o
    .clk                    (clk                              ), //i
    .reset                  (reset                            )  //i
  );
  PEWSOS_255 pe_mat_3_1 (
    .io_in_r_data           (pe_mat_3_0_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pe_mat_3_0_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pe_mat_3_0_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pe_mat_3_0_io_out_r_stall        ), //i
    .io_out_r_data          (pe_mat_3_1_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_3_1_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_3_1_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_3_1_io_out_r_stall        ), //o
    .io_in_c_data           (pe_mat_2_1_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pe_mat_2_1_io_out_c_is_stationary), //i
    .io_out_c_data          (pe_mat_3_1_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_3_1_io_out_c_is_stationary), //o
    .clk                    (clk                              ), //i
    .reset                  (reset                            )  //i
  );
  PEWSOS_255 pe_mat_3_2 (
    .io_in_r_data           (pe_mat_3_1_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pe_mat_3_1_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pe_mat_3_1_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pe_mat_3_1_io_out_r_stall        ), //i
    .io_out_r_data          (pe_mat_3_2_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_3_2_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_3_2_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_3_2_io_out_r_stall        ), //o
    .io_in_c_data           (pe_mat_2_2_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pe_mat_2_2_io_out_c_is_stationary), //i
    .io_out_c_data          (pe_mat_3_2_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_3_2_io_out_c_is_stationary), //o
    .clk                    (clk                              ), //i
    .reset                  (reset                            )  //i
  );
  PEWSOS_255 pe_mat_3_3 (
    .io_in_r_data           (pe_mat_3_2_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pe_mat_3_2_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pe_mat_3_2_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pe_mat_3_2_io_out_r_stall        ), //i
    .io_out_r_data          (pe_mat_3_3_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_3_3_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_3_3_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_3_3_io_out_r_stall        ), //o
    .io_in_c_data           (pe_mat_2_3_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pe_mat_2_3_io_out_c_is_stationary), //i
    .io_out_c_data          (pe_mat_3_3_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_3_3_io_out_c_is_stationary), //o
    .clk                    (clk                              ), //i
    .reset                  (reset                            )  //i
  );
  PEWSOS_255 pe_mat_3_4 (
    .io_in_r_data           (pe_mat_3_3_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pe_mat_3_3_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pe_mat_3_3_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pe_mat_3_3_io_out_r_stall        ), //i
    .io_out_r_data          (pe_mat_3_4_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_3_4_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_3_4_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_3_4_io_out_r_stall        ), //o
    .io_in_c_data           (pe_mat_2_4_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pe_mat_2_4_io_out_c_is_stationary), //i
    .io_out_c_data          (pe_mat_3_4_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_3_4_io_out_c_is_stationary), //o
    .clk                    (clk                              ), //i
    .reset                  (reset                            )  //i
  );
  PEWSOS_255 pe_mat_3_5 (
    .io_in_r_data           (pe_mat_3_4_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pe_mat_3_4_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pe_mat_3_4_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pe_mat_3_4_io_out_r_stall        ), //i
    .io_out_r_data          (pe_mat_3_5_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_3_5_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_3_5_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_3_5_io_out_r_stall        ), //o
    .io_in_c_data           (pe_mat_2_5_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pe_mat_2_5_io_out_c_is_stationary), //i
    .io_out_c_data          (pe_mat_3_5_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_3_5_io_out_c_is_stationary), //o
    .clk                    (clk                              ), //i
    .reset                  (reset                            )  //i
  );
  PEWSOS_255 pe_mat_3_6 (
    .io_in_r_data           (pe_mat_3_5_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pe_mat_3_5_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pe_mat_3_5_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pe_mat_3_5_io_out_r_stall        ), //i
    .io_out_r_data          (pe_mat_3_6_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_3_6_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_3_6_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_3_6_io_out_r_stall        ), //o
    .io_in_c_data           (pe_mat_2_6_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pe_mat_2_6_io_out_c_is_stationary), //i
    .io_out_c_data          (pe_mat_3_6_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_3_6_io_out_c_is_stationary), //o
    .clk                    (clk                              ), //i
    .reset                  (reset                            )  //i
  );
  PEWSOS_255 pe_mat_3_7 (
    .io_in_r_data           (pe_mat_3_6_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pe_mat_3_6_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pe_mat_3_6_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pe_mat_3_6_io_out_r_stall        ), //i
    .io_out_r_data          (pe_mat_3_7_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_3_7_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_3_7_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_3_7_io_out_r_stall        ), //o
    .io_in_c_data           (pe_mat_2_7_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pe_mat_2_7_io_out_c_is_stationary), //i
    .io_out_c_data          (pe_mat_3_7_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_3_7_io_out_c_is_stationary), //o
    .clk                    (clk                              ), //i
    .reset                  (reset                            )  //i
  );
  PEWSOS_255 pe_mat_3_8 (
    .io_in_r_data           (pe_mat_3_7_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pe_mat_3_7_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pe_mat_3_7_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pe_mat_3_7_io_out_r_stall        ), //i
    .io_out_r_data          (pe_mat_3_8_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_3_8_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_3_8_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_3_8_io_out_r_stall        ), //o
    .io_in_c_data           (pe_mat_2_8_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pe_mat_2_8_io_out_c_is_stationary), //i
    .io_out_c_data          (pe_mat_3_8_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_3_8_io_out_c_is_stationary), //o
    .clk                    (clk                              ), //i
    .reset                  (reset                            )  //i
  );
  PEWSOS_255 pe_mat_3_9 (
    .io_in_r_data           (pe_mat_3_8_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pe_mat_3_8_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pe_mat_3_8_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pe_mat_3_8_io_out_r_stall        ), //i
    .io_out_r_data          (pe_mat_3_9_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_3_9_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_3_9_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_3_9_io_out_r_stall        ), //o
    .io_in_c_data           (pe_mat_2_9_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pe_mat_2_9_io_out_c_is_stationary), //i
    .io_out_c_data          (pe_mat_3_9_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_3_9_io_out_c_is_stationary), //o
    .clk                    (clk                              ), //i
    .reset                  (reset                            )  //i
  );
  PEWSOS_255 pe_mat_3_10 (
    .io_in_r_data           (pe_mat_3_9_io_out_r_data[15:0]    ), //i
    .io_in_r_load_store     (pe_mat_3_9_io_out_r_load_store    ), //i
    .io_in_r_df_is_ws       (pe_mat_3_9_io_out_r_df_is_ws      ), //i
    .io_in_r_stall          (pe_mat_3_9_io_out_r_stall         ), //i
    .io_out_r_data          (pe_mat_3_10_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_3_10_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_3_10_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_3_10_io_out_r_stall        ), //o
    .io_in_c_data           (pe_mat_2_10_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pe_mat_2_10_io_out_c_is_stationary), //i
    .io_out_c_data          (pe_mat_3_10_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_3_10_io_out_c_is_stationary), //o
    .clk                    (clk                               ), //i
    .reset                  (reset                             )  //i
  );
  PEWSOS_255 pe_mat_3_11 (
    .io_in_r_data           (pe_mat_3_10_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pe_mat_3_10_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pe_mat_3_10_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pe_mat_3_10_io_out_r_stall        ), //i
    .io_out_r_data          (pe_mat_3_11_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_3_11_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_3_11_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_3_11_io_out_r_stall        ), //o
    .io_in_c_data           (pe_mat_2_11_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pe_mat_2_11_io_out_c_is_stationary), //i
    .io_out_c_data          (pe_mat_3_11_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_3_11_io_out_c_is_stationary), //o
    .clk                    (clk                               ), //i
    .reset                  (reset                             )  //i
  );
  PEWSOS_255 pe_mat_3_12 (
    .io_in_r_data           (pe_mat_3_11_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pe_mat_3_11_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pe_mat_3_11_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pe_mat_3_11_io_out_r_stall        ), //i
    .io_out_r_data          (pe_mat_3_12_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_3_12_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_3_12_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_3_12_io_out_r_stall        ), //o
    .io_in_c_data           (pe_mat_2_12_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pe_mat_2_12_io_out_c_is_stationary), //i
    .io_out_c_data          (pe_mat_3_12_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_3_12_io_out_c_is_stationary), //o
    .clk                    (clk                               ), //i
    .reset                  (reset                             )  //i
  );
  PEWSOS_255 pe_mat_3_13 (
    .io_in_r_data           (pe_mat_3_12_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pe_mat_3_12_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pe_mat_3_12_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pe_mat_3_12_io_out_r_stall        ), //i
    .io_out_r_data          (pe_mat_3_13_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_3_13_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_3_13_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_3_13_io_out_r_stall        ), //o
    .io_in_c_data           (pe_mat_2_13_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pe_mat_2_13_io_out_c_is_stationary), //i
    .io_out_c_data          (pe_mat_3_13_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_3_13_io_out_c_is_stationary), //o
    .clk                    (clk                               ), //i
    .reset                  (reset                             )  //i
  );
  PEWSOS_255 pe_mat_3_14 (
    .io_in_r_data           (pe_mat_3_13_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pe_mat_3_13_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pe_mat_3_13_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pe_mat_3_13_io_out_r_stall        ), //i
    .io_out_r_data          (pe_mat_3_14_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_3_14_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_3_14_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_3_14_io_out_r_stall        ), //o
    .io_in_c_data           (pe_mat_2_14_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pe_mat_2_14_io_out_c_is_stationary), //i
    .io_out_c_data          (pe_mat_3_14_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_3_14_io_out_c_is_stationary), //o
    .clk                    (clk                               ), //i
    .reset                  (reset                             )  //i
  );
  PEWSOS_255 pe_mat_3_15 (
    .io_in_r_data           (pe_mat_3_14_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pe_mat_3_14_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pe_mat_3_14_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pe_mat_3_14_io_out_r_stall        ), //i
    .io_out_r_data          (pe_mat_3_15_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_3_15_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_3_15_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_3_15_io_out_r_stall        ), //o
    .io_in_c_data           (pe_mat_2_15_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pe_mat_2_15_io_out_c_is_stationary), //i
    .io_out_c_data          (pe_mat_3_15_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_3_15_io_out_c_is_stationary), //o
    .clk                    (clk                               ), //i
    .reset                  (reset                             )  //i
  );
  PEWSOS_255 pe_mat_4_0 (
    .io_in_r_data           (io_in_r_4_data[15:0]             ), //i
    .io_in_r_load_store     (io_in_r_4_load_store             ), //i
    .io_in_r_df_is_ws       (io_in_r_4_df_is_ws               ), //i
    .io_in_r_stall          (io_in_r_4_stall                  ), //i
    .io_out_r_data          (pe_mat_4_0_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_4_0_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_4_0_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_4_0_io_out_r_stall        ), //o
    .io_in_c_data           (pe_mat_3_0_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pe_mat_3_0_io_out_c_is_stationary), //i
    .io_out_c_data          (pe_mat_4_0_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_4_0_io_out_c_is_stationary), //o
    .clk                    (clk                              ), //i
    .reset                  (reset                            )  //i
  );
  PEWSOS_255 pe_mat_4_1 (
    .io_in_r_data           (pe_mat_4_0_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pe_mat_4_0_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pe_mat_4_0_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pe_mat_4_0_io_out_r_stall        ), //i
    .io_out_r_data          (pe_mat_4_1_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_4_1_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_4_1_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_4_1_io_out_r_stall        ), //o
    .io_in_c_data           (pe_mat_3_1_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pe_mat_3_1_io_out_c_is_stationary), //i
    .io_out_c_data          (pe_mat_4_1_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_4_1_io_out_c_is_stationary), //o
    .clk                    (clk                              ), //i
    .reset                  (reset                            )  //i
  );
  PEWSOS_255 pe_mat_4_2 (
    .io_in_r_data           (pe_mat_4_1_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pe_mat_4_1_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pe_mat_4_1_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pe_mat_4_1_io_out_r_stall        ), //i
    .io_out_r_data          (pe_mat_4_2_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_4_2_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_4_2_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_4_2_io_out_r_stall        ), //o
    .io_in_c_data           (pe_mat_3_2_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pe_mat_3_2_io_out_c_is_stationary), //i
    .io_out_c_data          (pe_mat_4_2_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_4_2_io_out_c_is_stationary), //o
    .clk                    (clk                              ), //i
    .reset                  (reset                            )  //i
  );
  PEWSOS_255 pe_mat_4_3 (
    .io_in_r_data           (pe_mat_4_2_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pe_mat_4_2_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pe_mat_4_2_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pe_mat_4_2_io_out_r_stall        ), //i
    .io_out_r_data          (pe_mat_4_3_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_4_3_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_4_3_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_4_3_io_out_r_stall        ), //o
    .io_in_c_data           (pe_mat_3_3_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pe_mat_3_3_io_out_c_is_stationary), //i
    .io_out_c_data          (pe_mat_4_3_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_4_3_io_out_c_is_stationary), //o
    .clk                    (clk                              ), //i
    .reset                  (reset                            )  //i
  );
  PEWSOS_255 pe_mat_4_4 (
    .io_in_r_data           (pe_mat_4_3_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pe_mat_4_3_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pe_mat_4_3_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pe_mat_4_3_io_out_r_stall        ), //i
    .io_out_r_data          (pe_mat_4_4_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_4_4_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_4_4_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_4_4_io_out_r_stall        ), //o
    .io_in_c_data           (pe_mat_3_4_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pe_mat_3_4_io_out_c_is_stationary), //i
    .io_out_c_data          (pe_mat_4_4_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_4_4_io_out_c_is_stationary), //o
    .clk                    (clk                              ), //i
    .reset                  (reset                            )  //i
  );
  PEWSOS_255 pe_mat_4_5 (
    .io_in_r_data           (pe_mat_4_4_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pe_mat_4_4_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pe_mat_4_4_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pe_mat_4_4_io_out_r_stall        ), //i
    .io_out_r_data          (pe_mat_4_5_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_4_5_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_4_5_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_4_5_io_out_r_stall        ), //o
    .io_in_c_data           (pe_mat_3_5_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pe_mat_3_5_io_out_c_is_stationary), //i
    .io_out_c_data          (pe_mat_4_5_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_4_5_io_out_c_is_stationary), //o
    .clk                    (clk                              ), //i
    .reset                  (reset                            )  //i
  );
  PEWSOS_255 pe_mat_4_6 (
    .io_in_r_data           (pe_mat_4_5_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pe_mat_4_5_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pe_mat_4_5_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pe_mat_4_5_io_out_r_stall        ), //i
    .io_out_r_data          (pe_mat_4_6_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_4_6_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_4_6_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_4_6_io_out_r_stall        ), //o
    .io_in_c_data           (pe_mat_3_6_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pe_mat_3_6_io_out_c_is_stationary), //i
    .io_out_c_data          (pe_mat_4_6_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_4_6_io_out_c_is_stationary), //o
    .clk                    (clk                              ), //i
    .reset                  (reset                            )  //i
  );
  PEWSOS_255 pe_mat_4_7 (
    .io_in_r_data           (pe_mat_4_6_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pe_mat_4_6_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pe_mat_4_6_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pe_mat_4_6_io_out_r_stall        ), //i
    .io_out_r_data          (pe_mat_4_7_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_4_7_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_4_7_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_4_7_io_out_r_stall        ), //o
    .io_in_c_data           (pe_mat_3_7_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pe_mat_3_7_io_out_c_is_stationary), //i
    .io_out_c_data          (pe_mat_4_7_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_4_7_io_out_c_is_stationary), //o
    .clk                    (clk                              ), //i
    .reset                  (reset                            )  //i
  );
  PEWSOS_255 pe_mat_4_8 (
    .io_in_r_data           (pe_mat_4_7_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pe_mat_4_7_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pe_mat_4_7_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pe_mat_4_7_io_out_r_stall        ), //i
    .io_out_r_data          (pe_mat_4_8_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_4_8_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_4_8_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_4_8_io_out_r_stall        ), //o
    .io_in_c_data           (pe_mat_3_8_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pe_mat_3_8_io_out_c_is_stationary), //i
    .io_out_c_data          (pe_mat_4_8_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_4_8_io_out_c_is_stationary), //o
    .clk                    (clk                              ), //i
    .reset                  (reset                            )  //i
  );
  PEWSOS_255 pe_mat_4_9 (
    .io_in_r_data           (pe_mat_4_8_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pe_mat_4_8_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pe_mat_4_8_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pe_mat_4_8_io_out_r_stall        ), //i
    .io_out_r_data          (pe_mat_4_9_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_4_9_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_4_9_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_4_9_io_out_r_stall        ), //o
    .io_in_c_data           (pe_mat_3_9_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pe_mat_3_9_io_out_c_is_stationary), //i
    .io_out_c_data          (pe_mat_4_9_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_4_9_io_out_c_is_stationary), //o
    .clk                    (clk                              ), //i
    .reset                  (reset                            )  //i
  );
  PEWSOS_255 pe_mat_4_10 (
    .io_in_r_data           (pe_mat_4_9_io_out_r_data[15:0]    ), //i
    .io_in_r_load_store     (pe_mat_4_9_io_out_r_load_store    ), //i
    .io_in_r_df_is_ws       (pe_mat_4_9_io_out_r_df_is_ws      ), //i
    .io_in_r_stall          (pe_mat_4_9_io_out_r_stall         ), //i
    .io_out_r_data          (pe_mat_4_10_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_4_10_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_4_10_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_4_10_io_out_r_stall        ), //o
    .io_in_c_data           (pe_mat_3_10_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pe_mat_3_10_io_out_c_is_stationary), //i
    .io_out_c_data          (pe_mat_4_10_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_4_10_io_out_c_is_stationary), //o
    .clk                    (clk                               ), //i
    .reset                  (reset                             )  //i
  );
  PEWSOS_255 pe_mat_4_11 (
    .io_in_r_data           (pe_mat_4_10_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pe_mat_4_10_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pe_mat_4_10_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pe_mat_4_10_io_out_r_stall        ), //i
    .io_out_r_data          (pe_mat_4_11_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_4_11_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_4_11_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_4_11_io_out_r_stall        ), //o
    .io_in_c_data           (pe_mat_3_11_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pe_mat_3_11_io_out_c_is_stationary), //i
    .io_out_c_data          (pe_mat_4_11_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_4_11_io_out_c_is_stationary), //o
    .clk                    (clk                               ), //i
    .reset                  (reset                             )  //i
  );
  PEWSOS_255 pe_mat_4_12 (
    .io_in_r_data           (pe_mat_4_11_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pe_mat_4_11_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pe_mat_4_11_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pe_mat_4_11_io_out_r_stall        ), //i
    .io_out_r_data          (pe_mat_4_12_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_4_12_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_4_12_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_4_12_io_out_r_stall        ), //o
    .io_in_c_data           (pe_mat_3_12_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pe_mat_3_12_io_out_c_is_stationary), //i
    .io_out_c_data          (pe_mat_4_12_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_4_12_io_out_c_is_stationary), //o
    .clk                    (clk                               ), //i
    .reset                  (reset                             )  //i
  );
  PEWSOS_255 pe_mat_4_13 (
    .io_in_r_data           (pe_mat_4_12_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pe_mat_4_12_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pe_mat_4_12_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pe_mat_4_12_io_out_r_stall        ), //i
    .io_out_r_data          (pe_mat_4_13_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_4_13_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_4_13_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_4_13_io_out_r_stall        ), //o
    .io_in_c_data           (pe_mat_3_13_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pe_mat_3_13_io_out_c_is_stationary), //i
    .io_out_c_data          (pe_mat_4_13_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_4_13_io_out_c_is_stationary), //o
    .clk                    (clk                               ), //i
    .reset                  (reset                             )  //i
  );
  PEWSOS_255 pe_mat_4_14 (
    .io_in_r_data           (pe_mat_4_13_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pe_mat_4_13_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pe_mat_4_13_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pe_mat_4_13_io_out_r_stall        ), //i
    .io_out_r_data          (pe_mat_4_14_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_4_14_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_4_14_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_4_14_io_out_r_stall        ), //o
    .io_in_c_data           (pe_mat_3_14_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pe_mat_3_14_io_out_c_is_stationary), //i
    .io_out_c_data          (pe_mat_4_14_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_4_14_io_out_c_is_stationary), //o
    .clk                    (clk                               ), //i
    .reset                  (reset                             )  //i
  );
  PEWSOS_255 pe_mat_4_15 (
    .io_in_r_data           (pe_mat_4_14_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pe_mat_4_14_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pe_mat_4_14_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pe_mat_4_14_io_out_r_stall        ), //i
    .io_out_r_data          (pe_mat_4_15_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_4_15_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_4_15_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_4_15_io_out_r_stall        ), //o
    .io_in_c_data           (pe_mat_3_15_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pe_mat_3_15_io_out_c_is_stationary), //i
    .io_out_c_data          (pe_mat_4_15_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_4_15_io_out_c_is_stationary), //o
    .clk                    (clk                               ), //i
    .reset                  (reset                             )  //i
  );
  PEWSOS_255 pe_mat_5_0 (
    .io_in_r_data           (io_in_r_5_data[15:0]             ), //i
    .io_in_r_load_store     (io_in_r_5_load_store             ), //i
    .io_in_r_df_is_ws       (io_in_r_5_df_is_ws               ), //i
    .io_in_r_stall          (io_in_r_5_stall                  ), //i
    .io_out_r_data          (pe_mat_5_0_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_5_0_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_5_0_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_5_0_io_out_r_stall        ), //o
    .io_in_c_data           (pe_mat_4_0_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pe_mat_4_0_io_out_c_is_stationary), //i
    .io_out_c_data          (pe_mat_5_0_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_5_0_io_out_c_is_stationary), //o
    .clk                    (clk                              ), //i
    .reset                  (reset                            )  //i
  );
  PEWSOS_255 pe_mat_5_1 (
    .io_in_r_data           (pe_mat_5_0_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pe_mat_5_0_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pe_mat_5_0_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pe_mat_5_0_io_out_r_stall        ), //i
    .io_out_r_data          (pe_mat_5_1_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_5_1_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_5_1_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_5_1_io_out_r_stall        ), //o
    .io_in_c_data           (pe_mat_4_1_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pe_mat_4_1_io_out_c_is_stationary), //i
    .io_out_c_data          (pe_mat_5_1_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_5_1_io_out_c_is_stationary), //o
    .clk                    (clk                              ), //i
    .reset                  (reset                            )  //i
  );
  PEWSOS_255 pe_mat_5_2 (
    .io_in_r_data           (pe_mat_5_1_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pe_mat_5_1_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pe_mat_5_1_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pe_mat_5_1_io_out_r_stall        ), //i
    .io_out_r_data          (pe_mat_5_2_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_5_2_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_5_2_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_5_2_io_out_r_stall        ), //o
    .io_in_c_data           (pe_mat_4_2_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pe_mat_4_2_io_out_c_is_stationary), //i
    .io_out_c_data          (pe_mat_5_2_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_5_2_io_out_c_is_stationary), //o
    .clk                    (clk                              ), //i
    .reset                  (reset                            )  //i
  );
  PEWSOS_255 pe_mat_5_3 (
    .io_in_r_data           (pe_mat_5_2_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pe_mat_5_2_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pe_mat_5_2_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pe_mat_5_2_io_out_r_stall        ), //i
    .io_out_r_data          (pe_mat_5_3_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_5_3_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_5_3_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_5_3_io_out_r_stall        ), //o
    .io_in_c_data           (pe_mat_4_3_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pe_mat_4_3_io_out_c_is_stationary), //i
    .io_out_c_data          (pe_mat_5_3_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_5_3_io_out_c_is_stationary), //o
    .clk                    (clk                              ), //i
    .reset                  (reset                            )  //i
  );
  PEWSOS_255 pe_mat_5_4 (
    .io_in_r_data           (pe_mat_5_3_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pe_mat_5_3_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pe_mat_5_3_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pe_mat_5_3_io_out_r_stall        ), //i
    .io_out_r_data          (pe_mat_5_4_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_5_4_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_5_4_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_5_4_io_out_r_stall        ), //o
    .io_in_c_data           (pe_mat_4_4_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pe_mat_4_4_io_out_c_is_stationary), //i
    .io_out_c_data          (pe_mat_5_4_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_5_4_io_out_c_is_stationary), //o
    .clk                    (clk                              ), //i
    .reset                  (reset                            )  //i
  );
  PEWSOS_255 pe_mat_5_5 (
    .io_in_r_data           (pe_mat_5_4_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pe_mat_5_4_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pe_mat_5_4_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pe_mat_5_4_io_out_r_stall        ), //i
    .io_out_r_data          (pe_mat_5_5_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_5_5_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_5_5_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_5_5_io_out_r_stall        ), //o
    .io_in_c_data           (pe_mat_4_5_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pe_mat_4_5_io_out_c_is_stationary), //i
    .io_out_c_data          (pe_mat_5_5_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_5_5_io_out_c_is_stationary), //o
    .clk                    (clk                              ), //i
    .reset                  (reset                            )  //i
  );
  PEWSOS_255 pe_mat_5_6 (
    .io_in_r_data           (pe_mat_5_5_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pe_mat_5_5_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pe_mat_5_5_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pe_mat_5_5_io_out_r_stall        ), //i
    .io_out_r_data          (pe_mat_5_6_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_5_6_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_5_6_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_5_6_io_out_r_stall        ), //o
    .io_in_c_data           (pe_mat_4_6_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pe_mat_4_6_io_out_c_is_stationary), //i
    .io_out_c_data          (pe_mat_5_6_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_5_6_io_out_c_is_stationary), //o
    .clk                    (clk                              ), //i
    .reset                  (reset                            )  //i
  );
  PEWSOS_255 pe_mat_5_7 (
    .io_in_r_data           (pe_mat_5_6_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pe_mat_5_6_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pe_mat_5_6_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pe_mat_5_6_io_out_r_stall        ), //i
    .io_out_r_data          (pe_mat_5_7_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_5_7_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_5_7_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_5_7_io_out_r_stall        ), //o
    .io_in_c_data           (pe_mat_4_7_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pe_mat_4_7_io_out_c_is_stationary), //i
    .io_out_c_data          (pe_mat_5_7_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_5_7_io_out_c_is_stationary), //o
    .clk                    (clk                              ), //i
    .reset                  (reset                            )  //i
  );
  PEWSOS_255 pe_mat_5_8 (
    .io_in_r_data           (pe_mat_5_7_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pe_mat_5_7_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pe_mat_5_7_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pe_mat_5_7_io_out_r_stall        ), //i
    .io_out_r_data          (pe_mat_5_8_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_5_8_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_5_8_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_5_8_io_out_r_stall        ), //o
    .io_in_c_data           (pe_mat_4_8_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pe_mat_4_8_io_out_c_is_stationary), //i
    .io_out_c_data          (pe_mat_5_8_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_5_8_io_out_c_is_stationary), //o
    .clk                    (clk                              ), //i
    .reset                  (reset                            )  //i
  );
  PEWSOS_255 pe_mat_5_9 (
    .io_in_r_data           (pe_mat_5_8_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pe_mat_5_8_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pe_mat_5_8_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pe_mat_5_8_io_out_r_stall        ), //i
    .io_out_r_data          (pe_mat_5_9_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_5_9_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_5_9_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_5_9_io_out_r_stall        ), //o
    .io_in_c_data           (pe_mat_4_9_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pe_mat_4_9_io_out_c_is_stationary), //i
    .io_out_c_data          (pe_mat_5_9_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_5_9_io_out_c_is_stationary), //o
    .clk                    (clk                              ), //i
    .reset                  (reset                            )  //i
  );
  PEWSOS_255 pe_mat_5_10 (
    .io_in_r_data           (pe_mat_5_9_io_out_r_data[15:0]    ), //i
    .io_in_r_load_store     (pe_mat_5_9_io_out_r_load_store    ), //i
    .io_in_r_df_is_ws       (pe_mat_5_9_io_out_r_df_is_ws      ), //i
    .io_in_r_stall          (pe_mat_5_9_io_out_r_stall         ), //i
    .io_out_r_data          (pe_mat_5_10_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_5_10_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_5_10_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_5_10_io_out_r_stall        ), //o
    .io_in_c_data           (pe_mat_4_10_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pe_mat_4_10_io_out_c_is_stationary), //i
    .io_out_c_data          (pe_mat_5_10_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_5_10_io_out_c_is_stationary), //o
    .clk                    (clk                               ), //i
    .reset                  (reset                             )  //i
  );
  PEWSOS_255 pe_mat_5_11 (
    .io_in_r_data           (pe_mat_5_10_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pe_mat_5_10_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pe_mat_5_10_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pe_mat_5_10_io_out_r_stall        ), //i
    .io_out_r_data          (pe_mat_5_11_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_5_11_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_5_11_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_5_11_io_out_r_stall        ), //o
    .io_in_c_data           (pe_mat_4_11_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pe_mat_4_11_io_out_c_is_stationary), //i
    .io_out_c_data          (pe_mat_5_11_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_5_11_io_out_c_is_stationary), //o
    .clk                    (clk                               ), //i
    .reset                  (reset                             )  //i
  );
  PEWSOS_255 pe_mat_5_12 (
    .io_in_r_data           (pe_mat_5_11_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pe_mat_5_11_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pe_mat_5_11_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pe_mat_5_11_io_out_r_stall        ), //i
    .io_out_r_data          (pe_mat_5_12_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_5_12_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_5_12_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_5_12_io_out_r_stall        ), //o
    .io_in_c_data           (pe_mat_4_12_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pe_mat_4_12_io_out_c_is_stationary), //i
    .io_out_c_data          (pe_mat_5_12_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_5_12_io_out_c_is_stationary), //o
    .clk                    (clk                               ), //i
    .reset                  (reset                             )  //i
  );
  PEWSOS_255 pe_mat_5_13 (
    .io_in_r_data           (pe_mat_5_12_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pe_mat_5_12_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pe_mat_5_12_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pe_mat_5_12_io_out_r_stall        ), //i
    .io_out_r_data          (pe_mat_5_13_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_5_13_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_5_13_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_5_13_io_out_r_stall        ), //o
    .io_in_c_data           (pe_mat_4_13_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pe_mat_4_13_io_out_c_is_stationary), //i
    .io_out_c_data          (pe_mat_5_13_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_5_13_io_out_c_is_stationary), //o
    .clk                    (clk                               ), //i
    .reset                  (reset                             )  //i
  );
  PEWSOS_255 pe_mat_5_14 (
    .io_in_r_data           (pe_mat_5_13_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pe_mat_5_13_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pe_mat_5_13_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pe_mat_5_13_io_out_r_stall        ), //i
    .io_out_r_data          (pe_mat_5_14_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_5_14_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_5_14_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_5_14_io_out_r_stall        ), //o
    .io_in_c_data           (pe_mat_4_14_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pe_mat_4_14_io_out_c_is_stationary), //i
    .io_out_c_data          (pe_mat_5_14_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_5_14_io_out_c_is_stationary), //o
    .clk                    (clk                               ), //i
    .reset                  (reset                             )  //i
  );
  PEWSOS_255 pe_mat_5_15 (
    .io_in_r_data           (pe_mat_5_14_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pe_mat_5_14_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pe_mat_5_14_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pe_mat_5_14_io_out_r_stall        ), //i
    .io_out_r_data          (pe_mat_5_15_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_5_15_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_5_15_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_5_15_io_out_r_stall        ), //o
    .io_in_c_data           (pe_mat_4_15_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pe_mat_4_15_io_out_c_is_stationary), //i
    .io_out_c_data          (pe_mat_5_15_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_5_15_io_out_c_is_stationary), //o
    .clk                    (clk                               ), //i
    .reset                  (reset                             )  //i
  );
  PEWSOS_255 pe_mat_6_0 (
    .io_in_r_data           (io_in_r_6_data[15:0]             ), //i
    .io_in_r_load_store     (io_in_r_6_load_store             ), //i
    .io_in_r_df_is_ws       (io_in_r_6_df_is_ws               ), //i
    .io_in_r_stall          (io_in_r_6_stall                  ), //i
    .io_out_r_data          (pe_mat_6_0_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_6_0_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_6_0_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_6_0_io_out_r_stall        ), //o
    .io_in_c_data           (pe_mat_5_0_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pe_mat_5_0_io_out_c_is_stationary), //i
    .io_out_c_data          (pe_mat_6_0_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_6_0_io_out_c_is_stationary), //o
    .clk                    (clk                              ), //i
    .reset                  (reset                            )  //i
  );
  PEWSOS_255 pe_mat_6_1 (
    .io_in_r_data           (pe_mat_6_0_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pe_mat_6_0_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pe_mat_6_0_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pe_mat_6_0_io_out_r_stall        ), //i
    .io_out_r_data          (pe_mat_6_1_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_6_1_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_6_1_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_6_1_io_out_r_stall        ), //o
    .io_in_c_data           (pe_mat_5_1_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pe_mat_5_1_io_out_c_is_stationary), //i
    .io_out_c_data          (pe_mat_6_1_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_6_1_io_out_c_is_stationary), //o
    .clk                    (clk                              ), //i
    .reset                  (reset                            )  //i
  );
  PEWSOS_255 pe_mat_6_2 (
    .io_in_r_data           (pe_mat_6_1_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pe_mat_6_1_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pe_mat_6_1_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pe_mat_6_1_io_out_r_stall        ), //i
    .io_out_r_data          (pe_mat_6_2_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_6_2_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_6_2_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_6_2_io_out_r_stall        ), //o
    .io_in_c_data           (pe_mat_5_2_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pe_mat_5_2_io_out_c_is_stationary), //i
    .io_out_c_data          (pe_mat_6_2_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_6_2_io_out_c_is_stationary), //o
    .clk                    (clk                              ), //i
    .reset                  (reset                            )  //i
  );
  PEWSOS_255 pe_mat_6_3 (
    .io_in_r_data           (pe_mat_6_2_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pe_mat_6_2_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pe_mat_6_2_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pe_mat_6_2_io_out_r_stall        ), //i
    .io_out_r_data          (pe_mat_6_3_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_6_3_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_6_3_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_6_3_io_out_r_stall        ), //o
    .io_in_c_data           (pe_mat_5_3_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pe_mat_5_3_io_out_c_is_stationary), //i
    .io_out_c_data          (pe_mat_6_3_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_6_3_io_out_c_is_stationary), //o
    .clk                    (clk                              ), //i
    .reset                  (reset                            )  //i
  );
  PEWSOS_255 pe_mat_6_4 (
    .io_in_r_data           (pe_mat_6_3_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pe_mat_6_3_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pe_mat_6_3_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pe_mat_6_3_io_out_r_stall        ), //i
    .io_out_r_data          (pe_mat_6_4_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_6_4_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_6_4_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_6_4_io_out_r_stall        ), //o
    .io_in_c_data           (pe_mat_5_4_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pe_mat_5_4_io_out_c_is_stationary), //i
    .io_out_c_data          (pe_mat_6_4_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_6_4_io_out_c_is_stationary), //o
    .clk                    (clk                              ), //i
    .reset                  (reset                            )  //i
  );
  PEWSOS_255 pe_mat_6_5 (
    .io_in_r_data           (pe_mat_6_4_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pe_mat_6_4_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pe_mat_6_4_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pe_mat_6_4_io_out_r_stall        ), //i
    .io_out_r_data          (pe_mat_6_5_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_6_5_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_6_5_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_6_5_io_out_r_stall        ), //o
    .io_in_c_data           (pe_mat_5_5_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pe_mat_5_5_io_out_c_is_stationary), //i
    .io_out_c_data          (pe_mat_6_5_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_6_5_io_out_c_is_stationary), //o
    .clk                    (clk                              ), //i
    .reset                  (reset                            )  //i
  );
  PEWSOS_255 pe_mat_6_6 (
    .io_in_r_data           (pe_mat_6_5_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pe_mat_6_5_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pe_mat_6_5_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pe_mat_6_5_io_out_r_stall        ), //i
    .io_out_r_data          (pe_mat_6_6_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_6_6_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_6_6_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_6_6_io_out_r_stall        ), //o
    .io_in_c_data           (pe_mat_5_6_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pe_mat_5_6_io_out_c_is_stationary), //i
    .io_out_c_data          (pe_mat_6_6_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_6_6_io_out_c_is_stationary), //o
    .clk                    (clk                              ), //i
    .reset                  (reset                            )  //i
  );
  PEWSOS_255 pe_mat_6_7 (
    .io_in_r_data           (pe_mat_6_6_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pe_mat_6_6_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pe_mat_6_6_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pe_mat_6_6_io_out_r_stall        ), //i
    .io_out_r_data          (pe_mat_6_7_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_6_7_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_6_7_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_6_7_io_out_r_stall        ), //o
    .io_in_c_data           (pe_mat_5_7_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pe_mat_5_7_io_out_c_is_stationary), //i
    .io_out_c_data          (pe_mat_6_7_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_6_7_io_out_c_is_stationary), //o
    .clk                    (clk                              ), //i
    .reset                  (reset                            )  //i
  );
  PEWSOS_255 pe_mat_6_8 (
    .io_in_r_data           (pe_mat_6_7_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pe_mat_6_7_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pe_mat_6_7_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pe_mat_6_7_io_out_r_stall        ), //i
    .io_out_r_data          (pe_mat_6_8_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_6_8_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_6_8_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_6_8_io_out_r_stall        ), //o
    .io_in_c_data           (pe_mat_5_8_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pe_mat_5_8_io_out_c_is_stationary), //i
    .io_out_c_data          (pe_mat_6_8_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_6_8_io_out_c_is_stationary), //o
    .clk                    (clk                              ), //i
    .reset                  (reset                            )  //i
  );
  PEWSOS_255 pe_mat_6_9 (
    .io_in_r_data           (pe_mat_6_8_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pe_mat_6_8_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pe_mat_6_8_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pe_mat_6_8_io_out_r_stall        ), //i
    .io_out_r_data          (pe_mat_6_9_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_6_9_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_6_9_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_6_9_io_out_r_stall        ), //o
    .io_in_c_data           (pe_mat_5_9_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pe_mat_5_9_io_out_c_is_stationary), //i
    .io_out_c_data          (pe_mat_6_9_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_6_9_io_out_c_is_stationary), //o
    .clk                    (clk                              ), //i
    .reset                  (reset                            )  //i
  );
  PEWSOS_255 pe_mat_6_10 (
    .io_in_r_data           (pe_mat_6_9_io_out_r_data[15:0]    ), //i
    .io_in_r_load_store     (pe_mat_6_9_io_out_r_load_store    ), //i
    .io_in_r_df_is_ws       (pe_mat_6_9_io_out_r_df_is_ws      ), //i
    .io_in_r_stall          (pe_mat_6_9_io_out_r_stall         ), //i
    .io_out_r_data          (pe_mat_6_10_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_6_10_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_6_10_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_6_10_io_out_r_stall        ), //o
    .io_in_c_data           (pe_mat_5_10_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pe_mat_5_10_io_out_c_is_stationary), //i
    .io_out_c_data          (pe_mat_6_10_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_6_10_io_out_c_is_stationary), //o
    .clk                    (clk                               ), //i
    .reset                  (reset                             )  //i
  );
  PEWSOS_255 pe_mat_6_11 (
    .io_in_r_data           (pe_mat_6_10_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pe_mat_6_10_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pe_mat_6_10_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pe_mat_6_10_io_out_r_stall        ), //i
    .io_out_r_data          (pe_mat_6_11_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_6_11_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_6_11_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_6_11_io_out_r_stall        ), //o
    .io_in_c_data           (pe_mat_5_11_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pe_mat_5_11_io_out_c_is_stationary), //i
    .io_out_c_data          (pe_mat_6_11_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_6_11_io_out_c_is_stationary), //o
    .clk                    (clk                               ), //i
    .reset                  (reset                             )  //i
  );
  PEWSOS_255 pe_mat_6_12 (
    .io_in_r_data           (pe_mat_6_11_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pe_mat_6_11_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pe_mat_6_11_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pe_mat_6_11_io_out_r_stall        ), //i
    .io_out_r_data          (pe_mat_6_12_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_6_12_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_6_12_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_6_12_io_out_r_stall        ), //o
    .io_in_c_data           (pe_mat_5_12_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pe_mat_5_12_io_out_c_is_stationary), //i
    .io_out_c_data          (pe_mat_6_12_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_6_12_io_out_c_is_stationary), //o
    .clk                    (clk                               ), //i
    .reset                  (reset                             )  //i
  );
  PEWSOS_255 pe_mat_6_13 (
    .io_in_r_data           (pe_mat_6_12_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pe_mat_6_12_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pe_mat_6_12_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pe_mat_6_12_io_out_r_stall        ), //i
    .io_out_r_data          (pe_mat_6_13_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_6_13_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_6_13_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_6_13_io_out_r_stall        ), //o
    .io_in_c_data           (pe_mat_5_13_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pe_mat_5_13_io_out_c_is_stationary), //i
    .io_out_c_data          (pe_mat_6_13_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_6_13_io_out_c_is_stationary), //o
    .clk                    (clk                               ), //i
    .reset                  (reset                             )  //i
  );
  PEWSOS_255 pe_mat_6_14 (
    .io_in_r_data           (pe_mat_6_13_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pe_mat_6_13_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pe_mat_6_13_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pe_mat_6_13_io_out_r_stall        ), //i
    .io_out_r_data          (pe_mat_6_14_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_6_14_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_6_14_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_6_14_io_out_r_stall        ), //o
    .io_in_c_data           (pe_mat_5_14_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pe_mat_5_14_io_out_c_is_stationary), //i
    .io_out_c_data          (pe_mat_6_14_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_6_14_io_out_c_is_stationary), //o
    .clk                    (clk                               ), //i
    .reset                  (reset                             )  //i
  );
  PEWSOS_255 pe_mat_6_15 (
    .io_in_r_data           (pe_mat_6_14_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pe_mat_6_14_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pe_mat_6_14_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pe_mat_6_14_io_out_r_stall        ), //i
    .io_out_r_data          (pe_mat_6_15_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_6_15_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_6_15_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_6_15_io_out_r_stall        ), //o
    .io_in_c_data           (pe_mat_5_15_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pe_mat_5_15_io_out_c_is_stationary), //i
    .io_out_c_data          (pe_mat_6_15_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_6_15_io_out_c_is_stationary), //o
    .clk                    (clk                               ), //i
    .reset                  (reset                             )  //i
  );
  PEWSOS_255 pe_mat_7_0 (
    .io_in_r_data           (io_in_r_7_data[15:0]             ), //i
    .io_in_r_load_store     (io_in_r_7_load_store             ), //i
    .io_in_r_df_is_ws       (io_in_r_7_df_is_ws               ), //i
    .io_in_r_stall          (io_in_r_7_stall                  ), //i
    .io_out_r_data          (pe_mat_7_0_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_7_0_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_7_0_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_7_0_io_out_r_stall        ), //o
    .io_in_c_data           (pe_mat_6_0_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pe_mat_6_0_io_out_c_is_stationary), //i
    .io_out_c_data          (pe_mat_7_0_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_7_0_io_out_c_is_stationary), //o
    .clk                    (clk                              ), //i
    .reset                  (reset                            )  //i
  );
  PEWSOS_255 pe_mat_7_1 (
    .io_in_r_data           (pe_mat_7_0_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pe_mat_7_0_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pe_mat_7_0_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pe_mat_7_0_io_out_r_stall        ), //i
    .io_out_r_data          (pe_mat_7_1_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_7_1_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_7_1_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_7_1_io_out_r_stall        ), //o
    .io_in_c_data           (pe_mat_6_1_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pe_mat_6_1_io_out_c_is_stationary), //i
    .io_out_c_data          (pe_mat_7_1_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_7_1_io_out_c_is_stationary), //o
    .clk                    (clk                              ), //i
    .reset                  (reset                            )  //i
  );
  PEWSOS_255 pe_mat_7_2 (
    .io_in_r_data           (pe_mat_7_1_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pe_mat_7_1_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pe_mat_7_1_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pe_mat_7_1_io_out_r_stall        ), //i
    .io_out_r_data          (pe_mat_7_2_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_7_2_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_7_2_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_7_2_io_out_r_stall        ), //o
    .io_in_c_data           (pe_mat_6_2_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pe_mat_6_2_io_out_c_is_stationary), //i
    .io_out_c_data          (pe_mat_7_2_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_7_2_io_out_c_is_stationary), //o
    .clk                    (clk                              ), //i
    .reset                  (reset                            )  //i
  );
  PEWSOS_255 pe_mat_7_3 (
    .io_in_r_data           (pe_mat_7_2_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pe_mat_7_2_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pe_mat_7_2_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pe_mat_7_2_io_out_r_stall        ), //i
    .io_out_r_data          (pe_mat_7_3_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_7_3_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_7_3_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_7_3_io_out_r_stall        ), //o
    .io_in_c_data           (pe_mat_6_3_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pe_mat_6_3_io_out_c_is_stationary), //i
    .io_out_c_data          (pe_mat_7_3_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_7_3_io_out_c_is_stationary), //o
    .clk                    (clk                              ), //i
    .reset                  (reset                            )  //i
  );
  PEWSOS_255 pe_mat_7_4 (
    .io_in_r_data           (pe_mat_7_3_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pe_mat_7_3_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pe_mat_7_3_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pe_mat_7_3_io_out_r_stall        ), //i
    .io_out_r_data          (pe_mat_7_4_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_7_4_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_7_4_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_7_4_io_out_r_stall        ), //o
    .io_in_c_data           (pe_mat_6_4_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pe_mat_6_4_io_out_c_is_stationary), //i
    .io_out_c_data          (pe_mat_7_4_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_7_4_io_out_c_is_stationary), //o
    .clk                    (clk                              ), //i
    .reset                  (reset                            )  //i
  );
  PEWSOS_255 pe_mat_7_5 (
    .io_in_r_data           (pe_mat_7_4_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pe_mat_7_4_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pe_mat_7_4_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pe_mat_7_4_io_out_r_stall        ), //i
    .io_out_r_data          (pe_mat_7_5_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_7_5_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_7_5_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_7_5_io_out_r_stall        ), //o
    .io_in_c_data           (pe_mat_6_5_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pe_mat_6_5_io_out_c_is_stationary), //i
    .io_out_c_data          (pe_mat_7_5_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_7_5_io_out_c_is_stationary), //o
    .clk                    (clk                              ), //i
    .reset                  (reset                            )  //i
  );
  PEWSOS_255 pe_mat_7_6 (
    .io_in_r_data           (pe_mat_7_5_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pe_mat_7_5_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pe_mat_7_5_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pe_mat_7_5_io_out_r_stall        ), //i
    .io_out_r_data          (pe_mat_7_6_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_7_6_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_7_6_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_7_6_io_out_r_stall        ), //o
    .io_in_c_data           (pe_mat_6_6_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pe_mat_6_6_io_out_c_is_stationary), //i
    .io_out_c_data          (pe_mat_7_6_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_7_6_io_out_c_is_stationary), //o
    .clk                    (clk                              ), //i
    .reset                  (reset                            )  //i
  );
  PEWSOS_255 pe_mat_7_7 (
    .io_in_r_data           (pe_mat_7_6_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pe_mat_7_6_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pe_mat_7_6_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pe_mat_7_6_io_out_r_stall        ), //i
    .io_out_r_data          (pe_mat_7_7_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_7_7_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_7_7_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_7_7_io_out_r_stall        ), //o
    .io_in_c_data           (pe_mat_6_7_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pe_mat_6_7_io_out_c_is_stationary), //i
    .io_out_c_data          (pe_mat_7_7_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_7_7_io_out_c_is_stationary), //o
    .clk                    (clk                              ), //i
    .reset                  (reset                            )  //i
  );
  PEWSOS_255 pe_mat_7_8 (
    .io_in_r_data           (pe_mat_7_7_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pe_mat_7_7_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pe_mat_7_7_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pe_mat_7_7_io_out_r_stall        ), //i
    .io_out_r_data          (pe_mat_7_8_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_7_8_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_7_8_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_7_8_io_out_r_stall        ), //o
    .io_in_c_data           (pe_mat_6_8_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pe_mat_6_8_io_out_c_is_stationary), //i
    .io_out_c_data          (pe_mat_7_8_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_7_8_io_out_c_is_stationary), //o
    .clk                    (clk                              ), //i
    .reset                  (reset                            )  //i
  );
  PEWSOS_255 pe_mat_7_9 (
    .io_in_r_data           (pe_mat_7_8_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pe_mat_7_8_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pe_mat_7_8_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pe_mat_7_8_io_out_r_stall        ), //i
    .io_out_r_data          (pe_mat_7_9_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_7_9_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_7_9_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_7_9_io_out_r_stall        ), //o
    .io_in_c_data           (pe_mat_6_9_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pe_mat_6_9_io_out_c_is_stationary), //i
    .io_out_c_data          (pe_mat_7_9_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_7_9_io_out_c_is_stationary), //o
    .clk                    (clk                              ), //i
    .reset                  (reset                            )  //i
  );
  PEWSOS_255 pe_mat_7_10 (
    .io_in_r_data           (pe_mat_7_9_io_out_r_data[15:0]    ), //i
    .io_in_r_load_store     (pe_mat_7_9_io_out_r_load_store    ), //i
    .io_in_r_df_is_ws       (pe_mat_7_9_io_out_r_df_is_ws      ), //i
    .io_in_r_stall          (pe_mat_7_9_io_out_r_stall         ), //i
    .io_out_r_data          (pe_mat_7_10_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_7_10_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_7_10_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_7_10_io_out_r_stall        ), //o
    .io_in_c_data           (pe_mat_6_10_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pe_mat_6_10_io_out_c_is_stationary), //i
    .io_out_c_data          (pe_mat_7_10_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_7_10_io_out_c_is_stationary), //o
    .clk                    (clk                               ), //i
    .reset                  (reset                             )  //i
  );
  PEWSOS_255 pe_mat_7_11 (
    .io_in_r_data           (pe_mat_7_10_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pe_mat_7_10_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pe_mat_7_10_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pe_mat_7_10_io_out_r_stall        ), //i
    .io_out_r_data          (pe_mat_7_11_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_7_11_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_7_11_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_7_11_io_out_r_stall        ), //o
    .io_in_c_data           (pe_mat_6_11_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pe_mat_6_11_io_out_c_is_stationary), //i
    .io_out_c_data          (pe_mat_7_11_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_7_11_io_out_c_is_stationary), //o
    .clk                    (clk                               ), //i
    .reset                  (reset                             )  //i
  );
  PEWSOS_255 pe_mat_7_12 (
    .io_in_r_data           (pe_mat_7_11_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pe_mat_7_11_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pe_mat_7_11_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pe_mat_7_11_io_out_r_stall        ), //i
    .io_out_r_data          (pe_mat_7_12_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_7_12_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_7_12_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_7_12_io_out_r_stall        ), //o
    .io_in_c_data           (pe_mat_6_12_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pe_mat_6_12_io_out_c_is_stationary), //i
    .io_out_c_data          (pe_mat_7_12_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_7_12_io_out_c_is_stationary), //o
    .clk                    (clk                               ), //i
    .reset                  (reset                             )  //i
  );
  PEWSOS_255 pe_mat_7_13 (
    .io_in_r_data           (pe_mat_7_12_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pe_mat_7_12_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pe_mat_7_12_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pe_mat_7_12_io_out_r_stall        ), //i
    .io_out_r_data          (pe_mat_7_13_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_7_13_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_7_13_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_7_13_io_out_r_stall        ), //o
    .io_in_c_data           (pe_mat_6_13_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pe_mat_6_13_io_out_c_is_stationary), //i
    .io_out_c_data          (pe_mat_7_13_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_7_13_io_out_c_is_stationary), //o
    .clk                    (clk                               ), //i
    .reset                  (reset                             )  //i
  );
  PEWSOS_255 pe_mat_7_14 (
    .io_in_r_data           (pe_mat_7_13_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pe_mat_7_13_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pe_mat_7_13_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pe_mat_7_13_io_out_r_stall        ), //i
    .io_out_r_data          (pe_mat_7_14_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_7_14_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_7_14_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_7_14_io_out_r_stall        ), //o
    .io_in_c_data           (pe_mat_6_14_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pe_mat_6_14_io_out_c_is_stationary), //i
    .io_out_c_data          (pe_mat_7_14_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_7_14_io_out_c_is_stationary), //o
    .clk                    (clk                               ), //i
    .reset                  (reset                             )  //i
  );
  PEWSOS_255 pe_mat_7_15 (
    .io_in_r_data           (pe_mat_7_14_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pe_mat_7_14_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pe_mat_7_14_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pe_mat_7_14_io_out_r_stall        ), //i
    .io_out_r_data          (pe_mat_7_15_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_7_15_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_7_15_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_7_15_io_out_r_stall        ), //o
    .io_in_c_data           (pe_mat_6_15_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pe_mat_6_15_io_out_c_is_stationary), //i
    .io_out_c_data          (pe_mat_7_15_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_7_15_io_out_c_is_stationary), //o
    .clk                    (clk                               ), //i
    .reset                  (reset                             )  //i
  );
  PEWSOS_255 pe_mat_8_0 (
    .io_in_r_data           (io_in_r_8_data[15:0]             ), //i
    .io_in_r_load_store     (io_in_r_8_load_store             ), //i
    .io_in_r_df_is_ws       (io_in_r_8_df_is_ws               ), //i
    .io_in_r_stall          (io_in_r_8_stall                  ), //i
    .io_out_r_data          (pe_mat_8_0_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_8_0_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_8_0_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_8_0_io_out_r_stall        ), //o
    .io_in_c_data           (pe_mat_7_0_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pe_mat_7_0_io_out_c_is_stationary), //i
    .io_out_c_data          (pe_mat_8_0_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_8_0_io_out_c_is_stationary), //o
    .clk                    (clk                              ), //i
    .reset                  (reset                            )  //i
  );
  PEWSOS_255 pe_mat_8_1 (
    .io_in_r_data           (pe_mat_8_0_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pe_mat_8_0_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pe_mat_8_0_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pe_mat_8_0_io_out_r_stall        ), //i
    .io_out_r_data          (pe_mat_8_1_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_8_1_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_8_1_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_8_1_io_out_r_stall        ), //o
    .io_in_c_data           (pe_mat_7_1_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pe_mat_7_1_io_out_c_is_stationary), //i
    .io_out_c_data          (pe_mat_8_1_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_8_1_io_out_c_is_stationary), //o
    .clk                    (clk                              ), //i
    .reset                  (reset                            )  //i
  );
  PEWSOS_255 pe_mat_8_2 (
    .io_in_r_data           (pe_mat_8_1_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pe_mat_8_1_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pe_mat_8_1_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pe_mat_8_1_io_out_r_stall        ), //i
    .io_out_r_data          (pe_mat_8_2_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_8_2_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_8_2_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_8_2_io_out_r_stall        ), //o
    .io_in_c_data           (pe_mat_7_2_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pe_mat_7_2_io_out_c_is_stationary), //i
    .io_out_c_data          (pe_mat_8_2_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_8_2_io_out_c_is_stationary), //o
    .clk                    (clk                              ), //i
    .reset                  (reset                            )  //i
  );
  PEWSOS_255 pe_mat_8_3 (
    .io_in_r_data           (pe_mat_8_2_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pe_mat_8_2_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pe_mat_8_2_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pe_mat_8_2_io_out_r_stall        ), //i
    .io_out_r_data          (pe_mat_8_3_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_8_3_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_8_3_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_8_3_io_out_r_stall        ), //o
    .io_in_c_data           (pe_mat_7_3_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pe_mat_7_3_io_out_c_is_stationary), //i
    .io_out_c_data          (pe_mat_8_3_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_8_3_io_out_c_is_stationary), //o
    .clk                    (clk                              ), //i
    .reset                  (reset                            )  //i
  );
  PEWSOS_255 pe_mat_8_4 (
    .io_in_r_data           (pe_mat_8_3_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pe_mat_8_3_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pe_mat_8_3_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pe_mat_8_3_io_out_r_stall        ), //i
    .io_out_r_data          (pe_mat_8_4_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_8_4_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_8_4_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_8_4_io_out_r_stall        ), //o
    .io_in_c_data           (pe_mat_7_4_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pe_mat_7_4_io_out_c_is_stationary), //i
    .io_out_c_data          (pe_mat_8_4_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_8_4_io_out_c_is_stationary), //o
    .clk                    (clk                              ), //i
    .reset                  (reset                            )  //i
  );
  PEWSOS_255 pe_mat_8_5 (
    .io_in_r_data           (pe_mat_8_4_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pe_mat_8_4_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pe_mat_8_4_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pe_mat_8_4_io_out_r_stall        ), //i
    .io_out_r_data          (pe_mat_8_5_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_8_5_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_8_5_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_8_5_io_out_r_stall        ), //o
    .io_in_c_data           (pe_mat_7_5_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pe_mat_7_5_io_out_c_is_stationary), //i
    .io_out_c_data          (pe_mat_8_5_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_8_5_io_out_c_is_stationary), //o
    .clk                    (clk                              ), //i
    .reset                  (reset                            )  //i
  );
  PEWSOS_255 pe_mat_8_6 (
    .io_in_r_data           (pe_mat_8_5_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pe_mat_8_5_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pe_mat_8_5_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pe_mat_8_5_io_out_r_stall        ), //i
    .io_out_r_data          (pe_mat_8_6_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_8_6_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_8_6_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_8_6_io_out_r_stall        ), //o
    .io_in_c_data           (pe_mat_7_6_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pe_mat_7_6_io_out_c_is_stationary), //i
    .io_out_c_data          (pe_mat_8_6_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_8_6_io_out_c_is_stationary), //o
    .clk                    (clk                              ), //i
    .reset                  (reset                            )  //i
  );
  PEWSOS_255 pe_mat_8_7 (
    .io_in_r_data           (pe_mat_8_6_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pe_mat_8_6_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pe_mat_8_6_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pe_mat_8_6_io_out_r_stall        ), //i
    .io_out_r_data          (pe_mat_8_7_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_8_7_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_8_7_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_8_7_io_out_r_stall        ), //o
    .io_in_c_data           (pe_mat_7_7_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pe_mat_7_7_io_out_c_is_stationary), //i
    .io_out_c_data          (pe_mat_8_7_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_8_7_io_out_c_is_stationary), //o
    .clk                    (clk                              ), //i
    .reset                  (reset                            )  //i
  );
  PEWSOS_255 pe_mat_8_8 (
    .io_in_r_data           (pe_mat_8_7_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pe_mat_8_7_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pe_mat_8_7_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pe_mat_8_7_io_out_r_stall        ), //i
    .io_out_r_data          (pe_mat_8_8_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_8_8_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_8_8_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_8_8_io_out_r_stall        ), //o
    .io_in_c_data           (pe_mat_7_8_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pe_mat_7_8_io_out_c_is_stationary), //i
    .io_out_c_data          (pe_mat_8_8_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_8_8_io_out_c_is_stationary), //o
    .clk                    (clk                              ), //i
    .reset                  (reset                            )  //i
  );
  PEWSOS_255 pe_mat_8_9 (
    .io_in_r_data           (pe_mat_8_8_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pe_mat_8_8_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pe_mat_8_8_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pe_mat_8_8_io_out_r_stall        ), //i
    .io_out_r_data          (pe_mat_8_9_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_8_9_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_8_9_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_8_9_io_out_r_stall        ), //o
    .io_in_c_data           (pe_mat_7_9_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pe_mat_7_9_io_out_c_is_stationary), //i
    .io_out_c_data          (pe_mat_8_9_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_8_9_io_out_c_is_stationary), //o
    .clk                    (clk                              ), //i
    .reset                  (reset                            )  //i
  );
  PEWSOS_255 pe_mat_8_10 (
    .io_in_r_data           (pe_mat_8_9_io_out_r_data[15:0]    ), //i
    .io_in_r_load_store     (pe_mat_8_9_io_out_r_load_store    ), //i
    .io_in_r_df_is_ws       (pe_mat_8_9_io_out_r_df_is_ws      ), //i
    .io_in_r_stall          (pe_mat_8_9_io_out_r_stall         ), //i
    .io_out_r_data          (pe_mat_8_10_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_8_10_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_8_10_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_8_10_io_out_r_stall        ), //o
    .io_in_c_data           (pe_mat_7_10_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pe_mat_7_10_io_out_c_is_stationary), //i
    .io_out_c_data          (pe_mat_8_10_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_8_10_io_out_c_is_stationary), //o
    .clk                    (clk                               ), //i
    .reset                  (reset                             )  //i
  );
  PEWSOS_255 pe_mat_8_11 (
    .io_in_r_data           (pe_mat_8_10_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pe_mat_8_10_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pe_mat_8_10_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pe_mat_8_10_io_out_r_stall        ), //i
    .io_out_r_data          (pe_mat_8_11_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_8_11_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_8_11_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_8_11_io_out_r_stall        ), //o
    .io_in_c_data           (pe_mat_7_11_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pe_mat_7_11_io_out_c_is_stationary), //i
    .io_out_c_data          (pe_mat_8_11_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_8_11_io_out_c_is_stationary), //o
    .clk                    (clk                               ), //i
    .reset                  (reset                             )  //i
  );
  PEWSOS_255 pe_mat_8_12 (
    .io_in_r_data           (pe_mat_8_11_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pe_mat_8_11_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pe_mat_8_11_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pe_mat_8_11_io_out_r_stall        ), //i
    .io_out_r_data          (pe_mat_8_12_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_8_12_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_8_12_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_8_12_io_out_r_stall        ), //o
    .io_in_c_data           (pe_mat_7_12_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pe_mat_7_12_io_out_c_is_stationary), //i
    .io_out_c_data          (pe_mat_8_12_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_8_12_io_out_c_is_stationary), //o
    .clk                    (clk                               ), //i
    .reset                  (reset                             )  //i
  );
  PEWSOS_255 pe_mat_8_13 (
    .io_in_r_data           (pe_mat_8_12_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pe_mat_8_12_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pe_mat_8_12_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pe_mat_8_12_io_out_r_stall        ), //i
    .io_out_r_data          (pe_mat_8_13_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_8_13_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_8_13_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_8_13_io_out_r_stall        ), //o
    .io_in_c_data           (pe_mat_7_13_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pe_mat_7_13_io_out_c_is_stationary), //i
    .io_out_c_data          (pe_mat_8_13_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_8_13_io_out_c_is_stationary), //o
    .clk                    (clk                               ), //i
    .reset                  (reset                             )  //i
  );
  PEWSOS_255 pe_mat_8_14 (
    .io_in_r_data           (pe_mat_8_13_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pe_mat_8_13_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pe_mat_8_13_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pe_mat_8_13_io_out_r_stall        ), //i
    .io_out_r_data          (pe_mat_8_14_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_8_14_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_8_14_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_8_14_io_out_r_stall        ), //o
    .io_in_c_data           (pe_mat_7_14_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pe_mat_7_14_io_out_c_is_stationary), //i
    .io_out_c_data          (pe_mat_8_14_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_8_14_io_out_c_is_stationary), //o
    .clk                    (clk                               ), //i
    .reset                  (reset                             )  //i
  );
  PEWSOS_255 pe_mat_8_15 (
    .io_in_r_data           (pe_mat_8_14_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pe_mat_8_14_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pe_mat_8_14_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pe_mat_8_14_io_out_r_stall        ), //i
    .io_out_r_data          (pe_mat_8_15_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_8_15_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_8_15_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_8_15_io_out_r_stall        ), //o
    .io_in_c_data           (pe_mat_7_15_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pe_mat_7_15_io_out_c_is_stationary), //i
    .io_out_c_data          (pe_mat_8_15_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_8_15_io_out_c_is_stationary), //o
    .clk                    (clk                               ), //i
    .reset                  (reset                             )  //i
  );
  PEWSOS_255 pe_mat_9_0 (
    .io_in_r_data           (io_in_r_9_data[15:0]             ), //i
    .io_in_r_load_store     (io_in_r_9_load_store             ), //i
    .io_in_r_df_is_ws       (io_in_r_9_df_is_ws               ), //i
    .io_in_r_stall          (io_in_r_9_stall                  ), //i
    .io_out_r_data          (pe_mat_9_0_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_9_0_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_9_0_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_9_0_io_out_r_stall        ), //o
    .io_in_c_data           (pe_mat_8_0_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pe_mat_8_0_io_out_c_is_stationary), //i
    .io_out_c_data          (pe_mat_9_0_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_9_0_io_out_c_is_stationary), //o
    .clk                    (clk                              ), //i
    .reset                  (reset                            )  //i
  );
  PEWSOS_255 pe_mat_9_1 (
    .io_in_r_data           (pe_mat_9_0_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pe_mat_9_0_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pe_mat_9_0_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pe_mat_9_0_io_out_r_stall        ), //i
    .io_out_r_data          (pe_mat_9_1_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_9_1_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_9_1_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_9_1_io_out_r_stall        ), //o
    .io_in_c_data           (pe_mat_8_1_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pe_mat_8_1_io_out_c_is_stationary), //i
    .io_out_c_data          (pe_mat_9_1_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_9_1_io_out_c_is_stationary), //o
    .clk                    (clk                              ), //i
    .reset                  (reset                            )  //i
  );
  PEWSOS_255 pe_mat_9_2 (
    .io_in_r_data           (pe_mat_9_1_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pe_mat_9_1_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pe_mat_9_1_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pe_mat_9_1_io_out_r_stall        ), //i
    .io_out_r_data          (pe_mat_9_2_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_9_2_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_9_2_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_9_2_io_out_r_stall        ), //o
    .io_in_c_data           (pe_mat_8_2_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pe_mat_8_2_io_out_c_is_stationary), //i
    .io_out_c_data          (pe_mat_9_2_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_9_2_io_out_c_is_stationary), //o
    .clk                    (clk                              ), //i
    .reset                  (reset                            )  //i
  );
  PEWSOS_255 pe_mat_9_3 (
    .io_in_r_data           (pe_mat_9_2_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pe_mat_9_2_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pe_mat_9_2_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pe_mat_9_2_io_out_r_stall        ), //i
    .io_out_r_data          (pe_mat_9_3_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_9_3_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_9_3_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_9_3_io_out_r_stall        ), //o
    .io_in_c_data           (pe_mat_8_3_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pe_mat_8_3_io_out_c_is_stationary), //i
    .io_out_c_data          (pe_mat_9_3_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_9_3_io_out_c_is_stationary), //o
    .clk                    (clk                              ), //i
    .reset                  (reset                            )  //i
  );
  PEWSOS_255 pe_mat_9_4 (
    .io_in_r_data           (pe_mat_9_3_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pe_mat_9_3_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pe_mat_9_3_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pe_mat_9_3_io_out_r_stall        ), //i
    .io_out_r_data          (pe_mat_9_4_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_9_4_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_9_4_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_9_4_io_out_r_stall        ), //o
    .io_in_c_data           (pe_mat_8_4_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pe_mat_8_4_io_out_c_is_stationary), //i
    .io_out_c_data          (pe_mat_9_4_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_9_4_io_out_c_is_stationary), //o
    .clk                    (clk                              ), //i
    .reset                  (reset                            )  //i
  );
  PEWSOS_255 pe_mat_9_5 (
    .io_in_r_data           (pe_mat_9_4_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pe_mat_9_4_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pe_mat_9_4_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pe_mat_9_4_io_out_r_stall        ), //i
    .io_out_r_data          (pe_mat_9_5_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_9_5_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_9_5_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_9_5_io_out_r_stall        ), //o
    .io_in_c_data           (pe_mat_8_5_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pe_mat_8_5_io_out_c_is_stationary), //i
    .io_out_c_data          (pe_mat_9_5_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_9_5_io_out_c_is_stationary), //o
    .clk                    (clk                              ), //i
    .reset                  (reset                            )  //i
  );
  PEWSOS_255 pe_mat_9_6 (
    .io_in_r_data           (pe_mat_9_5_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pe_mat_9_5_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pe_mat_9_5_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pe_mat_9_5_io_out_r_stall        ), //i
    .io_out_r_data          (pe_mat_9_6_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_9_6_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_9_6_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_9_6_io_out_r_stall        ), //o
    .io_in_c_data           (pe_mat_8_6_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pe_mat_8_6_io_out_c_is_stationary), //i
    .io_out_c_data          (pe_mat_9_6_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_9_6_io_out_c_is_stationary), //o
    .clk                    (clk                              ), //i
    .reset                  (reset                            )  //i
  );
  PEWSOS_255 pe_mat_9_7 (
    .io_in_r_data           (pe_mat_9_6_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pe_mat_9_6_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pe_mat_9_6_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pe_mat_9_6_io_out_r_stall        ), //i
    .io_out_r_data          (pe_mat_9_7_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_9_7_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_9_7_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_9_7_io_out_r_stall        ), //o
    .io_in_c_data           (pe_mat_8_7_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pe_mat_8_7_io_out_c_is_stationary), //i
    .io_out_c_data          (pe_mat_9_7_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_9_7_io_out_c_is_stationary), //o
    .clk                    (clk                              ), //i
    .reset                  (reset                            )  //i
  );
  PEWSOS_255 pe_mat_9_8 (
    .io_in_r_data           (pe_mat_9_7_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pe_mat_9_7_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pe_mat_9_7_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pe_mat_9_7_io_out_r_stall        ), //i
    .io_out_r_data          (pe_mat_9_8_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_9_8_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_9_8_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_9_8_io_out_r_stall        ), //o
    .io_in_c_data           (pe_mat_8_8_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pe_mat_8_8_io_out_c_is_stationary), //i
    .io_out_c_data          (pe_mat_9_8_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_9_8_io_out_c_is_stationary), //o
    .clk                    (clk                              ), //i
    .reset                  (reset                            )  //i
  );
  PEWSOS_255 pe_mat_9_9 (
    .io_in_r_data           (pe_mat_9_8_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pe_mat_9_8_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pe_mat_9_8_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pe_mat_9_8_io_out_r_stall        ), //i
    .io_out_r_data          (pe_mat_9_9_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_9_9_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_9_9_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_9_9_io_out_r_stall        ), //o
    .io_in_c_data           (pe_mat_8_9_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pe_mat_8_9_io_out_c_is_stationary), //i
    .io_out_c_data          (pe_mat_9_9_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_9_9_io_out_c_is_stationary), //o
    .clk                    (clk                              ), //i
    .reset                  (reset                            )  //i
  );
  PEWSOS_255 pe_mat_9_10 (
    .io_in_r_data           (pe_mat_9_9_io_out_r_data[15:0]    ), //i
    .io_in_r_load_store     (pe_mat_9_9_io_out_r_load_store    ), //i
    .io_in_r_df_is_ws       (pe_mat_9_9_io_out_r_df_is_ws      ), //i
    .io_in_r_stall          (pe_mat_9_9_io_out_r_stall         ), //i
    .io_out_r_data          (pe_mat_9_10_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_9_10_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_9_10_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_9_10_io_out_r_stall        ), //o
    .io_in_c_data           (pe_mat_8_10_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pe_mat_8_10_io_out_c_is_stationary), //i
    .io_out_c_data          (pe_mat_9_10_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_9_10_io_out_c_is_stationary), //o
    .clk                    (clk                               ), //i
    .reset                  (reset                             )  //i
  );
  PEWSOS_255 pe_mat_9_11 (
    .io_in_r_data           (pe_mat_9_10_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pe_mat_9_10_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pe_mat_9_10_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pe_mat_9_10_io_out_r_stall        ), //i
    .io_out_r_data          (pe_mat_9_11_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_9_11_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_9_11_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_9_11_io_out_r_stall        ), //o
    .io_in_c_data           (pe_mat_8_11_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pe_mat_8_11_io_out_c_is_stationary), //i
    .io_out_c_data          (pe_mat_9_11_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_9_11_io_out_c_is_stationary), //o
    .clk                    (clk                               ), //i
    .reset                  (reset                             )  //i
  );
  PEWSOS_255 pe_mat_9_12 (
    .io_in_r_data           (pe_mat_9_11_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pe_mat_9_11_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pe_mat_9_11_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pe_mat_9_11_io_out_r_stall        ), //i
    .io_out_r_data          (pe_mat_9_12_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_9_12_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_9_12_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_9_12_io_out_r_stall        ), //o
    .io_in_c_data           (pe_mat_8_12_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pe_mat_8_12_io_out_c_is_stationary), //i
    .io_out_c_data          (pe_mat_9_12_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_9_12_io_out_c_is_stationary), //o
    .clk                    (clk                               ), //i
    .reset                  (reset                             )  //i
  );
  PEWSOS_255 pe_mat_9_13 (
    .io_in_r_data           (pe_mat_9_12_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pe_mat_9_12_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pe_mat_9_12_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pe_mat_9_12_io_out_r_stall        ), //i
    .io_out_r_data          (pe_mat_9_13_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_9_13_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_9_13_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_9_13_io_out_r_stall        ), //o
    .io_in_c_data           (pe_mat_8_13_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pe_mat_8_13_io_out_c_is_stationary), //i
    .io_out_c_data          (pe_mat_9_13_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_9_13_io_out_c_is_stationary), //o
    .clk                    (clk                               ), //i
    .reset                  (reset                             )  //i
  );
  PEWSOS_255 pe_mat_9_14 (
    .io_in_r_data           (pe_mat_9_13_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pe_mat_9_13_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pe_mat_9_13_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pe_mat_9_13_io_out_r_stall        ), //i
    .io_out_r_data          (pe_mat_9_14_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_9_14_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_9_14_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_9_14_io_out_r_stall        ), //o
    .io_in_c_data           (pe_mat_8_14_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pe_mat_8_14_io_out_c_is_stationary), //i
    .io_out_c_data          (pe_mat_9_14_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_9_14_io_out_c_is_stationary), //o
    .clk                    (clk                               ), //i
    .reset                  (reset                             )  //i
  );
  PEWSOS_255 pe_mat_9_15 (
    .io_in_r_data           (pe_mat_9_14_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pe_mat_9_14_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pe_mat_9_14_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pe_mat_9_14_io_out_r_stall        ), //i
    .io_out_r_data          (pe_mat_9_15_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_9_15_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_9_15_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_9_15_io_out_r_stall        ), //o
    .io_in_c_data           (pe_mat_8_15_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pe_mat_8_15_io_out_c_is_stationary), //i
    .io_out_c_data          (pe_mat_9_15_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_9_15_io_out_c_is_stationary), //o
    .clk                    (clk                               ), //i
    .reset                  (reset                             )  //i
  );
  PEWSOS_255 pe_mat_10_0 (
    .io_in_r_data           (io_in_r_10_data[15:0]             ), //i
    .io_in_r_load_store     (io_in_r_10_load_store             ), //i
    .io_in_r_df_is_ws       (io_in_r_10_df_is_ws               ), //i
    .io_in_r_stall          (io_in_r_10_stall                  ), //i
    .io_out_r_data          (pe_mat_10_0_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_10_0_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_10_0_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_10_0_io_out_r_stall        ), //o
    .io_in_c_data           (pe_mat_9_0_io_out_c_data[15:0]    ), //i
    .io_in_c_is_stationary  (pe_mat_9_0_io_out_c_is_stationary ), //i
    .io_out_c_data          (pe_mat_10_0_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_10_0_io_out_c_is_stationary), //o
    .clk                    (clk                               ), //i
    .reset                  (reset                             )  //i
  );
  PEWSOS_255 pe_mat_10_1 (
    .io_in_r_data           (pe_mat_10_0_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pe_mat_10_0_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pe_mat_10_0_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pe_mat_10_0_io_out_r_stall        ), //i
    .io_out_r_data          (pe_mat_10_1_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_10_1_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_10_1_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_10_1_io_out_r_stall        ), //o
    .io_in_c_data           (pe_mat_9_1_io_out_c_data[15:0]    ), //i
    .io_in_c_is_stationary  (pe_mat_9_1_io_out_c_is_stationary ), //i
    .io_out_c_data          (pe_mat_10_1_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_10_1_io_out_c_is_stationary), //o
    .clk                    (clk                               ), //i
    .reset                  (reset                             )  //i
  );
  PEWSOS_255 pe_mat_10_2 (
    .io_in_r_data           (pe_mat_10_1_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pe_mat_10_1_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pe_mat_10_1_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pe_mat_10_1_io_out_r_stall        ), //i
    .io_out_r_data          (pe_mat_10_2_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_10_2_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_10_2_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_10_2_io_out_r_stall        ), //o
    .io_in_c_data           (pe_mat_9_2_io_out_c_data[15:0]    ), //i
    .io_in_c_is_stationary  (pe_mat_9_2_io_out_c_is_stationary ), //i
    .io_out_c_data          (pe_mat_10_2_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_10_2_io_out_c_is_stationary), //o
    .clk                    (clk                               ), //i
    .reset                  (reset                             )  //i
  );
  PEWSOS_255 pe_mat_10_3 (
    .io_in_r_data           (pe_mat_10_2_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pe_mat_10_2_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pe_mat_10_2_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pe_mat_10_2_io_out_r_stall        ), //i
    .io_out_r_data          (pe_mat_10_3_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_10_3_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_10_3_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_10_3_io_out_r_stall        ), //o
    .io_in_c_data           (pe_mat_9_3_io_out_c_data[15:0]    ), //i
    .io_in_c_is_stationary  (pe_mat_9_3_io_out_c_is_stationary ), //i
    .io_out_c_data          (pe_mat_10_3_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_10_3_io_out_c_is_stationary), //o
    .clk                    (clk                               ), //i
    .reset                  (reset                             )  //i
  );
  PEWSOS_255 pe_mat_10_4 (
    .io_in_r_data           (pe_mat_10_3_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pe_mat_10_3_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pe_mat_10_3_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pe_mat_10_3_io_out_r_stall        ), //i
    .io_out_r_data          (pe_mat_10_4_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_10_4_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_10_4_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_10_4_io_out_r_stall        ), //o
    .io_in_c_data           (pe_mat_9_4_io_out_c_data[15:0]    ), //i
    .io_in_c_is_stationary  (pe_mat_9_4_io_out_c_is_stationary ), //i
    .io_out_c_data          (pe_mat_10_4_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_10_4_io_out_c_is_stationary), //o
    .clk                    (clk                               ), //i
    .reset                  (reset                             )  //i
  );
  PEWSOS_255 pe_mat_10_5 (
    .io_in_r_data           (pe_mat_10_4_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pe_mat_10_4_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pe_mat_10_4_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pe_mat_10_4_io_out_r_stall        ), //i
    .io_out_r_data          (pe_mat_10_5_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_10_5_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_10_5_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_10_5_io_out_r_stall        ), //o
    .io_in_c_data           (pe_mat_9_5_io_out_c_data[15:0]    ), //i
    .io_in_c_is_stationary  (pe_mat_9_5_io_out_c_is_stationary ), //i
    .io_out_c_data          (pe_mat_10_5_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_10_5_io_out_c_is_stationary), //o
    .clk                    (clk                               ), //i
    .reset                  (reset                             )  //i
  );
  PEWSOS_255 pe_mat_10_6 (
    .io_in_r_data           (pe_mat_10_5_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pe_mat_10_5_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pe_mat_10_5_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pe_mat_10_5_io_out_r_stall        ), //i
    .io_out_r_data          (pe_mat_10_6_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_10_6_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_10_6_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_10_6_io_out_r_stall        ), //o
    .io_in_c_data           (pe_mat_9_6_io_out_c_data[15:0]    ), //i
    .io_in_c_is_stationary  (pe_mat_9_6_io_out_c_is_stationary ), //i
    .io_out_c_data          (pe_mat_10_6_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_10_6_io_out_c_is_stationary), //o
    .clk                    (clk                               ), //i
    .reset                  (reset                             )  //i
  );
  PEWSOS_255 pe_mat_10_7 (
    .io_in_r_data           (pe_mat_10_6_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pe_mat_10_6_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pe_mat_10_6_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pe_mat_10_6_io_out_r_stall        ), //i
    .io_out_r_data          (pe_mat_10_7_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_10_7_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_10_7_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_10_7_io_out_r_stall        ), //o
    .io_in_c_data           (pe_mat_9_7_io_out_c_data[15:0]    ), //i
    .io_in_c_is_stationary  (pe_mat_9_7_io_out_c_is_stationary ), //i
    .io_out_c_data          (pe_mat_10_7_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_10_7_io_out_c_is_stationary), //o
    .clk                    (clk                               ), //i
    .reset                  (reset                             )  //i
  );
  PEWSOS_255 pe_mat_10_8 (
    .io_in_r_data           (pe_mat_10_7_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pe_mat_10_7_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pe_mat_10_7_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pe_mat_10_7_io_out_r_stall        ), //i
    .io_out_r_data          (pe_mat_10_8_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_10_8_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_10_8_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_10_8_io_out_r_stall        ), //o
    .io_in_c_data           (pe_mat_9_8_io_out_c_data[15:0]    ), //i
    .io_in_c_is_stationary  (pe_mat_9_8_io_out_c_is_stationary ), //i
    .io_out_c_data          (pe_mat_10_8_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_10_8_io_out_c_is_stationary), //o
    .clk                    (clk                               ), //i
    .reset                  (reset                             )  //i
  );
  PEWSOS_255 pe_mat_10_9 (
    .io_in_r_data           (pe_mat_10_8_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pe_mat_10_8_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pe_mat_10_8_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pe_mat_10_8_io_out_r_stall        ), //i
    .io_out_r_data          (pe_mat_10_9_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_10_9_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_10_9_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_10_9_io_out_r_stall        ), //o
    .io_in_c_data           (pe_mat_9_9_io_out_c_data[15:0]    ), //i
    .io_in_c_is_stationary  (pe_mat_9_9_io_out_c_is_stationary ), //i
    .io_out_c_data          (pe_mat_10_9_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_10_9_io_out_c_is_stationary), //o
    .clk                    (clk                               ), //i
    .reset                  (reset                             )  //i
  );
  PEWSOS_255 pe_mat_10_10 (
    .io_in_r_data           (pe_mat_10_9_io_out_r_data[15:0]    ), //i
    .io_in_r_load_store     (pe_mat_10_9_io_out_r_load_store    ), //i
    .io_in_r_df_is_ws       (pe_mat_10_9_io_out_r_df_is_ws      ), //i
    .io_in_r_stall          (pe_mat_10_9_io_out_r_stall         ), //i
    .io_out_r_data          (pe_mat_10_10_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_10_10_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_10_10_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_10_10_io_out_r_stall        ), //o
    .io_in_c_data           (pe_mat_9_10_io_out_c_data[15:0]    ), //i
    .io_in_c_is_stationary  (pe_mat_9_10_io_out_c_is_stationary ), //i
    .io_out_c_data          (pe_mat_10_10_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_10_10_io_out_c_is_stationary), //o
    .clk                    (clk                                ), //i
    .reset                  (reset                              )  //i
  );
  PEWSOS_255 pe_mat_10_11 (
    .io_in_r_data           (pe_mat_10_10_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pe_mat_10_10_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pe_mat_10_10_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pe_mat_10_10_io_out_r_stall        ), //i
    .io_out_r_data          (pe_mat_10_11_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_10_11_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_10_11_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_10_11_io_out_r_stall        ), //o
    .io_in_c_data           (pe_mat_9_11_io_out_c_data[15:0]    ), //i
    .io_in_c_is_stationary  (pe_mat_9_11_io_out_c_is_stationary ), //i
    .io_out_c_data          (pe_mat_10_11_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_10_11_io_out_c_is_stationary), //o
    .clk                    (clk                                ), //i
    .reset                  (reset                              )  //i
  );
  PEWSOS_255 pe_mat_10_12 (
    .io_in_r_data           (pe_mat_10_11_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pe_mat_10_11_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pe_mat_10_11_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pe_mat_10_11_io_out_r_stall        ), //i
    .io_out_r_data          (pe_mat_10_12_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_10_12_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_10_12_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_10_12_io_out_r_stall        ), //o
    .io_in_c_data           (pe_mat_9_12_io_out_c_data[15:0]    ), //i
    .io_in_c_is_stationary  (pe_mat_9_12_io_out_c_is_stationary ), //i
    .io_out_c_data          (pe_mat_10_12_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_10_12_io_out_c_is_stationary), //o
    .clk                    (clk                                ), //i
    .reset                  (reset                              )  //i
  );
  PEWSOS_255 pe_mat_10_13 (
    .io_in_r_data           (pe_mat_10_12_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pe_mat_10_12_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pe_mat_10_12_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pe_mat_10_12_io_out_r_stall        ), //i
    .io_out_r_data          (pe_mat_10_13_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_10_13_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_10_13_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_10_13_io_out_r_stall        ), //o
    .io_in_c_data           (pe_mat_9_13_io_out_c_data[15:0]    ), //i
    .io_in_c_is_stationary  (pe_mat_9_13_io_out_c_is_stationary ), //i
    .io_out_c_data          (pe_mat_10_13_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_10_13_io_out_c_is_stationary), //o
    .clk                    (clk                                ), //i
    .reset                  (reset                              )  //i
  );
  PEWSOS_255 pe_mat_10_14 (
    .io_in_r_data           (pe_mat_10_13_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pe_mat_10_13_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pe_mat_10_13_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pe_mat_10_13_io_out_r_stall        ), //i
    .io_out_r_data          (pe_mat_10_14_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_10_14_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_10_14_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_10_14_io_out_r_stall        ), //o
    .io_in_c_data           (pe_mat_9_14_io_out_c_data[15:0]    ), //i
    .io_in_c_is_stationary  (pe_mat_9_14_io_out_c_is_stationary ), //i
    .io_out_c_data          (pe_mat_10_14_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_10_14_io_out_c_is_stationary), //o
    .clk                    (clk                                ), //i
    .reset                  (reset                              )  //i
  );
  PEWSOS_255 pe_mat_10_15 (
    .io_in_r_data           (pe_mat_10_14_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pe_mat_10_14_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pe_mat_10_14_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pe_mat_10_14_io_out_r_stall        ), //i
    .io_out_r_data          (pe_mat_10_15_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_10_15_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_10_15_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_10_15_io_out_r_stall        ), //o
    .io_in_c_data           (pe_mat_9_15_io_out_c_data[15:0]    ), //i
    .io_in_c_is_stationary  (pe_mat_9_15_io_out_c_is_stationary ), //i
    .io_out_c_data          (pe_mat_10_15_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_10_15_io_out_c_is_stationary), //o
    .clk                    (clk                                ), //i
    .reset                  (reset                              )  //i
  );
  PEWSOS_255 pe_mat_11_0 (
    .io_in_r_data           (io_in_r_11_data[15:0]             ), //i
    .io_in_r_load_store     (io_in_r_11_load_store             ), //i
    .io_in_r_df_is_ws       (io_in_r_11_df_is_ws               ), //i
    .io_in_r_stall          (io_in_r_11_stall                  ), //i
    .io_out_r_data          (pe_mat_11_0_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_11_0_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_11_0_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_11_0_io_out_r_stall        ), //o
    .io_in_c_data           (pe_mat_10_0_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pe_mat_10_0_io_out_c_is_stationary), //i
    .io_out_c_data          (pe_mat_11_0_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_11_0_io_out_c_is_stationary), //o
    .clk                    (clk                               ), //i
    .reset                  (reset                             )  //i
  );
  PEWSOS_255 pe_mat_11_1 (
    .io_in_r_data           (pe_mat_11_0_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pe_mat_11_0_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pe_mat_11_0_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pe_mat_11_0_io_out_r_stall        ), //i
    .io_out_r_data          (pe_mat_11_1_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_11_1_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_11_1_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_11_1_io_out_r_stall        ), //o
    .io_in_c_data           (pe_mat_10_1_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pe_mat_10_1_io_out_c_is_stationary), //i
    .io_out_c_data          (pe_mat_11_1_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_11_1_io_out_c_is_stationary), //o
    .clk                    (clk                               ), //i
    .reset                  (reset                             )  //i
  );
  PEWSOS_255 pe_mat_11_2 (
    .io_in_r_data           (pe_mat_11_1_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pe_mat_11_1_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pe_mat_11_1_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pe_mat_11_1_io_out_r_stall        ), //i
    .io_out_r_data          (pe_mat_11_2_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_11_2_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_11_2_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_11_2_io_out_r_stall        ), //o
    .io_in_c_data           (pe_mat_10_2_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pe_mat_10_2_io_out_c_is_stationary), //i
    .io_out_c_data          (pe_mat_11_2_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_11_2_io_out_c_is_stationary), //o
    .clk                    (clk                               ), //i
    .reset                  (reset                             )  //i
  );
  PEWSOS_255 pe_mat_11_3 (
    .io_in_r_data           (pe_mat_11_2_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pe_mat_11_2_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pe_mat_11_2_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pe_mat_11_2_io_out_r_stall        ), //i
    .io_out_r_data          (pe_mat_11_3_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_11_3_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_11_3_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_11_3_io_out_r_stall        ), //o
    .io_in_c_data           (pe_mat_10_3_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pe_mat_10_3_io_out_c_is_stationary), //i
    .io_out_c_data          (pe_mat_11_3_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_11_3_io_out_c_is_stationary), //o
    .clk                    (clk                               ), //i
    .reset                  (reset                             )  //i
  );
  PEWSOS_255 pe_mat_11_4 (
    .io_in_r_data           (pe_mat_11_3_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pe_mat_11_3_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pe_mat_11_3_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pe_mat_11_3_io_out_r_stall        ), //i
    .io_out_r_data          (pe_mat_11_4_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_11_4_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_11_4_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_11_4_io_out_r_stall        ), //o
    .io_in_c_data           (pe_mat_10_4_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pe_mat_10_4_io_out_c_is_stationary), //i
    .io_out_c_data          (pe_mat_11_4_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_11_4_io_out_c_is_stationary), //o
    .clk                    (clk                               ), //i
    .reset                  (reset                             )  //i
  );
  PEWSOS_255 pe_mat_11_5 (
    .io_in_r_data           (pe_mat_11_4_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pe_mat_11_4_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pe_mat_11_4_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pe_mat_11_4_io_out_r_stall        ), //i
    .io_out_r_data          (pe_mat_11_5_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_11_5_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_11_5_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_11_5_io_out_r_stall        ), //o
    .io_in_c_data           (pe_mat_10_5_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pe_mat_10_5_io_out_c_is_stationary), //i
    .io_out_c_data          (pe_mat_11_5_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_11_5_io_out_c_is_stationary), //o
    .clk                    (clk                               ), //i
    .reset                  (reset                             )  //i
  );
  PEWSOS_255 pe_mat_11_6 (
    .io_in_r_data           (pe_mat_11_5_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pe_mat_11_5_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pe_mat_11_5_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pe_mat_11_5_io_out_r_stall        ), //i
    .io_out_r_data          (pe_mat_11_6_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_11_6_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_11_6_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_11_6_io_out_r_stall        ), //o
    .io_in_c_data           (pe_mat_10_6_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pe_mat_10_6_io_out_c_is_stationary), //i
    .io_out_c_data          (pe_mat_11_6_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_11_6_io_out_c_is_stationary), //o
    .clk                    (clk                               ), //i
    .reset                  (reset                             )  //i
  );
  PEWSOS_255 pe_mat_11_7 (
    .io_in_r_data           (pe_mat_11_6_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pe_mat_11_6_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pe_mat_11_6_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pe_mat_11_6_io_out_r_stall        ), //i
    .io_out_r_data          (pe_mat_11_7_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_11_7_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_11_7_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_11_7_io_out_r_stall        ), //o
    .io_in_c_data           (pe_mat_10_7_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pe_mat_10_7_io_out_c_is_stationary), //i
    .io_out_c_data          (pe_mat_11_7_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_11_7_io_out_c_is_stationary), //o
    .clk                    (clk                               ), //i
    .reset                  (reset                             )  //i
  );
  PEWSOS_255 pe_mat_11_8 (
    .io_in_r_data           (pe_mat_11_7_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pe_mat_11_7_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pe_mat_11_7_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pe_mat_11_7_io_out_r_stall        ), //i
    .io_out_r_data          (pe_mat_11_8_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_11_8_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_11_8_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_11_8_io_out_r_stall        ), //o
    .io_in_c_data           (pe_mat_10_8_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pe_mat_10_8_io_out_c_is_stationary), //i
    .io_out_c_data          (pe_mat_11_8_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_11_8_io_out_c_is_stationary), //o
    .clk                    (clk                               ), //i
    .reset                  (reset                             )  //i
  );
  PEWSOS_255 pe_mat_11_9 (
    .io_in_r_data           (pe_mat_11_8_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pe_mat_11_8_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pe_mat_11_8_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pe_mat_11_8_io_out_r_stall        ), //i
    .io_out_r_data          (pe_mat_11_9_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_11_9_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_11_9_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_11_9_io_out_r_stall        ), //o
    .io_in_c_data           (pe_mat_10_9_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pe_mat_10_9_io_out_c_is_stationary), //i
    .io_out_c_data          (pe_mat_11_9_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_11_9_io_out_c_is_stationary), //o
    .clk                    (clk                               ), //i
    .reset                  (reset                             )  //i
  );
  PEWSOS_255 pe_mat_11_10 (
    .io_in_r_data           (pe_mat_11_9_io_out_r_data[15:0]    ), //i
    .io_in_r_load_store     (pe_mat_11_9_io_out_r_load_store    ), //i
    .io_in_r_df_is_ws       (pe_mat_11_9_io_out_r_df_is_ws      ), //i
    .io_in_r_stall          (pe_mat_11_9_io_out_r_stall         ), //i
    .io_out_r_data          (pe_mat_11_10_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_11_10_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_11_10_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_11_10_io_out_r_stall        ), //o
    .io_in_c_data           (pe_mat_10_10_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pe_mat_10_10_io_out_c_is_stationary), //i
    .io_out_c_data          (pe_mat_11_10_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_11_10_io_out_c_is_stationary), //o
    .clk                    (clk                                ), //i
    .reset                  (reset                              )  //i
  );
  PEWSOS_255 pe_mat_11_11 (
    .io_in_r_data           (pe_mat_11_10_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pe_mat_11_10_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pe_mat_11_10_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pe_mat_11_10_io_out_r_stall        ), //i
    .io_out_r_data          (pe_mat_11_11_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_11_11_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_11_11_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_11_11_io_out_r_stall        ), //o
    .io_in_c_data           (pe_mat_10_11_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pe_mat_10_11_io_out_c_is_stationary), //i
    .io_out_c_data          (pe_mat_11_11_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_11_11_io_out_c_is_stationary), //o
    .clk                    (clk                                ), //i
    .reset                  (reset                              )  //i
  );
  PEWSOS_255 pe_mat_11_12 (
    .io_in_r_data           (pe_mat_11_11_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pe_mat_11_11_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pe_mat_11_11_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pe_mat_11_11_io_out_r_stall        ), //i
    .io_out_r_data          (pe_mat_11_12_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_11_12_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_11_12_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_11_12_io_out_r_stall        ), //o
    .io_in_c_data           (pe_mat_10_12_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pe_mat_10_12_io_out_c_is_stationary), //i
    .io_out_c_data          (pe_mat_11_12_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_11_12_io_out_c_is_stationary), //o
    .clk                    (clk                                ), //i
    .reset                  (reset                              )  //i
  );
  PEWSOS_255 pe_mat_11_13 (
    .io_in_r_data           (pe_mat_11_12_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pe_mat_11_12_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pe_mat_11_12_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pe_mat_11_12_io_out_r_stall        ), //i
    .io_out_r_data          (pe_mat_11_13_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_11_13_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_11_13_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_11_13_io_out_r_stall        ), //o
    .io_in_c_data           (pe_mat_10_13_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pe_mat_10_13_io_out_c_is_stationary), //i
    .io_out_c_data          (pe_mat_11_13_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_11_13_io_out_c_is_stationary), //o
    .clk                    (clk                                ), //i
    .reset                  (reset                              )  //i
  );
  PEWSOS_255 pe_mat_11_14 (
    .io_in_r_data           (pe_mat_11_13_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pe_mat_11_13_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pe_mat_11_13_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pe_mat_11_13_io_out_r_stall        ), //i
    .io_out_r_data          (pe_mat_11_14_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_11_14_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_11_14_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_11_14_io_out_r_stall        ), //o
    .io_in_c_data           (pe_mat_10_14_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pe_mat_10_14_io_out_c_is_stationary), //i
    .io_out_c_data          (pe_mat_11_14_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_11_14_io_out_c_is_stationary), //o
    .clk                    (clk                                ), //i
    .reset                  (reset                              )  //i
  );
  PEWSOS_255 pe_mat_11_15 (
    .io_in_r_data           (pe_mat_11_14_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pe_mat_11_14_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pe_mat_11_14_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pe_mat_11_14_io_out_r_stall        ), //i
    .io_out_r_data          (pe_mat_11_15_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_11_15_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_11_15_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_11_15_io_out_r_stall        ), //o
    .io_in_c_data           (pe_mat_10_15_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pe_mat_10_15_io_out_c_is_stationary), //i
    .io_out_c_data          (pe_mat_11_15_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_11_15_io_out_c_is_stationary), //o
    .clk                    (clk                                ), //i
    .reset                  (reset                              )  //i
  );
  PEWSOS_255 pe_mat_12_0 (
    .io_in_r_data           (io_in_r_12_data[15:0]             ), //i
    .io_in_r_load_store     (io_in_r_12_load_store             ), //i
    .io_in_r_df_is_ws       (io_in_r_12_df_is_ws               ), //i
    .io_in_r_stall          (io_in_r_12_stall                  ), //i
    .io_out_r_data          (pe_mat_12_0_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_12_0_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_12_0_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_12_0_io_out_r_stall        ), //o
    .io_in_c_data           (pe_mat_11_0_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pe_mat_11_0_io_out_c_is_stationary), //i
    .io_out_c_data          (pe_mat_12_0_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_12_0_io_out_c_is_stationary), //o
    .clk                    (clk                               ), //i
    .reset                  (reset                             )  //i
  );
  PEWSOS_255 pe_mat_12_1 (
    .io_in_r_data           (pe_mat_12_0_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pe_mat_12_0_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pe_mat_12_0_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pe_mat_12_0_io_out_r_stall        ), //i
    .io_out_r_data          (pe_mat_12_1_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_12_1_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_12_1_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_12_1_io_out_r_stall        ), //o
    .io_in_c_data           (pe_mat_11_1_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pe_mat_11_1_io_out_c_is_stationary), //i
    .io_out_c_data          (pe_mat_12_1_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_12_1_io_out_c_is_stationary), //o
    .clk                    (clk                               ), //i
    .reset                  (reset                             )  //i
  );
  PEWSOS_255 pe_mat_12_2 (
    .io_in_r_data           (pe_mat_12_1_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pe_mat_12_1_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pe_mat_12_1_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pe_mat_12_1_io_out_r_stall        ), //i
    .io_out_r_data          (pe_mat_12_2_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_12_2_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_12_2_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_12_2_io_out_r_stall        ), //o
    .io_in_c_data           (pe_mat_11_2_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pe_mat_11_2_io_out_c_is_stationary), //i
    .io_out_c_data          (pe_mat_12_2_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_12_2_io_out_c_is_stationary), //o
    .clk                    (clk                               ), //i
    .reset                  (reset                             )  //i
  );
  PEWSOS_255 pe_mat_12_3 (
    .io_in_r_data           (pe_mat_12_2_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pe_mat_12_2_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pe_mat_12_2_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pe_mat_12_2_io_out_r_stall        ), //i
    .io_out_r_data          (pe_mat_12_3_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_12_3_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_12_3_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_12_3_io_out_r_stall        ), //o
    .io_in_c_data           (pe_mat_11_3_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pe_mat_11_3_io_out_c_is_stationary), //i
    .io_out_c_data          (pe_mat_12_3_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_12_3_io_out_c_is_stationary), //o
    .clk                    (clk                               ), //i
    .reset                  (reset                             )  //i
  );
  PEWSOS_255 pe_mat_12_4 (
    .io_in_r_data           (pe_mat_12_3_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pe_mat_12_3_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pe_mat_12_3_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pe_mat_12_3_io_out_r_stall        ), //i
    .io_out_r_data          (pe_mat_12_4_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_12_4_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_12_4_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_12_4_io_out_r_stall        ), //o
    .io_in_c_data           (pe_mat_11_4_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pe_mat_11_4_io_out_c_is_stationary), //i
    .io_out_c_data          (pe_mat_12_4_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_12_4_io_out_c_is_stationary), //o
    .clk                    (clk                               ), //i
    .reset                  (reset                             )  //i
  );
  PEWSOS_255 pe_mat_12_5 (
    .io_in_r_data           (pe_mat_12_4_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pe_mat_12_4_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pe_mat_12_4_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pe_mat_12_4_io_out_r_stall        ), //i
    .io_out_r_data          (pe_mat_12_5_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_12_5_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_12_5_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_12_5_io_out_r_stall        ), //o
    .io_in_c_data           (pe_mat_11_5_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pe_mat_11_5_io_out_c_is_stationary), //i
    .io_out_c_data          (pe_mat_12_5_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_12_5_io_out_c_is_stationary), //o
    .clk                    (clk                               ), //i
    .reset                  (reset                             )  //i
  );
  PEWSOS_255 pe_mat_12_6 (
    .io_in_r_data           (pe_mat_12_5_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pe_mat_12_5_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pe_mat_12_5_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pe_mat_12_5_io_out_r_stall        ), //i
    .io_out_r_data          (pe_mat_12_6_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_12_6_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_12_6_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_12_6_io_out_r_stall        ), //o
    .io_in_c_data           (pe_mat_11_6_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pe_mat_11_6_io_out_c_is_stationary), //i
    .io_out_c_data          (pe_mat_12_6_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_12_6_io_out_c_is_stationary), //o
    .clk                    (clk                               ), //i
    .reset                  (reset                             )  //i
  );
  PEWSOS_255 pe_mat_12_7 (
    .io_in_r_data           (pe_mat_12_6_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pe_mat_12_6_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pe_mat_12_6_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pe_mat_12_6_io_out_r_stall        ), //i
    .io_out_r_data          (pe_mat_12_7_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_12_7_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_12_7_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_12_7_io_out_r_stall        ), //o
    .io_in_c_data           (pe_mat_11_7_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pe_mat_11_7_io_out_c_is_stationary), //i
    .io_out_c_data          (pe_mat_12_7_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_12_7_io_out_c_is_stationary), //o
    .clk                    (clk                               ), //i
    .reset                  (reset                             )  //i
  );
  PEWSOS_255 pe_mat_12_8 (
    .io_in_r_data           (pe_mat_12_7_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pe_mat_12_7_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pe_mat_12_7_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pe_mat_12_7_io_out_r_stall        ), //i
    .io_out_r_data          (pe_mat_12_8_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_12_8_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_12_8_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_12_8_io_out_r_stall        ), //o
    .io_in_c_data           (pe_mat_11_8_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pe_mat_11_8_io_out_c_is_stationary), //i
    .io_out_c_data          (pe_mat_12_8_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_12_8_io_out_c_is_stationary), //o
    .clk                    (clk                               ), //i
    .reset                  (reset                             )  //i
  );
  PEWSOS_255 pe_mat_12_9 (
    .io_in_r_data           (pe_mat_12_8_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pe_mat_12_8_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pe_mat_12_8_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pe_mat_12_8_io_out_r_stall        ), //i
    .io_out_r_data          (pe_mat_12_9_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_12_9_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_12_9_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_12_9_io_out_r_stall        ), //o
    .io_in_c_data           (pe_mat_11_9_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pe_mat_11_9_io_out_c_is_stationary), //i
    .io_out_c_data          (pe_mat_12_9_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_12_9_io_out_c_is_stationary), //o
    .clk                    (clk                               ), //i
    .reset                  (reset                             )  //i
  );
  PEWSOS_255 pe_mat_12_10 (
    .io_in_r_data           (pe_mat_12_9_io_out_r_data[15:0]    ), //i
    .io_in_r_load_store     (pe_mat_12_9_io_out_r_load_store    ), //i
    .io_in_r_df_is_ws       (pe_mat_12_9_io_out_r_df_is_ws      ), //i
    .io_in_r_stall          (pe_mat_12_9_io_out_r_stall         ), //i
    .io_out_r_data          (pe_mat_12_10_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_12_10_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_12_10_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_12_10_io_out_r_stall        ), //o
    .io_in_c_data           (pe_mat_11_10_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pe_mat_11_10_io_out_c_is_stationary), //i
    .io_out_c_data          (pe_mat_12_10_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_12_10_io_out_c_is_stationary), //o
    .clk                    (clk                                ), //i
    .reset                  (reset                              )  //i
  );
  PEWSOS_255 pe_mat_12_11 (
    .io_in_r_data           (pe_mat_12_10_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pe_mat_12_10_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pe_mat_12_10_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pe_mat_12_10_io_out_r_stall        ), //i
    .io_out_r_data          (pe_mat_12_11_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_12_11_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_12_11_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_12_11_io_out_r_stall        ), //o
    .io_in_c_data           (pe_mat_11_11_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pe_mat_11_11_io_out_c_is_stationary), //i
    .io_out_c_data          (pe_mat_12_11_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_12_11_io_out_c_is_stationary), //o
    .clk                    (clk                                ), //i
    .reset                  (reset                              )  //i
  );
  PEWSOS_255 pe_mat_12_12 (
    .io_in_r_data           (pe_mat_12_11_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pe_mat_12_11_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pe_mat_12_11_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pe_mat_12_11_io_out_r_stall        ), //i
    .io_out_r_data          (pe_mat_12_12_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_12_12_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_12_12_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_12_12_io_out_r_stall        ), //o
    .io_in_c_data           (pe_mat_11_12_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pe_mat_11_12_io_out_c_is_stationary), //i
    .io_out_c_data          (pe_mat_12_12_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_12_12_io_out_c_is_stationary), //o
    .clk                    (clk                                ), //i
    .reset                  (reset                              )  //i
  );
  PEWSOS_255 pe_mat_12_13 (
    .io_in_r_data           (pe_mat_12_12_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pe_mat_12_12_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pe_mat_12_12_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pe_mat_12_12_io_out_r_stall        ), //i
    .io_out_r_data          (pe_mat_12_13_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_12_13_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_12_13_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_12_13_io_out_r_stall        ), //o
    .io_in_c_data           (pe_mat_11_13_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pe_mat_11_13_io_out_c_is_stationary), //i
    .io_out_c_data          (pe_mat_12_13_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_12_13_io_out_c_is_stationary), //o
    .clk                    (clk                                ), //i
    .reset                  (reset                              )  //i
  );
  PEWSOS_255 pe_mat_12_14 (
    .io_in_r_data           (pe_mat_12_13_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pe_mat_12_13_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pe_mat_12_13_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pe_mat_12_13_io_out_r_stall        ), //i
    .io_out_r_data          (pe_mat_12_14_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_12_14_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_12_14_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_12_14_io_out_r_stall        ), //o
    .io_in_c_data           (pe_mat_11_14_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pe_mat_11_14_io_out_c_is_stationary), //i
    .io_out_c_data          (pe_mat_12_14_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_12_14_io_out_c_is_stationary), //o
    .clk                    (clk                                ), //i
    .reset                  (reset                              )  //i
  );
  PEWSOS_255 pe_mat_12_15 (
    .io_in_r_data           (pe_mat_12_14_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pe_mat_12_14_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pe_mat_12_14_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pe_mat_12_14_io_out_r_stall        ), //i
    .io_out_r_data          (pe_mat_12_15_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_12_15_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_12_15_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_12_15_io_out_r_stall        ), //o
    .io_in_c_data           (pe_mat_11_15_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pe_mat_11_15_io_out_c_is_stationary), //i
    .io_out_c_data          (pe_mat_12_15_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_12_15_io_out_c_is_stationary), //o
    .clk                    (clk                                ), //i
    .reset                  (reset                              )  //i
  );
  PEWSOS_255 pe_mat_13_0 (
    .io_in_r_data           (io_in_r_13_data[15:0]             ), //i
    .io_in_r_load_store     (io_in_r_13_load_store             ), //i
    .io_in_r_df_is_ws       (io_in_r_13_df_is_ws               ), //i
    .io_in_r_stall          (io_in_r_13_stall                  ), //i
    .io_out_r_data          (pe_mat_13_0_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_13_0_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_13_0_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_13_0_io_out_r_stall        ), //o
    .io_in_c_data           (pe_mat_12_0_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pe_mat_12_0_io_out_c_is_stationary), //i
    .io_out_c_data          (pe_mat_13_0_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_13_0_io_out_c_is_stationary), //o
    .clk                    (clk                               ), //i
    .reset                  (reset                             )  //i
  );
  PEWSOS_255 pe_mat_13_1 (
    .io_in_r_data           (pe_mat_13_0_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pe_mat_13_0_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pe_mat_13_0_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pe_mat_13_0_io_out_r_stall        ), //i
    .io_out_r_data          (pe_mat_13_1_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_13_1_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_13_1_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_13_1_io_out_r_stall        ), //o
    .io_in_c_data           (pe_mat_12_1_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pe_mat_12_1_io_out_c_is_stationary), //i
    .io_out_c_data          (pe_mat_13_1_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_13_1_io_out_c_is_stationary), //o
    .clk                    (clk                               ), //i
    .reset                  (reset                             )  //i
  );
  PEWSOS_255 pe_mat_13_2 (
    .io_in_r_data           (pe_mat_13_1_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pe_mat_13_1_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pe_mat_13_1_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pe_mat_13_1_io_out_r_stall        ), //i
    .io_out_r_data          (pe_mat_13_2_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_13_2_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_13_2_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_13_2_io_out_r_stall        ), //o
    .io_in_c_data           (pe_mat_12_2_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pe_mat_12_2_io_out_c_is_stationary), //i
    .io_out_c_data          (pe_mat_13_2_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_13_2_io_out_c_is_stationary), //o
    .clk                    (clk                               ), //i
    .reset                  (reset                             )  //i
  );
  PEWSOS_255 pe_mat_13_3 (
    .io_in_r_data           (pe_mat_13_2_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pe_mat_13_2_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pe_mat_13_2_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pe_mat_13_2_io_out_r_stall        ), //i
    .io_out_r_data          (pe_mat_13_3_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_13_3_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_13_3_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_13_3_io_out_r_stall        ), //o
    .io_in_c_data           (pe_mat_12_3_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pe_mat_12_3_io_out_c_is_stationary), //i
    .io_out_c_data          (pe_mat_13_3_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_13_3_io_out_c_is_stationary), //o
    .clk                    (clk                               ), //i
    .reset                  (reset                             )  //i
  );
  PEWSOS_255 pe_mat_13_4 (
    .io_in_r_data           (pe_mat_13_3_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pe_mat_13_3_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pe_mat_13_3_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pe_mat_13_3_io_out_r_stall        ), //i
    .io_out_r_data          (pe_mat_13_4_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_13_4_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_13_4_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_13_4_io_out_r_stall        ), //o
    .io_in_c_data           (pe_mat_12_4_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pe_mat_12_4_io_out_c_is_stationary), //i
    .io_out_c_data          (pe_mat_13_4_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_13_4_io_out_c_is_stationary), //o
    .clk                    (clk                               ), //i
    .reset                  (reset                             )  //i
  );
  PEWSOS_255 pe_mat_13_5 (
    .io_in_r_data           (pe_mat_13_4_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pe_mat_13_4_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pe_mat_13_4_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pe_mat_13_4_io_out_r_stall        ), //i
    .io_out_r_data          (pe_mat_13_5_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_13_5_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_13_5_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_13_5_io_out_r_stall        ), //o
    .io_in_c_data           (pe_mat_12_5_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pe_mat_12_5_io_out_c_is_stationary), //i
    .io_out_c_data          (pe_mat_13_5_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_13_5_io_out_c_is_stationary), //o
    .clk                    (clk                               ), //i
    .reset                  (reset                             )  //i
  );
  PEWSOS_255 pe_mat_13_6 (
    .io_in_r_data           (pe_mat_13_5_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pe_mat_13_5_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pe_mat_13_5_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pe_mat_13_5_io_out_r_stall        ), //i
    .io_out_r_data          (pe_mat_13_6_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_13_6_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_13_6_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_13_6_io_out_r_stall        ), //o
    .io_in_c_data           (pe_mat_12_6_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pe_mat_12_6_io_out_c_is_stationary), //i
    .io_out_c_data          (pe_mat_13_6_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_13_6_io_out_c_is_stationary), //o
    .clk                    (clk                               ), //i
    .reset                  (reset                             )  //i
  );
  PEWSOS_255 pe_mat_13_7 (
    .io_in_r_data           (pe_mat_13_6_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pe_mat_13_6_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pe_mat_13_6_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pe_mat_13_6_io_out_r_stall        ), //i
    .io_out_r_data          (pe_mat_13_7_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_13_7_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_13_7_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_13_7_io_out_r_stall        ), //o
    .io_in_c_data           (pe_mat_12_7_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pe_mat_12_7_io_out_c_is_stationary), //i
    .io_out_c_data          (pe_mat_13_7_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_13_7_io_out_c_is_stationary), //o
    .clk                    (clk                               ), //i
    .reset                  (reset                             )  //i
  );
  PEWSOS_255 pe_mat_13_8 (
    .io_in_r_data           (pe_mat_13_7_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pe_mat_13_7_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pe_mat_13_7_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pe_mat_13_7_io_out_r_stall        ), //i
    .io_out_r_data          (pe_mat_13_8_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_13_8_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_13_8_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_13_8_io_out_r_stall        ), //o
    .io_in_c_data           (pe_mat_12_8_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pe_mat_12_8_io_out_c_is_stationary), //i
    .io_out_c_data          (pe_mat_13_8_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_13_8_io_out_c_is_stationary), //o
    .clk                    (clk                               ), //i
    .reset                  (reset                             )  //i
  );
  PEWSOS_255 pe_mat_13_9 (
    .io_in_r_data           (pe_mat_13_8_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pe_mat_13_8_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pe_mat_13_8_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pe_mat_13_8_io_out_r_stall        ), //i
    .io_out_r_data          (pe_mat_13_9_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_13_9_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_13_9_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_13_9_io_out_r_stall        ), //o
    .io_in_c_data           (pe_mat_12_9_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pe_mat_12_9_io_out_c_is_stationary), //i
    .io_out_c_data          (pe_mat_13_9_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_13_9_io_out_c_is_stationary), //o
    .clk                    (clk                               ), //i
    .reset                  (reset                             )  //i
  );
  PEWSOS_255 pe_mat_13_10 (
    .io_in_r_data           (pe_mat_13_9_io_out_r_data[15:0]    ), //i
    .io_in_r_load_store     (pe_mat_13_9_io_out_r_load_store    ), //i
    .io_in_r_df_is_ws       (pe_mat_13_9_io_out_r_df_is_ws      ), //i
    .io_in_r_stall          (pe_mat_13_9_io_out_r_stall         ), //i
    .io_out_r_data          (pe_mat_13_10_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_13_10_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_13_10_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_13_10_io_out_r_stall        ), //o
    .io_in_c_data           (pe_mat_12_10_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pe_mat_12_10_io_out_c_is_stationary), //i
    .io_out_c_data          (pe_mat_13_10_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_13_10_io_out_c_is_stationary), //o
    .clk                    (clk                                ), //i
    .reset                  (reset                              )  //i
  );
  PEWSOS_255 pe_mat_13_11 (
    .io_in_r_data           (pe_mat_13_10_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pe_mat_13_10_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pe_mat_13_10_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pe_mat_13_10_io_out_r_stall        ), //i
    .io_out_r_data          (pe_mat_13_11_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_13_11_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_13_11_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_13_11_io_out_r_stall        ), //o
    .io_in_c_data           (pe_mat_12_11_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pe_mat_12_11_io_out_c_is_stationary), //i
    .io_out_c_data          (pe_mat_13_11_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_13_11_io_out_c_is_stationary), //o
    .clk                    (clk                                ), //i
    .reset                  (reset                              )  //i
  );
  PEWSOS_255 pe_mat_13_12 (
    .io_in_r_data           (pe_mat_13_11_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pe_mat_13_11_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pe_mat_13_11_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pe_mat_13_11_io_out_r_stall        ), //i
    .io_out_r_data          (pe_mat_13_12_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_13_12_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_13_12_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_13_12_io_out_r_stall        ), //o
    .io_in_c_data           (pe_mat_12_12_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pe_mat_12_12_io_out_c_is_stationary), //i
    .io_out_c_data          (pe_mat_13_12_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_13_12_io_out_c_is_stationary), //o
    .clk                    (clk                                ), //i
    .reset                  (reset                              )  //i
  );
  PEWSOS_255 pe_mat_13_13 (
    .io_in_r_data           (pe_mat_13_12_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pe_mat_13_12_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pe_mat_13_12_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pe_mat_13_12_io_out_r_stall        ), //i
    .io_out_r_data          (pe_mat_13_13_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_13_13_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_13_13_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_13_13_io_out_r_stall        ), //o
    .io_in_c_data           (pe_mat_12_13_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pe_mat_12_13_io_out_c_is_stationary), //i
    .io_out_c_data          (pe_mat_13_13_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_13_13_io_out_c_is_stationary), //o
    .clk                    (clk                                ), //i
    .reset                  (reset                              )  //i
  );
  PEWSOS_255 pe_mat_13_14 (
    .io_in_r_data           (pe_mat_13_13_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pe_mat_13_13_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pe_mat_13_13_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pe_mat_13_13_io_out_r_stall        ), //i
    .io_out_r_data          (pe_mat_13_14_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_13_14_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_13_14_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_13_14_io_out_r_stall        ), //o
    .io_in_c_data           (pe_mat_12_14_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pe_mat_12_14_io_out_c_is_stationary), //i
    .io_out_c_data          (pe_mat_13_14_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_13_14_io_out_c_is_stationary), //o
    .clk                    (clk                                ), //i
    .reset                  (reset                              )  //i
  );
  PEWSOS_255 pe_mat_13_15 (
    .io_in_r_data           (pe_mat_13_14_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pe_mat_13_14_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pe_mat_13_14_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pe_mat_13_14_io_out_r_stall        ), //i
    .io_out_r_data          (pe_mat_13_15_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_13_15_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_13_15_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_13_15_io_out_r_stall        ), //o
    .io_in_c_data           (pe_mat_12_15_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pe_mat_12_15_io_out_c_is_stationary), //i
    .io_out_c_data          (pe_mat_13_15_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_13_15_io_out_c_is_stationary), //o
    .clk                    (clk                                ), //i
    .reset                  (reset                              )  //i
  );
  PEWSOS_255 pe_mat_14_0 (
    .io_in_r_data           (io_in_r_14_data[15:0]             ), //i
    .io_in_r_load_store     (io_in_r_14_load_store             ), //i
    .io_in_r_df_is_ws       (io_in_r_14_df_is_ws               ), //i
    .io_in_r_stall          (io_in_r_14_stall                  ), //i
    .io_out_r_data          (pe_mat_14_0_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_14_0_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_14_0_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_14_0_io_out_r_stall        ), //o
    .io_in_c_data           (pe_mat_13_0_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pe_mat_13_0_io_out_c_is_stationary), //i
    .io_out_c_data          (pe_mat_14_0_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_14_0_io_out_c_is_stationary), //o
    .clk                    (clk                               ), //i
    .reset                  (reset                             )  //i
  );
  PEWSOS_255 pe_mat_14_1 (
    .io_in_r_data           (pe_mat_14_0_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pe_mat_14_0_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pe_mat_14_0_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pe_mat_14_0_io_out_r_stall        ), //i
    .io_out_r_data          (pe_mat_14_1_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_14_1_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_14_1_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_14_1_io_out_r_stall        ), //o
    .io_in_c_data           (pe_mat_13_1_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pe_mat_13_1_io_out_c_is_stationary), //i
    .io_out_c_data          (pe_mat_14_1_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_14_1_io_out_c_is_stationary), //o
    .clk                    (clk                               ), //i
    .reset                  (reset                             )  //i
  );
  PEWSOS_255 pe_mat_14_2 (
    .io_in_r_data           (pe_mat_14_1_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pe_mat_14_1_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pe_mat_14_1_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pe_mat_14_1_io_out_r_stall        ), //i
    .io_out_r_data          (pe_mat_14_2_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_14_2_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_14_2_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_14_2_io_out_r_stall        ), //o
    .io_in_c_data           (pe_mat_13_2_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pe_mat_13_2_io_out_c_is_stationary), //i
    .io_out_c_data          (pe_mat_14_2_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_14_2_io_out_c_is_stationary), //o
    .clk                    (clk                               ), //i
    .reset                  (reset                             )  //i
  );
  PEWSOS_255 pe_mat_14_3 (
    .io_in_r_data           (pe_mat_14_2_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pe_mat_14_2_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pe_mat_14_2_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pe_mat_14_2_io_out_r_stall        ), //i
    .io_out_r_data          (pe_mat_14_3_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_14_3_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_14_3_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_14_3_io_out_r_stall        ), //o
    .io_in_c_data           (pe_mat_13_3_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pe_mat_13_3_io_out_c_is_stationary), //i
    .io_out_c_data          (pe_mat_14_3_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_14_3_io_out_c_is_stationary), //o
    .clk                    (clk                               ), //i
    .reset                  (reset                             )  //i
  );
  PEWSOS_255 pe_mat_14_4 (
    .io_in_r_data           (pe_mat_14_3_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pe_mat_14_3_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pe_mat_14_3_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pe_mat_14_3_io_out_r_stall        ), //i
    .io_out_r_data          (pe_mat_14_4_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_14_4_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_14_4_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_14_4_io_out_r_stall        ), //o
    .io_in_c_data           (pe_mat_13_4_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pe_mat_13_4_io_out_c_is_stationary), //i
    .io_out_c_data          (pe_mat_14_4_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_14_4_io_out_c_is_stationary), //o
    .clk                    (clk                               ), //i
    .reset                  (reset                             )  //i
  );
  PEWSOS_255 pe_mat_14_5 (
    .io_in_r_data           (pe_mat_14_4_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pe_mat_14_4_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pe_mat_14_4_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pe_mat_14_4_io_out_r_stall        ), //i
    .io_out_r_data          (pe_mat_14_5_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_14_5_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_14_5_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_14_5_io_out_r_stall        ), //o
    .io_in_c_data           (pe_mat_13_5_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pe_mat_13_5_io_out_c_is_stationary), //i
    .io_out_c_data          (pe_mat_14_5_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_14_5_io_out_c_is_stationary), //o
    .clk                    (clk                               ), //i
    .reset                  (reset                             )  //i
  );
  PEWSOS_255 pe_mat_14_6 (
    .io_in_r_data           (pe_mat_14_5_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pe_mat_14_5_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pe_mat_14_5_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pe_mat_14_5_io_out_r_stall        ), //i
    .io_out_r_data          (pe_mat_14_6_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_14_6_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_14_6_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_14_6_io_out_r_stall        ), //o
    .io_in_c_data           (pe_mat_13_6_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pe_mat_13_6_io_out_c_is_stationary), //i
    .io_out_c_data          (pe_mat_14_6_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_14_6_io_out_c_is_stationary), //o
    .clk                    (clk                               ), //i
    .reset                  (reset                             )  //i
  );
  PEWSOS_255 pe_mat_14_7 (
    .io_in_r_data           (pe_mat_14_6_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pe_mat_14_6_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pe_mat_14_6_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pe_mat_14_6_io_out_r_stall        ), //i
    .io_out_r_data          (pe_mat_14_7_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_14_7_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_14_7_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_14_7_io_out_r_stall        ), //o
    .io_in_c_data           (pe_mat_13_7_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pe_mat_13_7_io_out_c_is_stationary), //i
    .io_out_c_data          (pe_mat_14_7_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_14_7_io_out_c_is_stationary), //o
    .clk                    (clk                               ), //i
    .reset                  (reset                             )  //i
  );
  PEWSOS_255 pe_mat_14_8 (
    .io_in_r_data           (pe_mat_14_7_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pe_mat_14_7_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pe_mat_14_7_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pe_mat_14_7_io_out_r_stall        ), //i
    .io_out_r_data          (pe_mat_14_8_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_14_8_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_14_8_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_14_8_io_out_r_stall        ), //o
    .io_in_c_data           (pe_mat_13_8_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pe_mat_13_8_io_out_c_is_stationary), //i
    .io_out_c_data          (pe_mat_14_8_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_14_8_io_out_c_is_stationary), //o
    .clk                    (clk                               ), //i
    .reset                  (reset                             )  //i
  );
  PEWSOS_255 pe_mat_14_9 (
    .io_in_r_data           (pe_mat_14_8_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pe_mat_14_8_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pe_mat_14_8_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pe_mat_14_8_io_out_r_stall        ), //i
    .io_out_r_data          (pe_mat_14_9_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_14_9_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_14_9_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_14_9_io_out_r_stall        ), //o
    .io_in_c_data           (pe_mat_13_9_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pe_mat_13_9_io_out_c_is_stationary), //i
    .io_out_c_data          (pe_mat_14_9_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_14_9_io_out_c_is_stationary), //o
    .clk                    (clk                               ), //i
    .reset                  (reset                             )  //i
  );
  PEWSOS_255 pe_mat_14_10 (
    .io_in_r_data           (pe_mat_14_9_io_out_r_data[15:0]    ), //i
    .io_in_r_load_store     (pe_mat_14_9_io_out_r_load_store    ), //i
    .io_in_r_df_is_ws       (pe_mat_14_9_io_out_r_df_is_ws      ), //i
    .io_in_r_stall          (pe_mat_14_9_io_out_r_stall         ), //i
    .io_out_r_data          (pe_mat_14_10_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_14_10_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_14_10_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_14_10_io_out_r_stall        ), //o
    .io_in_c_data           (pe_mat_13_10_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pe_mat_13_10_io_out_c_is_stationary), //i
    .io_out_c_data          (pe_mat_14_10_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_14_10_io_out_c_is_stationary), //o
    .clk                    (clk                                ), //i
    .reset                  (reset                              )  //i
  );
  PEWSOS_255 pe_mat_14_11 (
    .io_in_r_data           (pe_mat_14_10_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pe_mat_14_10_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pe_mat_14_10_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pe_mat_14_10_io_out_r_stall        ), //i
    .io_out_r_data          (pe_mat_14_11_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_14_11_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_14_11_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_14_11_io_out_r_stall        ), //o
    .io_in_c_data           (pe_mat_13_11_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pe_mat_13_11_io_out_c_is_stationary), //i
    .io_out_c_data          (pe_mat_14_11_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_14_11_io_out_c_is_stationary), //o
    .clk                    (clk                                ), //i
    .reset                  (reset                              )  //i
  );
  PEWSOS_255 pe_mat_14_12 (
    .io_in_r_data           (pe_mat_14_11_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pe_mat_14_11_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pe_mat_14_11_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pe_mat_14_11_io_out_r_stall        ), //i
    .io_out_r_data          (pe_mat_14_12_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_14_12_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_14_12_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_14_12_io_out_r_stall        ), //o
    .io_in_c_data           (pe_mat_13_12_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pe_mat_13_12_io_out_c_is_stationary), //i
    .io_out_c_data          (pe_mat_14_12_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_14_12_io_out_c_is_stationary), //o
    .clk                    (clk                                ), //i
    .reset                  (reset                              )  //i
  );
  PEWSOS_255 pe_mat_14_13 (
    .io_in_r_data           (pe_mat_14_12_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pe_mat_14_12_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pe_mat_14_12_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pe_mat_14_12_io_out_r_stall        ), //i
    .io_out_r_data          (pe_mat_14_13_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_14_13_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_14_13_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_14_13_io_out_r_stall        ), //o
    .io_in_c_data           (pe_mat_13_13_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pe_mat_13_13_io_out_c_is_stationary), //i
    .io_out_c_data          (pe_mat_14_13_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_14_13_io_out_c_is_stationary), //o
    .clk                    (clk                                ), //i
    .reset                  (reset                              )  //i
  );
  PEWSOS_255 pe_mat_14_14 (
    .io_in_r_data           (pe_mat_14_13_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pe_mat_14_13_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pe_mat_14_13_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pe_mat_14_13_io_out_r_stall        ), //i
    .io_out_r_data          (pe_mat_14_14_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_14_14_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_14_14_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_14_14_io_out_r_stall        ), //o
    .io_in_c_data           (pe_mat_13_14_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pe_mat_13_14_io_out_c_is_stationary), //i
    .io_out_c_data          (pe_mat_14_14_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_14_14_io_out_c_is_stationary), //o
    .clk                    (clk                                ), //i
    .reset                  (reset                              )  //i
  );
  PEWSOS_255 pe_mat_14_15 (
    .io_in_r_data           (pe_mat_14_14_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pe_mat_14_14_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pe_mat_14_14_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pe_mat_14_14_io_out_r_stall        ), //i
    .io_out_r_data          (pe_mat_14_15_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_14_15_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_14_15_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_14_15_io_out_r_stall        ), //o
    .io_in_c_data           (pe_mat_13_15_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pe_mat_13_15_io_out_c_is_stationary), //i
    .io_out_c_data          (pe_mat_14_15_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_14_15_io_out_c_is_stationary), //o
    .clk                    (clk                                ), //i
    .reset                  (reset                              )  //i
  );
  PEWSOS_255 pe_mat_15_0 (
    .io_in_r_data           (io_in_r_15_data[15:0]             ), //i
    .io_in_r_load_store     (io_in_r_15_load_store             ), //i
    .io_in_r_df_is_ws       (io_in_r_15_df_is_ws               ), //i
    .io_in_r_stall          (io_in_r_15_stall                  ), //i
    .io_out_r_data          (pe_mat_15_0_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_15_0_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_15_0_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_15_0_io_out_r_stall        ), //o
    .io_in_c_data           (pe_mat_14_0_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pe_mat_14_0_io_out_c_is_stationary), //i
    .io_out_c_data          (pe_mat_15_0_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_15_0_io_out_c_is_stationary), //o
    .clk                    (clk                               ), //i
    .reset                  (reset                             )  //i
  );
  PEWSOS_255 pe_mat_15_1 (
    .io_in_r_data           (pe_mat_15_0_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pe_mat_15_0_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pe_mat_15_0_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pe_mat_15_0_io_out_r_stall        ), //i
    .io_out_r_data          (pe_mat_15_1_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_15_1_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_15_1_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_15_1_io_out_r_stall        ), //o
    .io_in_c_data           (pe_mat_14_1_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pe_mat_14_1_io_out_c_is_stationary), //i
    .io_out_c_data          (pe_mat_15_1_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_15_1_io_out_c_is_stationary), //o
    .clk                    (clk                               ), //i
    .reset                  (reset                             )  //i
  );
  PEWSOS_255 pe_mat_15_2 (
    .io_in_r_data           (pe_mat_15_1_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pe_mat_15_1_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pe_mat_15_1_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pe_mat_15_1_io_out_r_stall        ), //i
    .io_out_r_data          (pe_mat_15_2_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_15_2_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_15_2_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_15_2_io_out_r_stall        ), //o
    .io_in_c_data           (pe_mat_14_2_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pe_mat_14_2_io_out_c_is_stationary), //i
    .io_out_c_data          (pe_mat_15_2_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_15_2_io_out_c_is_stationary), //o
    .clk                    (clk                               ), //i
    .reset                  (reset                             )  //i
  );
  PEWSOS_255 pe_mat_15_3 (
    .io_in_r_data           (pe_mat_15_2_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pe_mat_15_2_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pe_mat_15_2_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pe_mat_15_2_io_out_r_stall        ), //i
    .io_out_r_data          (pe_mat_15_3_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_15_3_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_15_3_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_15_3_io_out_r_stall        ), //o
    .io_in_c_data           (pe_mat_14_3_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pe_mat_14_3_io_out_c_is_stationary), //i
    .io_out_c_data          (pe_mat_15_3_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_15_3_io_out_c_is_stationary), //o
    .clk                    (clk                               ), //i
    .reset                  (reset                             )  //i
  );
  PEWSOS_255 pe_mat_15_4 (
    .io_in_r_data           (pe_mat_15_3_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pe_mat_15_3_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pe_mat_15_3_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pe_mat_15_3_io_out_r_stall        ), //i
    .io_out_r_data          (pe_mat_15_4_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_15_4_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_15_4_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_15_4_io_out_r_stall        ), //o
    .io_in_c_data           (pe_mat_14_4_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pe_mat_14_4_io_out_c_is_stationary), //i
    .io_out_c_data          (pe_mat_15_4_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_15_4_io_out_c_is_stationary), //o
    .clk                    (clk                               ), //i
    .reset                  (reset                             )  //i
  );
  PEWSOS_255 pe_mat_15_5 (
    .io_in_r_data           (pe_mat_15_4_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pe_mat_15_4_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pe_mat_15_4_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pe_mat_15_4_io_out_r_stall        ), //i
    .io_out_r_data          (pe_mat_15_5_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_15_5_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_15_5_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_15_5_io_out_r_stall        ), //o
    .io_in_c_data           (pe_mat_14_5_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pe_mat_14_5_io_out_c_is_stationary), //i
    .io_out_c_data          (pe_mat_15_5_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_15_5_io_out_c_is_stationary), //o
    .clk                    (clk                               ), //i
    .reset                  (reset                             )  //i
  );
  PEWSOS_255 pe_mat_15_6 (
    .io_in_r_data           (pe_mat_15_5_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pe_mat_15_5_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pe_mat_15_5_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pe_mat_15_5_io_out_r_stall        ), //i
    .io_out_r_data          (pe_mat_15_6_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_15_6_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_15_6_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_15_6_io_out_r_stall        ), //o
    .io_in_c_data           (pe_mat_14_6_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pe_mat_14_6_io_out_c_is_stationary), //i
    .io_out_c_data          (pe_mat_15_6_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_15_6_io_out_c_is_stationary), //o
    .clk                    (clk                               ), //i
    .reset                  (reset                             )  //i
  );
  PEWSOS_255 pe_mat_15_7 (
    .io_in_r_data           (pe_mat_15_6_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pe_mat_15_6_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pe_mat_15_6_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pe_mat_15_6_io_out_r_stall        ), //i
    .io_out_r_data          (pe_mat_15_7_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_15_7_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_15_7_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_15_7_io_out_r_stall        ), //o
    .io_in_c_data           (pe_mat_14_7_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pe_mat_14_7_io_out_c_is_stationary), //i
    .io_out_c_data          (pe_mat_15_7_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_15_7_io_out_c_is_stationary), //o
    .clk                    (clk                               ), //i
    .reset                  (reset                             )  //i
  );
  PEWSOS_255 pe_mat_15_8 (
    .io_in_r_data           (pe_mat_15_7_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pe_mat_15_7_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pe_mat_15_7_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pe_mat_15_7_io_out_r_stall        ), //i
    .io_out_r_data          (pe_mat_15_8_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_15_8_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_15_8_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_15_8_io_out_r_stall        ), //o
    .io_in_c_data           (pe_mat_14_8_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pe_mat_14_8_io_out_c_is_stationary), //i
    .io_out_c_data          (pe_mat_15_8_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_15_8_io_out_c_is_stationary), //o
    .clk                    (clk                               ), //i
    .reset                  (reset                             )  //i
  );
  PEWSOS_255 pe_mat_15_9 (
    .io_in_r_data           (pe_mat_15_8_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pe_mat_15_8_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pe_mat_15_8_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pe_mat_15_8_io_out_r_stall        ), //i
    .io_out_r_data          (pe_mat_15_9_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_15_9_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_15_9_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_15_9_io_out_r_stall        ), //o
    .io_in_c_data           (pe_mat_14_9_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pe_mat_14_9_io_out_c_is_stationary), //i
    .io_out_c_data          (pe_mat_15_9_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_15_9_io_out_c_is_stationary), //o
    .clk                    (clk                               ), //i
    .reset                  (reset                             )  //i
  );
  PEWSOS_255 pe_mat_15_10 (
    .io_in_r_data           (pe_mat_15_9_io_out_r_data[15:0]    ), //i
    .io_in_r_load_store     (pe_mat_15_9_io_out_r_load_store    ), //i
    .io_in_r_df_is_ws       (pe_mat_15_9_io_out_r_df_is_ws      ), //i
    .io_in_r_stall          (pe_mat_15_9_io_out_r_stall         ), //i
    .io_out_r_data          (pe_mat_15_10_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_15_10_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_15_10_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_15_10_io_out_r_stall        ), //o
    .io_in_c_data           (pe_mat_14_10_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pe_mat_14_10_io_out_c_is_stationary), //i
    .io_out_c_data          (pe_mat_15_10_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_15_10_io_out_c_is_stationary), //o
    .clk                    (clk                                ), //i
    .reset                  (reset                              )  //i
  );
  PEWSOS_255 pe_mat_15_11 (
    .io_in_r_data           (pe_mat_15_10_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pe_mat_15_10_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pe_mat_15_10_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pe_mat_15_10_io_out_r_stall        ), //i
    .io_out_r_data          (pe_mat_15_11_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_15_11_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_15_11_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_15_11_io_out_r_stall        ), //o
    .io_in_c_data           (pe_mat_14_11_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pe_mat_14_11_io_out_c_is_stationary), //i
    .io_out_c_data          (pe_mat_15_11_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_15_11_io_out_c_is_stationary), //o
    .clk                    (clk                                ), //i
    .reset                  (reset                              )  //i
  );
  PEWSOS_255 pe_mat_15_12 (
    .io_in_r_data           (pe_mat_15_11_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pe_mat_15_11_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pe_mat_15_11_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pe_mat_15_11_io_out_r_stall        ), //i
    .io_out_r_data          (pe_mat_15_12_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_15_12_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_15_12_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_15_12_io_out_r_stall        ), //o
    .io_in_c_data           (pe_mat_14_12_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pe_mat_14_12_io_out_c_is_stationary), //i
    .io_out_c_data          (pe_mat_15_12_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_15_12_io_out_c_is_stationary), //o
    .clk                    (clk                                ), //i
    .reset                  (reset                              )  //i
  );
  PEWSOS_255 pe_mat_15_13 (
    .io_in_r_data           (pe_mat_15_12_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pe_mat_15_12_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pe_mat_15_12_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pe_mat_15_12_io_out_r_stall        ), //i
    .io_out_r_data          (pe_mat_15_13_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_15_13_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_15_13_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_15_13_io_out_r_stall        ), //o
    .io_in_c_data           (pe_mat_14_13_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pe_mat_14_13_io_out_c_is_stationary), //i
    .io_out_c_data          (pe_mat_15_13_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_15_13_io_out_c_is_stationary), //o
    .clk                    (clk                                ), //i
    .reset                  (reset                              )  //i
  );
  PEWSOS_255 pe_mat_15_14 (
    .io_in_r_data           (pe_mat_15_13_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pe_mat_15_13_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pe_mat_15_13_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pe_mat_15_13_io_out_r_stall        ), //i
    .io_out_r_data          (pe_mat_15_14_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_15_14_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_15_14_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_15_14_io_out_r_stall        ), //o
    .io_in_c_data           (pe_mat_14_14_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pe_mat_14_14_io_out_c_is_stationary), //i
    .io_out_c_data          (pe_mat_15_14_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_15_14_io_out_c_is_stationary), //o
    .clk                    (clk                                ), //i
    .reset                  (reset                              )  //i
  );
  PEWSOS_255 pe_mat_15_15 (
    .io_in_r_data           (pe_mat_15_14_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pe_mat_15_14_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pe_mat_15_14_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pe_mat_15_14_io_out_r_stall        ), //i
    .io_out_r_data          (pe_mat_15_15_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pe_mat_15_15_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pe_mat_15_15_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pe_mat_15_15_io_out_r_stall        ), //o
    .io_in_c_data           (pe_mat_14_15_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pe_mat_14_15_io_out_c_is_stationary), //i
    .io_out_c_data          (pe_mat_15_15_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pe_mat_15_15_io_out_c_is_stationary), //o
    .clk                    (clk                                ), //i
    .reset                  (reset                              )  //i
  );
  assign io_out_r_0_data = pe_mat_0_15_io_out_r_data; // @[SystolicConnect.scala 50:16]
  assign io_out_r_0_load_store = pe_mat_0_15_io_out_r_load_store; // @[SystolicConnect.scala 50:16]
  assign io_out_r_0_df_is_ws = pe_mat_0_15_io_out_r_df_is_ws; // @[SystolicConnect.scala 50:16]
  assign io_out_r_0_stall = pe_mat_0_15_io_out_r_stall; // @[SystolicConnect.scala 50:16]
  assign io_out_r_1_data = pe_mat_1_15_io_out_r_data; // @[SystolicConnect.scala 50:16]
  assign io_out_r_1_load_store = pe_mat_1_15_io_out_r_load_store; // @[SystolicConnect.scala 50:16]
  assign io_out_r_1_df_is_ws = pe_mat_1_15_io_out_r_df_is_ws; // @[SystolicConnect.scala 50:16]
  assign io_out_r_1_stall = pe_mat_1_15_io_out_r_stall; // @[SystolicConnect.scala 50:16]
  assign io_out_r_2_data = pe_mat_2_15_io_out_r_data; // @[SystolicConnect.scala 50:16]
  assign io_out_r_2_load_store = pe_mat_2_15_io_out_r_load_store; // @[SystolicConnect.scala 50:16]
  assign io_out_r_2_df_is_ws = pe_mat_2_15_io_out_r_df_is_ws; // @[SystolicConnect.scala 50:16]
  assign io_out_r_2_stall = pe_mat_2_15_io_out_r_stall; // @[SystolicConnect.scala 50:16]
  assign io_out_r_3_data = pe_mat_3_15_io_out_r_data; // @[SystolicConnect.scala 50:16]
  assign io_out_r_3_load_store = pe_mat_3_15_io_out_r_load_store; // @[SystolicConnect.scala 50:16]
  assign io_out_r_3_df_is_ws = pe_mat_3_15_io_out_r_df_is_ws; // @[SystolicConnect.scala 50:16]
  assign io_out_r_3_stall = pe_mat_3_15_io_out_r_stall; // @[SystolicConnect.scala 50:16]
  assign io_out_r_4_data = pe_mat_4_15_io_out_r_data; // @[SystolicConnect.scala 50:16]
  assign io_out_r_4_load_store = pe_mat_4_15_io_out_r_load_store; // @[SystolicConnect.scala 50:16]
  assign io_out_r_4_df_is_ws = pe_mat_4_15_io_out_r_df_is_ws; // @[SystolicConnect.scala 50:16]
  assign io_out_r_4_stall = pe_mat_4_15_io_out_r_stall; // @[SystolicConnect.scala 50:16]
  assign io_out_r_5_data = pe_mat_5_15_io_out_r_data; // @[SystolicConnect.scala 50:16]
  assign io_out_r_5_load_store = pe_mat_5_15_io_out_r_load_store; // @[SystolicConnect.scala 50:16]
  assign io_out_r_5_df_is_ws = pe_mat_5_15_io_out_r_df_is_ws; // @[SystolicConnect.scala 50:16]
  assign io_out_r_5_stall = pe_mat_5_15_io_out_r_stall; // @[SystolicConnect.scala 50:16]
  assign io_out_r_6_data = pe_mat_6_15_io_out_r_data; // @[SystolicConnect.scala 50:16]
  assign io_out_r_6_load_store = pe_mat_6_15_io_out_r_load_store; // @[SystolicConnect.scala 50:16]
  assign io_out_r_6_df_is_ws = pe_mat_6_15_io_out_r_df_is_ws; // @[SystolicConnect.scala 50:16]
  assign io_out_r_6_stall = pe_mat_6_15_io_out_r_stall; // @[SystolicConnect.scala 50:16]
  assign io_out_r_7_data = pe_mat_7_15_io_out_r_data; // @[SystolicConnect.scala 50:16]
  assign io_out_r_7_load_store = pe_mat_7_15_io_out_r_load_store; // @[SystolicConnect.scala 50:16]
  assign io_out_r_7_df_is_ws = pe_mat_7_15_io_out_r_df_is_ws; // @[SystolicConnect.scala 50:16]
  assign io_out_r_7_stall = pe_mat_7_15_io_out_r_stall; // @[SystolicConnect.scala 50:16]
  assign io_out_r_8_data = pe_mat_8_15_io_out_r_data; // @[SystolicConnect.scala 50:16]
  assign io_out_r_8_load_store = pe_mat_8_15_io_out_r_load_store; // @[SystolicConnect.scala 50:16]
  assign io_out_r_8_df_is_ws = pe_mat_8_15_io_out_r_df_is_ws; // @[SystolicConnect.scala 50:16]
  assign io_out_r_8_stall = pe_mat_8_15_io_out_r_stall; // @[SystolicConnect.scala 50:16]
  assign io_out_r_9_data = pe_mat_9_15_io_out_r_data; // @[SystolicConnect.scala 50:16]
  assign io_out_r_9_load_store = pe_mat_9_15_io_out_r_load_store; // @[SystolicConnect.scala 50:16]
  assign io_out_r_9_df_is_ws = pe_mat_9_15_io_out_r_df_is_ws; // @[SystolicConnect.scala 50:16]
  assign io_out_r_9_stall = pe_mat_9_15_io_out_r_stall; // @[SystolicConnect.scala 50:16]
  assign io_out_r_10_data = pe_mat_10_15_io_out_r_data; // @[SystolicConnect.scala 50:16]
  assign io_out_r_10_load_store = pe_mat_10_15_io_out_r_load_store; // @[SystolicConnect.scala 50:16]
  assign io_out_r_10_df_is_ws = pe_mat_10_15_io_out_r_df_is_ws; // @[SystolicConnect.scala 50:16]
  assign io_out_r_10_stall = pe_mat_10_15_io_out_r_stall; // @[SystolicConnect.scala 50:16]
  assign io_out_r_11_data = pe_mat_11_15_io_out_r_data; // @[SystolicConnect.scala 50:16]
  assign io_out_r_11_load_store = pe_mat_11_15_io_out_r_load_store; // @[SystolicConnect.scala 50:16]
  assign io_out_r_11_df_is_ws = pe_mat_11_15_io_out_r_df_is_ws; // @[SystolicConnect.scala 50:16]
  assign io_out_r_11_stall = pe_mat_11_15_io_out_r_stall; // @[SystolicConnect.scala 50:16]
  assign io_out_r_12_data = pe_mat_12_15_io_out_r_data; // @[SystolicConnect.scala 50:16]
  assign io_out_r_12_load_store = pe_mat_12_15_io_out_r_load_store; // @[SystolicConnect.scala 50:16]
  assign io_out_r_12_df_is_ws = pe_mat_12_15_io_out_r_df_is_ws; // @[SystolicConnect.scala 50:16]
  assign io_out_r_12_stall = pe_mat_12_15_io_out_r_stall; // @[SystolicConnect.scala 50:16]
  assign io_out_r_13_data = pe_mat_13_15_io_out_r_data; // @[SystolicConnect.scala 50:16]
  assign io_out_r_13_load_store = pe_mat_13_15_io_out_r_load_store; // @[SystolicConnect.scala 50:16]
  assign io_out_r_13_df_is_ws = pe_mat_13_15_io_out_r_df_is_ws; // @[SystolicConnect.scala 50:16]
  assign io_out_r_13_stall = pe_mat_13_15_io_out_r_stall; // @[SystolicConnect.scala 50:16]
  assign io_out_r_14_data = pe_mat_14_15_io_out_r_data; // @[SystolicConnect.scala 50:16]
  assign io_out_r_14_load_store = pe_mat_14_15_io_out_r_load_store; // @[SystolicConnect.scala 50:16]
  assign io_out_r_14_df_is_ws = pe_mat_14_15_io_out_r_df_is_ws; // @[SystolicConnect.scala 50:16]
  assign io_out_r_14_stall = pe_mat_14_15_io_out_r_stall; // @[SystolicConnect.scala 50:16]
  assign io_out_r_15_data = pe_mat_15_15_io_out_r_data; // @[SystolicConnect.scala 50:16]
  assign io_out_r_15_load_store = pe_mat_15_15_io_out_r_load_store; // @[SystolicConnect.scala 50:16]
  assign io_out_r_15_df_is_ws = pe_mat_15_15_io_out_r_df_is_ws; // @[SystolicConnect.scala 50:16]
  assign io_out_r_15_stall = pe_mat_15_15_io_out_r_stall; // @[SystolicConnect.scala 50:16]
  assign io_out_c_0_data = pe_mat_15_0_io_out_c_data; // @[SystolicConnect.scala 56:16]
  assign io_out_c_0_is_stationary = pe_mat_15_0_io_out_c_is_stationary; // @[SystolicConnect.scala 56:16]
  assign io_out_c_1_data = pe_mat_15_1_io_out_c_data; // @[SystolicConnect.scala 56:16]
  assign io_out_c_1_is_stationary = pe_mat_15_1_io_out_c_is_stationary; // @[SystolicConnect.scala 56:16]
  assign io_out_c_2_data = pe_mat_15_2_io_out_c_data; // @[SystolicConnect.scala 56:16]
  assign io_out_c_2_is_stationary = pe_mat_15_2_io_out_c_is_stationary; // @[SystolicConnect.scala 56:16]
  assign io_out_c_3_data = pe_mat_15_3_io_out_c_data; // @[SystolicConnect.scala 56:16]
  assign io_out_c_3_is_stationary = pe_mat_15_3_io_out_c_is_stationary; // @[SystolicConnect.scala 56:16]
  assign io_out_c_4_data = pe_mat_15_4_io_out_c_data; // @[SystolicConnect.scala 56:16]
  assign io_out_c_4_is_stationary = pe_mat_15_4_io_out_c_is_stationary; // @[SystolicConnect.scala 56:16]
  assign io_out_c_5_data = pe_mat_15_5_io_out_c_data; // @[SystolicConnect.scala 56:16]
  assign io_out_c_5_is_stationary = pe_mat_15_5_io_out_c_is_stationary; // @[SystolicConnect.scala 56:16]
  assign io_out_c_6_data = pe_mat_15_6_io_out_c_data; // @[SystolicConnect.scala 56:16]
  assign io_out_c_6_is_stationary = pe_mat_15_6_io_out_c_is_stationary; // @[SystolicConnect.scala 56:16]
  assign io_out_c_7_data = pe_mat_15_7_io_out_c_data; // @[SystolicConnect.scala 56:16]
  assign io_out_c_7_is_stationary = pe_mat_15_7_io_out_c_is_stationary; // @[SystolicConnect.scala 56:16]
  assign io_out_c_8_data = pe_mat_15_8_io_out_c_data; // @[SystolicConnect.scala 56:16]
  assign io_out_c_8_is_stationary = pe_mat_15_8_io_out_c_is_stationary; // @[SystolicConnect.scala 56:16]
  assign io_out_c_9_data = pe_mat_15_9_io_out_c_data; // @[SystolicConnect.scala 56:16]
  assign io_out_c_9_is_stationary = pe_mat_15_9_io_out_c_is_stationary; // @[SystolicConnect.scala 56:16]
  assign io_out_c_10_data = pe_mat_15_10_io_out_c_data; // @[SystolicConnect.scala 56:16]
  assign io_out_c_10_is_stationary = pe_mat_15_10_io_out_c_is_stationary; // @[SystolicConnect.scala 56:16]
  assign io_out_c_11_data = pe_mat_15_11_io_out_c_data; // @[SystolicConnect.scala 56:16]
  assign io_out_c_11_is_stationary = pe_mat_15_11_io_out_c_is_stationary; // @[SystolicConnect.scala 56:16]
  assign io_out_c_12_data = pe_mat_15_12_io_out_c_data; // @[SystolicConnect.scala 56:16]
  assign io_out_c_12_is_stationary = pe_mat_15_12_io_out_c_is_stationary; // @[SystolicConnect.scala 56:16]
  assign io_out_c_13_data = pe_mat_15_13_io_out_c_data; // @[SystolicConnect.scala 56:16]
  assign io_out_c_13_is_stationary = pe_mat_15_13_io_out_c_is_stationary; // @[SystolicConnect.scala 56:16]
  assign io_out_c_14_data = pe_mat_15_14_io_out_c_data; // @[SystolicConnect.scala 56:16]
  assign io_out_c_14_is_stationary = pe_mat_15_14_io_out_c_is_stationary; // @[SystolicConnect.scala 56:16]
  assign io_out_c_15_data = pe_mat_15_15_io_out_c_data; // @[SystolicConnect.scala 56:16]
  assign io_out_c_15_is_stationary = pe_mat_15_15_io_out_c_is_stationary; // @[SystolicConnect.scala 56:16]

endmodule

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

//PEWSOS_255 replaced by PEWSOS_255

module PEWSOS_255 (
  input      [15:0]   io_in_r_data,
  input               io_in_r_load_store,
  input               io_in_r_df_is_ws,
  input               io_in_r_stall,
  output     [15:0]   io_out_r_data,
  output              io_out_r_load_store,
  output              io_out_r_df_is_ws,
  output              io_out_r_stall,
  input      [15:0]   io_in_c_data,
  input               io_in_c_is_stationary,
  output     [15:0]   io_out_c_data,
  output              io_out_c_is_stationary,
  input               clk,
  input               reset
);

  wire       [15:0]   mac_256_io_psum;
  wire       [15:0]   mac_256_io_weight;
  wire       [15:0]   mac_256_io_result;
  wire                not_stall;
  wire       [15:0]   mac_result;
  reg        [15:0]   stationary;
  reg                 stationary_en;
  wire                when_PEWSOS_l68;
  reg        [15:0]   stationary_reg;
  reg                 io_in_r_stall_regNext;
  reg        [15:0]   io_in_r_data_regNextWhen;
  reg                 io_in_r_load_store_regNextWhen;
  reg                 io_in_r_df_is_ws_regNextWhen;
  reg        [15:0]   out_c_data;
  reg                 out_c_is_stationary;
  wire                when_PEWSOS_l87;
  wire                when_PEWSOS_l95;
  reg        [15:0]   out_c_data_regNextWhen;
  reg                 out_c_is_stationary_regNextWhen;

  Mac_255 mac_256 (
    .io_psum            (mac_256_io_psum[15:0]  ), //i
    .io_weight          (mac_256_io_weight[15:0]), //i
    .io_inputActivation (io_in_r_data[15:0]     ), //i
    .io_result          (mac_256_io_result[15:0])  //o
  );
  assign not_stall = (! io_in_r_stall); // @[BaseType.scala 299:24]
  always @(*) begin
    if(io_in_r_df_is_ws) begin
      stationary = io_in_c_data; // @[PEWSOS.scala 57:16]
    end else begin
      if(io_in_c_is_stationary) begin
        stationary = 16'h0; // @[PEWSOS.scala 61:18]
      end else begin
        stationary = mac_result; // @[PEWSOS.scala 64:18]
      end
    end
  end

  always @(*) begin
    if(io_in_r_df_is_ws) begin
      stationary_en = io_in_r_load_store; // @[PEWSOS.scala 58:19]
    end else begin
      if(io_in_c_is_stationary) begin
        stationary_en = io_in_r_load_store; // @[PEWSOS.scala 62:21]
      end else begin
        stationary_en = 1'b1; // @[PEWSOS.scala 65:21]
      end
    end
  end

  assign when_PEWSOS_l68 = (stationary_en && not_stall); // @[BaseType.scala 305:24]
  assign mac_256_io_psum = (io_in_r_df_is_ws ? io_in_c_data : stationary_reg); // @[PEWSOS.scala 72:15]
  assign mac_256_io_weight = (io_in_r_df_is_ws ? stationary_reg : io_in_c_data); // @[PEWSOS.scala 73:17]
  assign mac_result = mac_256_io_result; // @[PEWSOS.scala 75:14]
  assign io_out_r_stall = io_in_r_stall_regNext; // @[PEWSOS.scala 78:18]
  assign io_out_r_data = io_in_r_data_regNextWhen; // @[PEWSOS.scala 79:17]
  assign io_out_r_load_store = io_in_r_load_store_regNextWhen; // @[PEWSOS.scala 80:23]
  assign io_out_r_df_is_ws = io_in_r_df_is_ws_regNextWhen; // @[PEWSOS.scala 81:21]
  assign when_PEWSOS_l87 = (io_in_c_is_stationary && (! io_in_r_load_store)); // @[BaseType.scala 305:24]
  always @(*) begin
    if(io_in_r_df_is_ws) begin
      if(when_PEWSOS_l87) begin
        out_c_data = io_in_c_data; // @[PEWSOS.scala 88:18]
      end else begin
        out_c_data = mac_result; // @[PEWSOS.scala 91:18]
      end
    end else begin
      if(when_PEWSOS_l95) begin
        out_c_data = io_in_c_data; // @[PEWSOS.scala 96:18]
      end else begin
        if(io_in_r_load_store) begin
          out_c_data = stationary_reg; // @[PEWSOS.scala 99:18]
        end else begin
          out_c_data = io_in_c_data; // @[PEWSOS.scala 102:18]
        end
      end
    end
  end

  always @(*) begin
    if(io_in_r_df_is_ws) begin
      if(when_PEWSOS_l87) begin
        out_c_is_stationary = 1'b1; // @[PEWSOS.scala 89:27]
      end else begin
        out_c_is_stationary = 1'b0; // @[PEWSOS.scala 92:27]
      end
    end else begin
      if(when_PEWSOS_l95) begin
        out_c_is_stationary = 1'b1; // @[PEWSOS.scala 97:27]
      end else begin
        if(io_in_r_load_store) begin
          out_c_is_stationary = 1'b1; // @[PEWSOS.scala 100:27]
        end else begin
          out_c_is_stationary = 1'b0; // @[PEWSOS.scala 103:27]
        end
      end
    end
  end

  assign when_PEWSOS_l95 = (io_in_c_is_stationary && (! io_in_r_load_store)); // @[BaseType.scala 305:24]
  assign io_out_c_data = out_c_data_regNextWhen; // @[PEWSOS.scala 106:17]
  assign io_out_c_is_stationary = out_c_is_stationary_regNextWhen; // @[PEWSOS.scala 107:26]
  always @(posedge clk) begin
    if(when_PEWSOS_l68) begin
      stationary_reg <= stationary; // @[PEWSOS.scala 68:35]
    end
    io_in_r_stall_regNext <= io_in_r_stall; // @[Reg.scala 39:30]
    if(not_stall) begin
      io_in_r_data_regNextWhen <= io_in_r_data; // @[PEWSOS.scala 79:31]
    end
    if(not_stall) begin
      io_in_r_load_store_regNextWhen <= io_in_r_load_store; // @[PEWSOS.scala 80:37]
    end
    if(not_stall) begin
      io_in_r_df_is_ws_regNextWhen <= io_in_r_df_is_ws; // @[PEWSOS.scala 81:35]
    end
    if(not_stall) begin
      out_c_data_regNextWhen <= out_c_data; // @[PEWSOS.scala 106:31]
    end
    if(not_stall) begin
      out_c_is_stationary_regNextWhen <= out_c_is_stationary; // @[PEWSOS.scala 107:40]
    end
  end


endmodule

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

//Mac_255 replaced by Mac_255

module Mac_255 (
  input      [15:0]   io_psum,
  input      [15:0]   io_weight,
  input      [15:0]   io_inputActivation,
  output     [15:0]   io_result
);

  wire       [31:0]   _zz_io_result;
  wire       [31:0]   _zz_io_result_1;
  wire       [31:0]   _zz_io_result_2;

  assign _zz_io_result = ($signed(_zz_io_result_1) + $signed(_zz_io_result_2));
  assign _zz_io_result_1 = ($signed(io_inputActivation) * $signed(io_weight));
  assign _zz_io_result_2 = {{16{io_psum[15]}}, io_psum};
  assign io_result = _zz_io_result[15:0]; // @[Mac.scala 14:31]

endmodule
