// Generator : SpinalHDL v1.8.0    git head : 4e3563a282582b41f4eaafc503787757251d23ea
// Component : ArraySARA
// Git hash  : aeab30821bf33dec846c2049cebcf2d24a28afa4

`timescale 1ns/1ps

module ArraySARA (
  input      [15:0]   io_in_r_0_data_0_data,
  input               io_in_r_0_data_0_load_store,
  input               io_in_r_0_data_0_df_is_ws,
  input               io_in_r_0_data_0_stall,
  input      [15:0]   io_in_r_0_data_1_data,
  input               io_in_r_0_data_1_load_store,
  input               io_in_r_0_data_1_df_is_ws,
  input               io_in_r_0_data_1_stall,
  input      [15:0]   io_in_r_0_data_2_data,
  input               io_in_r_0_data_2_load_store,
  input               io_in_r_0_data_2_df_is_ws,
  input               io_in_r_0_data_2_stall,
  input      [15:0]   io_in_r_0_data_3_data,
  input               io_in_r_0_data_3_load_store,
  input               io_in_r_0_data_3_df_is_ws,
  input               io_in_r_0_data_3_stall,
  input      [15:0]   io_in_r_0_bypass_0_0_data,
  input               io_in_r_0_bypass_0_0_load_store,
  input               io_in_r_0_bypass_0_0_df_is_ws,
  input               io_in_r_0_bypass_0_0_stall,
  input      [15:0]   io_in_r_0_bypass_0_1_data,
  input               io_in_r_0_bypass_0_1_load_store,
  input               io_in_r_0_bypass_0_1_df_is_ws,
  input               io_in_r_0_bypass_0_1_stall,
  input      [15:0]   io_in_r_0_bypass_0_2_data,
  input               io_in_r_0_bypass_0_2_load_store,
  input               io_in_r_0_bypass_0_2_df_is_ws,
  input               io_in_r_0_bypass_0_2_stall,
  input      [15:0]   io_in_r_0_bypass_0_3_data,
  input               io_in_r_0_bypass_0_3_load_store,
  input               io_in_r_0_bypass_0_3_df_is_ws,
  input               io_in_r_0_bypass_0_3_stall,
  input      [15:0]   io_in_r_0_bypass_1_0_data,
  input               io_in_r_0_bypass_1_0_load_store,
  input               io_in_r_0_bypass_1_0_df_is_ws,
  input               io_in_r_0_bypass_1_0_stall,
  input      [15:0]   io_in_r_0_bypass_1_1_data,
  input               io_in_r_0_bypass_1_1_load_store,
  input               io_in_r_0_bypass_1_1_df_is_ws,
  input               io_in_r_0_bypass_1_1_stall,
  input      [15:0]   io_in_r_0_bypass_1_2_data,
  input               io_in_r_0_bypass_1_2_load_store,
  input               io_in_r_0_bypass_1_2_df_is_ws,
  input               io_in_r_0_bypass_1_2_stall,
  input      [15:0]   io_in_r_0_bypass_1_3_data,
  input               io_in_r_0_bypass_1_3_load_store,
  input               io_in_r_0_bypass_1_3_df_is_ws,
  input               io_in_r_0_bypass_1_3_stall,
  input               io_in_r_0_input_from_bypass_0,
  input               io_in_r_0_input_from_bypass_1,
  input      [15:0]   io_in_r_1_data_0_data,
  input               io_in_r_1_data_0_load_store,
  input               io_in_r_1_data_0_df_is_ws,
  input               io_in_r_1_data_0_stall,
  input      [15:0]   io_in_r_1_data_1_data,
  input               io_in_r_1_data_1_load_store,
  input               io_in_r_1_data_1_df_is_ws,
  input               io_in_r_1_data_1_stall,
  input      [15:0]   io_in_r_1_data_2_data,
  input               io_in_r_1_data_2_load_store,
  input               io_in_r_1_data_2_df_is_ws,
  input               io_in_r_1_data_2_stall,
  input      [15:0]   io_in_r_1_data_3_data,
  input               io_in_r_1_data_3_load_store,
  input               io_in_r_1_data_3_df_is_ws,
  input               io_in_r_1_data_3_stall,
  input      [15:0]   io_in_r_1_bypass_0_0_data,
  input               io_in_r_1_bypass_0_0_load_store,
  input               io_in_r_1_bypass_0_0_df_is_ws,
  input               io_in_r_1_bypass_0_0_stall,
  input      [15:0]   io_in_r_1_bypass_0_1_data,
  input               io_in_r_1_bypass_0_1_load_store,
  input               io_in_r_1_bypass_0_1_df_is_ws,
  input               io_in_r_1_bypass_0_1_stall,
  input      [15:0]   io_in_r_1_bypass_0_2_data,
  input               io_in_r_1_bypass_0_2_load_store,
  input               io_in_r_1_bypass_0_2_df_is_ws,
  input               io_in_r_1_bypass_0_2_stall,
  input      [15:0]   io_in_r_1_bypass_0_3_data,
  input               io_in_r_1_bypass_0_3_load_store,
  input               io_in_r_1_bypass_0_3_df_is_ws,
  input               io_in_r_1_bypass_0_3_stall,
  input      [15:0]   io_in_r_1_bypass_1_0_data,
  input               io_in_r_1_bypass_1_0_load_store,
  input               io_in_r_1_bypass_1_0_df_is_ws,
  input               io_in_r_1_bypass_1_0_stall,
  input      [15:0]   io_in_r_1_bypass_1_1_data,
  input               io_in_r_1_bypass_1_1_load_store,
  input               io_in_r_1_bypass_1_1_df_is_ws,
  input               io_in_r_1_bypass_1_1_stall,
  input      [15:0]   io_in_r_1_bypass_1_2_data,
  input               io_in_r_1_bypass_1_2_load_store,
  input               io_in_r_1_bypass_1_2_df_is_ws,
  input               io_in_r_1_bypass_1_2_stall,
  input      [15:0]   io_in_r_1_bypass_1_3_data,
  input               io_in_r_1_bypass_1_3_load_store,
  input               io_in_r_1_bypass_1_3_df_is_ws,
  input               io_in_r_1_bypass_1_3_stall,
  input               io_in_r_1_input_from_bypass_0,
  input               io_in_r_1_input_from_bypass_1,
  output     [15:0]   io_out_r_0_data_0_data,
  output              io_out_r_0_data_0_load_store,
  output              io_out_r_0_data_0_df_is_ws,
  output              io_out_r_0_data_0_stall,
  output     [15:0]   io_out_r_0_data_1_data,
  output              io_out_r_0_data_1_load_store,
  output              io_out_r_0_data_1_df_is_ws,
  output              io_out_r_0_data_1_stall,
  output     [15:0]   io_out_r_0_data_2_data,
  output              io_out_r_0_data_2_load_store,
  output              io_out_r_0_data_2_df_is_ws,
  output              io_out_r_0_data_2_stall,
  output     [15:0]   io_out_r_0_data_3_data,
  output              io_out_r_0_data_3_load_store,
  output              io_out_r_0_data_3_df_is_ws,
  output              io_out_r_0_data_3_stall,
  output     [15:0]   io_out_r_0_bypass_0_0_data,
  output              io_out_r_0_bypass_0_0_load_store,
  output              io_out_r_0_bypass_0_0_df_is_ws,
  output              io_out_r_0_bypass_0_0_stall,
  output     [15:0]   io_out_r_0_bypass_0_1_data,
  output              io_out_r_0_bypass_0_1_load_store,
  output              io_out_r_0_bypass_0_1_df_is_ws,
  output              io_out_r_0_bypass_0_1_stall,
  output     [15:0]   io_out_r_0_bypass_0_2_data,
  output              io_out_r_0_bypass_0_2_load_store,
  output              io_out_r_0_bypass_0_2_df_is_ws,
  output              io_out_r_0_bypass_0_2_stall,
  output     [15:0]   io_out_r_0_bypass_0_3_data,
  output              io_out_r_0_bypass_0_3_load_store,
  output              io_out_r_0_bypass_0_3_df_is_ws,
  output              io_out_r_0_bypass_0_3_stall,
  output     [15:0]   io_out_r_0_bypass_1_0_data,
  output              io_out_r_0_bypass_1_0_load_store,
  output              io_out_r_0_bypass_1_0_df_is_ws,
  output              io_out_r_0_bypass_1_0_stall,
  output     [15:0]   io_out_r_0_bypass_1_1_data,
  output              io_out_r_0_bypass_1_1_load_store,
  output              io_out_r_0_bypass_1_1_df_is_ws,
  output              io_out_r_0_bypass_1_1_stall,
  output     [15:0]   io_out_r_0_bypass_1_2_data,
  output              io_out_r_0_bypass_1_2_load_store,
  output              io_out_r_0_bypass_1_2_df_is_ws,
  output              io_out_r_0_bypass_1_2_stall,
  output     [15:0]   io_out_r_0_bypass_1_3_data,
  output              io_out_r_0_bypass_1_3_load_store,
  output              io_out_r_0_bypass_1_3_df_is_ws,
  output              io_out_r_0_bypass_1_3_stall,
  output              io_out_r_0_input_from_bypass_0,
  output              io_out_r_0_input_from_bypass_1,
  output     [15:0]   io_out_r_1_data_0_data,
  output              io_out_r_1_data_0_load_store,
  output              io_out_r_1_data_0_df_is_ws,
  output              io_out_r_1_data_0_stall,
  output     [15:0]   io_out_r_1_data_1_data,
  output              io_out_r_1_data_1_load_store,
  output              io_out_r_1_data_1_df_is_ws,
  output              io_out_r_1_data_1_stall,
  output     [15:0]   io_out_r_1_data_2_data,
  output              io_out_r_1_data_2_load_store,
  output              io_out_r_1_data_2_df_is_ws,
  output              io_out_r_1_data_2_stall,
  output     [15:0]   io_out_r_1_data_3_data,
  output              io_out_r_1_data_3_load_store,
  output              io_out_r_1_data_3_df_is_ws,
  output              io_out_r_1_data_3_stall,
  output     [15:0]   io_out_r_1_bypass_0_0_data,
  output              io_out_r_1_bypass_0_0_load_store,
  output              io_out_r_1_bypass_0_0_df_is_ws,
  output              io_out_r_1_bypass_0_0_stall,
  output     [15:0]   io_out_r_1_bypass_0_1_data,
  output              io_out_r_1_bypass_0_1_load_store,
  output              io_out_r_1_bypass_0_1_df_is_ws,
  output              io_out_r_1_bypass_0_1_stall,
  output     [15:0]   io_out_r_1_bypass_0_2_data,
  output              io_out_r_1_bypass_0_2_load_store,
  output              io_out_r_1_bypass_0_2_df_is_ws,
  output              io_out_r_1_bypass_0_2_stall,
  output     [15:0]   io_out_r_1_bypass_0_3_data,
  output              io_out_r_1_bypass_0_3_load_store,
  output              io_out_r_1_bypass_0_3_df_is_ws,
  output              io_out_r_1_bypass_0_3_stall,
  output     [15:0]   io_out_r_1_bypass_1_0_data,
  output              io_out_r_1_bypass_1_0_load_store,
  output              io_out_r_1_bypass_1_0_df_is_ws,
  output              io_out_r_1_bypass_1_0_stall,
  output     [15:0]   io_out_r_1_bypass_1_1_data,
  output              io_out_r_1_bypass_1_1_load_store,
  output              io_out_r_1_bypass_1_1_df_is_ws,
  output              io_out_r_1_bypass_1_1_stall,
  output     [15:0]   io_out_r_1_bypass_1_2_data,
  output              io_out_r_1_bypass_1_2_load_store,
  output              io_out_r_1_bypass_1_2_df_is_ws,
  output              io_out_r_1_bypass_1_2_stall,
  output     [15:0]   io_out_r_1_bypass_1_3_data,
  output              io_out_r_1_bypass_1_3_load_store,
  output              io_out_r_1_bypass_1_3_df_is_ws,
  output              io_out_r_1_bypass_1_3_stall,
  output              io_out_r_1_input_from_bypass_0,
  output              io_out_r_1_input_from_bypass_1,
  input      [15:0]   io_in_c_0_data_0_data,
  input               io_in_c_0_data_0_is_stationary,
  input      [15:0]   io_in_c_0_data_1_data,
  input               io_in_c_0_data_1_is_stationary,
  input      [15:0]   io_in_c_0_data_2_data,
  input               io_in_c_0_data_2_is_stationary,
  input      [15:0]   io_in_c_0_data_3_data,
  input               io_in_c_0_data_3_is_stationary,
  input      [15:0]   io_in_c_0_bypass_0_0_data,
  input               io_in_c_0_bypass_0_0_is_stationary,
  input      [15:0]   io_in_c_0_bypass_0_1_data,
  input               io_in_c_0_bypass_0_1_is_stationary,
  input      [15:0]   io_in_c_0_bypass_0_2_data,
  input               io_in_c_0_bypass_0_2_is_stationary,
  input      [15:0]   io_in_c_0_bypass_0_3_data,
  input               io_in_c_0_bypass_0_3_is_stationary,
  input      [15:0]   io_in_c_0_bypass_1_0_data,
  input               io_in_c_0_bypass_1_0_is_stationary,
  input      [15:0]   io_in_c_0_bypass_1_1_data,
  input               io_in_c_0_bypass_1_1_is_stationary,
  input      [15:0]   io_in_c_0_bypass_1_2_data,
  input               io_in_c_0_bypass_1_2_is_stationary,
  input      [15:0]   io_in_c_0_bypass_1_3_data,
  input               io_in_c_0_bypass_1_3_is_stationary,
  input               io_in_c_0_input_from_bypass_0,
  input               io_in_c_0_input_from_bypass_1,
  input      [15:0]   io_in_c_1_data_0_data,
  input               io_in_c_1_data_0_is_stationary,
  input      [15:0]   io_in_c_1_data_1_data,
  input               io_in_c_1_data_1_is_stationary,
  input      [15:0]   io_in_c_1_data_2_data,
  input               io_in_c_1_data_2_is_stationary,
  input      [15:0]   io_in_c_1_data_3_data,
  input               io_in_c_1_data_3_is_stationary,
  input      [15:0]   io_in_c_1_bypass_0_0_data,
  input               io_in_c_1_bypass_0_0_is_stationary,
  input      [15:0]   io_in_c_1_bypass_0_1_data,
  input               io_in_c_1_bypass_0_1_is_stationary,
  input      [15:0]   io_in_c_1_bypass_0_2_data,
  input               io_in_c_1_bypass_0_2_is_stationary,
  input      [15:0]   io_in_c_1_bypass_0_3_data,
  input               io_in_c_1_bypass_0_3_is_stationary,
  input      [15:0]   io_in_c_1_bypass_1_0_data,
  input               io_in_c_1_bypass_1_0_is_stationary,
  input      [15:0]   io_in_c_1_bypass_1_1_data,
  input               io_in_c_1_bypass_1_1_is_stationary,
  input      [15:0]   io_in_c_1_bypass_1_2_data,
  input               io_in_c_1_bypass_1_2_is_stationary,
  input      [15:0]   io_in_c_1_bypass_1_3_data,
  input               io_in_c_1_bypass_1_3_is_stationary,
  input               io_in_c_1_input_from_bypass_0,
  input               io_in_c_1_input_from_bypass_1,
  output     [15:0]   io_out_c_0_data_0_data,
  output              io_out_c_0_data_0_is_stationary,
  output     [15:0]   io_out_c_0_data_1_data,
  output              io_out_c_0_data_1_is_stationary,
  output     [15:0]   io_out_c_0_data_2_data,
  output              io_out_c_0_data_2_is_stationary,
  output     [15:0]   io_out_c_0_data_3_data,
  output              io_out_c_0_data_3_is_stationary,
  output     [15:0]   io_out_c_0_bypass_0_0_data,
  output              io_out_c_0_bypass_0_0_is_stationary,
  output     [15:0]   io_out_c_0_bypass_0_1_data,
  output              io_out_c_0_bypass_0_1_is_stationary,
  output     [15:0]   io_out_c_0_bypass_0_2_data,
  output              io_out_c_0_bypass_0_2_is_stationary,
  output     [15:0]   io_out_c_0_bypass_0_3_data,
  output              io_out_c_0_bypass_0_3_is_stationary,
  output     [15:0]   io_out_c_0_bypass_1_0_data,
  output              io_out_c_0_bypass_1_0_is_stationary,
  output     [15:0]   io_out_c_0_bypass_1_1_data,
  output              io_out_c_0_bypass_1_1_is_stationary,
  output     [15:0]   io_out_c_0_bypass_1_2_data,
  output              io_out_c_0_bypass_1_2_is_stationary,
  output     [15:0]   io_out_c_0_bypass_1_3_data,
  output              io_out_c_0_bypass_1_3_is_stationary,
  output              io_out_c_0_input_from_bypass_0,
  output              io_out_c_0_input_from_bypass_1,
  output     [15:0]   io_out_c_1_data_0_data,
  output              io_out_c_1_data_0_is_stationary,
  output     [15:0]   io_out_c_1_data_1_data,
  output              io_out_c_1_data_1_is_stationary,
  output     [15:0]   io_out_c_1_data_2_data,
  output              io_out_c_1_data_2_is_stationary,
  output     [15:0]   io_out_c_1_data_3_data,
  output              io_out_c_1_data_3_is_stationary,
  output     [15:0]   io_out_c_1_bypass_0_0_data,
  output              io_out_c_1_bypass_0_0_is_stationary,
  output     [15:0]   io_out_c_1_bypass_0_1_data,
  output              io_out_c_1_bypass_0_1_is_stationary,
  output     [15:0]   io_out_c_1_bypass_0_2_data,
  output              io_out_c_1_bypass_0_2_is_stationary,
  output     [15:0]   io_out_c_1_bypass_0_3_data,
  output              io_out_c_1_bypass_0_3_is_stationary,
  output     [15:0]   io_out_c_1_bypass_1_0_data,
  output              io_out_c_1_bypass_1_0_is_stationary,
  output     [15:0]   io_out_c_1_bypass_1_1_data,
  output              io_out_c_1_bypass_1_1_is_stationary,
  output     [15:0]   io_out_c_1_bypass_1_2_data,
  output              io_out_c_1_bypass_1_2_is_stationary,
  output     [15:0]   io_out_c_1_bypass_1_3_data,
  output              io_out_c_1_bypass_1_3_is_stationary,
  output              io_out_c_1_input_from_bypass_0,
  output              io_out_c_1_input_from_bypass_1,
  input               clk,
  input               reset
);

  wire       [15:0]   cellSARA_8_io_in_r_data_0_data;
  wire                cellSARA_8_io_in_r_data_0_load_store;
  wire                cellSARA_8_io_in_r_data_0_df_is_ws;
  wire                cellSARA_8_io_in_r_data_0_stall;
  wire       [15:0]   cellSARA_8_io_in_r_data_1_data;
  wire                cellSARA_8_io_in_r_data_1_load_store;
  wire                cellSARA_8_io_in_r_data_1_df_is_ws;
  wire                cellSARA_8_io_in_r_data_1_stall;
  wire       [15:0]   cellSARA_8_io_in_r_data_2_data;
  wire                cellSARA_8_io_in_r_data_2_load_store;
  wire                cellSARA_8_io_in_r_data_2_df_is_ws;
  wire                cellSARA_8_io_in_r_data_2_stall;
  wire       [15:0]   cellSARA_8_io_in_r_data_3_data;
  wire                cellSARA_8_io_in_r_data_3_load_store;
  wire                cellSARA_8_io_in_r_data_3_df_is_ws;
  wire                cellSARA_8_io_in_r_data_3_stall;
  wire       [15:0]   cellSARA_8_io_in_r_bypass_0_0_data;
  wire                cellSARA_8_io_in_r_bypass_0_0_load_store;
  wire                cellSARA_8_io_in_r_bypass_0_0_df_is_ws;
  wire                cellSARA_8_io_in_r_bypass_0_0_stall;
  wire       [15:0]   cellSARA_8_io_in_r_bypass_0_1_data;
  wire                cellSARA_8_io_in_r_bypass_0_1_load_store;
  wire                cellSARA_8_io_in_r_bypass_0_1_df_is_ws;
  wire                cellSARA_8_io_in_r_bypass_0_1_stall;
  wire       [15:0]   cellSARA_8_io_in_r_bypass_0_2_data;
  wire                cellSARA_8_io_in_r_bypass_0_2_load_store;
  wire                cellSARA_8_io_in_r_bypass_0_2_df_is_ws;
  wire                cellSARA_8_io_in_r_bypass_0_2_stall;
  wire       [15:0]   cellSARA_8_io_in_r_bypass_0_3_data;
  wire                cellSARA_8_io_in_r_bypass_0_3_load_store;
  wire                cellSARA_8_io_in_r_bypass_0_3_df_is_ws;
  wire                cellSARA_8_io_in_r_bypass_0_3_stall;
  wire       [15:0]   cellSARA_8_io_in_r_bypass_1_0_data;
  wire                cellSARA_8_io_in_r_bypass_1_0_load_store;
  wire                cellSARA_8_io_in_r_bypass_1_0_df_is_ws;
  wire                cellSARA_8_io_in_r_bypass_1_0_stall;
  wire       [15:0]   cellSARA_8_io_in_r_bypass_1_1_data;
  wire                cellSARA_8_io_in_r_bypass_1_1_load_store;
  wire                cellSARA_8_io_in_r_bypass_1_1_df_is_ws;
  wire                cellSARA_8_io_in_r_bypass_1_1_stall;
  wire       [15:0]   cellSARA_8_io_in_r_bypass_1_2_data;
  wire                cellSARA_8_io_in_r_bypass_1_2_load_store;
  wire                cellSARA_8_io_in_r_bypass_1_2_df_is_ws;
  wire                cellSARA_8_io_in_r_bypass_1_2_stall;
  wire       [15:0]   cellSARA_8_io_in_r_bypass_1_3_data;
  wire                cellSARA_8_io_in_r_bypass_1_3_load_store;
  wire                cellSARA_8_io_in_r_bypass_1_3_df_is_ws;
  wire                cellSARA_8_io_in_r_bypass_1_3_stall;
  wire                cellSARA_8_io_in_r_input_from_bypass_0;
  wire                cellSARA_8_io_in_r_input_from_bypass_1;
  wire       [15:0]   cellSARA_8_io_in_c_data_0_data;
  wire                cellSARA_8_io_in_c_data_0_is_stationary;
  wire       [15:0]   cellSARA_8_io_in_c_data_1_data;
  wire                cellSARA_8_io_in_c_data_1_is_stationary;
  wire       [15:0]   cellSARA_8_io_in_c_data_2_data;
  wire                cellSARA_8_io_in_c_data_2_is_stationary;
  wire       [15:0]   cellSARA_8_io_in_c_data_3_data;
  wire                cellSARA_8_io_in_c_data_3_is_stationary;
  wire       [15:0]   cellSARA_8_io_in_c_bypass_0_0_data;
  wire                cellSARA_8_io_in_c_bypass_0_0_is_stationary;
  wire       [15:0]   cellSARA_8_io_in_c_bypass_0_1_data;
  wire                cellSARA_8_io_in_c_bypass_0_1_is_stationary;
  wire       [15:0]   cellSARA_8_io_in_c_bypass_0_2_data;
  wire                cellSARA_8_io_in_c_bypass_0_2_is_stationary;
  wire       [15:0]   cellSARA_8_io_in_c_bypass_0_3_data;
  wire                cellSARA_8_io_in_c_bypass_0_3_is_stationary;
  wire       [15:0]   cellSARA_8_io_in_c_bypass_1_0_data;
  wire                cellSARA_8_io_in_c_bypass_1_0_is_stationary;
  wire       [15:0]   cellSARA_8_io_in_c_bypass_1_1_data;
  wire                cellSARA_8_io_in_c_bypass_1_1_is_stationary;
  wire       [15:0]   cellSARA_8_io_in_c_bypass_1_2_data;
  wire                cellSARA_8_io_in_c_bypass_1_2_is_stationary;
  wire       [15:0]   cellSARA_8_io_in_c_bypass_1_3_data;
  wire                cellSARA_8_io_in_c_bypass_1_3_is_stationary;
  wire                cellSARA_8_io_in_c_input_from_bypass_0;
  wire                cellSARA_8_io_in_c_input_from_bypass_1;
  wire       [15:0]   cellSARA_9_io_in_r_data_0_data;
  wire                cellSARA_9_io_in_r_data_0_load_store;
  wire                cellSARA_9_io_in_r_data_0_df_is_ws;
  wire                cellSARA_9_io_in_r_data_0_stall;
  wire       [15:0]   cellSARA_9_io_in_r_data_1_data;
  wire                cellSARA_9_io_in_r_data_1_load_store;
  wire                cellSARA_9_io_in_r_data_1_df_is_ws;
  wire                cellSARA_9_io_in_r_data_1_stall;
  wire       [15:0]   cellSARA_9_io_in_r_data_2_data;
  wire                cellSARA_9_io_in_r_data_2_load_store;
  wire                cellSARA_9_io_in_r_data_2_df_is_ws;
  wire                cellSARA_9_io_in_r_data_2_stall;
  wire       [15:0]   cellSARA_9_io_in_r_data_3_data;
  wire                cellSARA_9_io_in_r_data_3_load_store;
  wire                cellSARA_9_io_in_r_data_3_df_is_ws;
  wire                cellSARA_9_io_in_r_data_3_stall;
  wire       [15:0]   cellSARA_9_io_in_r_bypass_0_0_data;
  wire                cellSARA_9_io_in_r_bypass_0_0_load_store;
  wire                cellSARA_9_io_in_r_bypass_0_0_df_is_ws;
  wire                cellSARA_9_io_in_r_bypass_0_0_stall;
  wire       [15:0]   cellSARA_9_io_in_r_bypass_0_1_data;
  wire                cellSARA_9_io_in_r_bypass_0_1_load_store;
  wire                cellSARA_9_io_in_r_bypass_0_1_df_is_ws;
  wire                cellSARA_9_io_in_r_bypass_0_1_stall;
  wire       [15:0]   cellSARA_9_io_in_r_bypass_0_2_data;
  wire                cellSARA_9_io_in_r_bypass_0_2_load_store;
  wire                cellSARA_9_io_in_r_bypass_0_2_df_is_ws;
  wire                cellSARA_9_io_in_r_bypass_0_2_stall;
  wire       [15:0]   cellSARA_9_io_in_r_bypass_0_3_data;
  wire                cellSARA_9_io_in_r_bypass_0_3_load_store;
  wire                cellSARA_9_io_in_r_bypass_0_3_df_is_ws;
  wire                cellSARA_9_io_in_r_bypass_0_3_stall;
  wire       [15:0]   cellSARA_9_io_in_r_bypass_1_0_data;
  wire                cellSARA_9_io_in_r_bypass_1_0_load_store;
  wire                cellSARA_9_io_in_r_bypass_1_0_df_is_ws;
  wire                cellSARA_9_io_in_r_bypass_1_0_stall;
  wire       [15:0]   cellSARA_9_io_in_r_bypass_1_1_data;
  wire                cellSARA_9_io_in_r_bypass_1_1_load_store;
  wire                cellSARA_9_io_in_r_bypass_1_1_df_is_ws;
  wire                cellSARA_9_io_in_r_bypass_1_1_stall;
  wire       [15:0]   cellSARA_9_io_in_r_bypass_1_2_data;
  wire                cellSARA_9_io_in_r_bypass_1_2_load_store;
  wire                cellSARA_9_io_in_r_bypass_1_2_df_is_ws;
  wire                cellSARA_9_io_in_r_bypass_1_2_stall;
  wire       [15:0]   cellSARA_9_io_in_r_bypass_1_3_data;
  wire                cellSARA_9_io_in_r_bypass_1_3_load_store;
  wire                cellSARA_9_io_in_r_bypass_1_3_df_is_ws;
  wire                cellSARA_9_io_in_r_bypass_1_3_stall;
  wire                cellSARA_9_io_in_r_input_from_bypass_0;
  wire                cellSARA_9_io_in_r_input_from_bypass_1;
  wire       [15:0]   cellSARA_9_io_in_c_data_0_data;
  wire                cellSARA_9_io_in_c_data_0_is_stationary;
  wire       [15:0]   cellSARA_9_io_in_c_data_1_data;
  wire                cellSARA_9_io_in_c_data_1_is_stationary;
  wire       [15:0]   cellSARA_9_io_in_c_data_2_data;
  wire                cellSARA_9_io_in_c_data_2_is_stationary;
  wire       [15:0]   cellSARA_9_io_in_c_data_3_data;
  wire                cellSARA_9_io_in_c_data_3_is_stationary;
  wire       [15:0]   cellSARA_9_io_in_c_bypass_0_0_data;
  wire                cellSARA_9_io_in_c_bypass_0_0_is_stationary;
  wire       [15:0]   cellSARA_9_io_in_c_bypass_0_1_data;
  wire                cellSARA_9_io_in_c_bypass_0_1_is_stationary;
  wire       [15:0]   cellSARA_9_io_in_c_bypass_0_2_data;
  wire                cellSARA_9_io_in_c_bypass_0_2_is_stationary;
  wire       [15:0]   cellSARA_9_io_in_c_bypass_0_3_data;
  wire                cellSARA_9_io_in_c_bypass_0_3_is_stationary;
  wire       [15:0]   cellSARA_9_io_in_c_bypass_1_0_data;
  wire                cellSARA_9_io_in_c_bypass_1_0_is_stationary;
  wire       [15:0]   cellSARA_9_io_in_c_bypass_1_1_data;
  wire                cellSARA_9_io_in_c_bypass_1_1_is_stationary;
  wire       [15:0]   cellSARA_9_io_in_c_bypass_1_2_data;
  wire                cellSARA_9_io_in_c_bypass_1_2_is_stationary;
  wire       [15:0]   cellSARA_9_io_in_c_bypass_1_3_data;
  wire                cellSARA_9_io_in_c_bypass_1_3_is_stationary;
  wire                cellSARA_9_io_in_c_input_from_bypass_0;
  wire                cellSARA_9_io_in_c_input_from_bypass_1;
  wire       [15:0]   cellSARA_10_io_in_r_data_0_data;
  wire                cellSARA_10_io_in_r_data_0_load_store;
  wire                cellSARA_10_io_in_r_data_0_df_is_ws;
  wire                cellSARA_10_io_in_r_data_0_stall;
  wire       [15:0]   cellSARA_10_io_in_r_data_1_data;
  wire                cellSARA_10_io_in_r_data_1_load_store;
  wire                cellSARA_10_io_in_r_data_1_df_is_ws;
  wire                cellSARA_10_io_in_r_data_1_stall;
  wire       [15:0]   cellSARA_10_io_in_r_data_2_data;
  wire                cellSARA_10_io_in_r_data_2_load_store;
  wire                cellSARA_10_io_in_r_data_2_df_is_ws;
  wire                cellSARA_10_io_in_r_data_2_stall;
  wire       [15:0]   cellSARA_10_io_in_r_data_3_data;
  wire                cellSARA_10_io_in_r_data_3_load_store;
  wire                cellSARA_10_io_in_r_data_3_df_is_ws;
  wire                cellSARA_10_io_in_r_data_3_stall;
  wire       [15:0]   cellSARA_10_io_in_r_bypass_0_0_data;
  wire                cellSARA_10_io_in_r_bypass_0_0_load_store;
  wire                cellSARA_10_io_in_r_bypass_0_0_df_is_ws;
  wire                cellSARA_10_io_in_r_bypass_0_0_stall;
  wire       [15:0]   cellSARA_10_io_in_r_bypass_0_1_data;
  wire                cellSARA_10_io_in_r_bypass_0_1_load_store;
  wire                cellSARA_10_io_in_r_bypass_0_1_df_is_ws;
  wire                cellSARA_10_io_in_r_bypass_0_1_stall;
  wire       [15:0]   cellSARA_10_io_in_r_bypass_0_2_data;
  wire                cellSARA_10_io_in_r_bypass_0_2_load_store;
  wire                cellSARA_10_io_in_r_bypass_0_2_df_is_ws;
  wire                cellSARA_10_io_in_r_bypass_0_2_stall;
  wire       [15:0]   cellSARA_10_io_in_r_bypass_0_3_data;
  wire                cellSARA_10_io_in_r_bypass_0_3_load_store;
  wire                cellSARA_10_io_in_r_bypass_0_3_df_is_ws;
  wire                cellSARA_10_io_in_r_bypass_0_3_stall;
  wire       [15:0]   cellSARA_10_io_in_r_bypass_1_0_data;
  wire                cellSARA_10_io_in_r_bypass_1_0_load_store;
  wire                cellSARA_10_io_in_r_bypass_1_0_df_is_ws;
  wire                cellSARA_10_io_in_r_bypass_1_0_stall;
  wire       [15:0]   cellSARA_10_io_in_r_bypass_1_1_data;
  wire                cellSARA_10_io_in_r_bypass_1_1_load_store;
  wire                cellSARA_10_io_in_r_bypass_1_1_df_is_ws;
  wire                cellSARA_10_io_in_r_bypass_1_1_stall;
  wire       [15:0]   cellSARA_10_io_in_r_bypass_1_2_data;
  wire                cellSARA_10_io_in_r_bypass_1_2_load_store;
  wire                cellSARA_10_io_in_r_bypass_1_2_df_is_ws;
  wire                cellSARA_10_io_in_r_bypass_1_2_stall;
  wire       [15:0]   cellSARA_10_io_in_r_bypass_1_3_data;
  wire                cellSARA_10_io_in_r_bypass_1_3_load_store;
  wire                cellSARA_10_io_in_r_bypass_1_3_df_is_ws;
  wire                cellSARA_10_io_in_r_bypass_1_3_stall;
  wire                cellSARA_10_io_in_r_input_from_bypass_0;
  wire                cellSARA_10_io_in_r_input_from_bypass_1;
  wire       [15:0]   cellSARA_10_io_in_c_data_0_data;
  wire                cellSARA_10_io_in_c_data_0_is_stationary;
  wire       [15:0]   cellSARA_10_io_in_c_data_1_data;
  wire                cellSARA_10_io_in_c_data_1_is_stationary;
  wire       [15:0]   cellSARA_10_io_in_c_data_2_data;
  wire                cellSARA_10_io_in_c_data_2_is_stationary;
  wire       [15:0]   cellSARA_10_io_in_c_data_3_data;
  wire                cellSARA_10_io_in_c_data_3_is_stationary;
  wire       [15:0]   cellSARA_10_io_in_c_bypass_0_0_data;
  wire                cellSARA_10_io_in_c_bypass_0_0_is_stationary;
  wire       [15:0]   cellSARA_10_io_in_c_bypass_0_1_data;
  wire                cellSARA_10_io_in_c_bypass_0_1_is_stationary;
  wire       [15:0]   cellSARA_10_io_in_c_bypass_0_2_data;
  wire                cellSARA_10_io_in_c_bypass_0_2_is_stationary;
  wire       [15:0]   cellSARA_10_io_in_c_bypass_0_3_data;
  wire                cellSARA_10_io_in_c_bypass_0_3_is_stationary;
  wire       [15:0]   cellSARA_10_io_in_c_bypass_1_0_data;
  wire                cellSARA_10_io_in_c_bypass_1_0_is_stationary;
  wire       [15:0]   cellSARA_10_io_in_c_bypass_1_1_data;
  wire                cellSARA_10_io_in_c_bypass_1_1_is_stationary;
  wire       [15:0]   cellSARA_10_io_in_c_bypass_1_2_data;
  wire                cellSARA_10_io_in_c_bypass_1_2_is_stationary;
  wire       [15:0]   cellSARA_10_io_in_c_bypass_1_3_data;
  wire                cellSARA_10_io_in_c_bypass_1_3_is_stationary;
  wire                cellSARA_10_io_in_c_input_from_bypass_0;
  wire                cellSARA_10_io_in_c_input_from_bypass_1;
  wire       [15:0]   cellSARA_11_io_in_r_data_0_data;
  wire                cellSARA_11_io_in_r_data_0_load_store;
  wire                cellSARA_11_io_in_r_data_0_df_is_ws;
  wire                cellSARA_11_io_in_r_data_0_stall;
  wire       [15:0]   cellSARA_11_io_in_r_data_1_data;
  wire                cellSARA_11_io_in_r_data_1_load_store;
  wire                cellSARA_11_io_in_r_data_1_df_is_ws;
  wire                cellSARA_11_io_in_r_data_1_stall;
  wire       [15:0]   cellSARA_11_io_in_r_data_2_data;
  wire                cellSARA_11_io_in_r_data_2_load_store;
  wire                cellSARA_11_io_in_r_data_2_df_is_ws;
  wire                cellSARA_11_io_in_r_data_2_stall;
  wire       [15:0]   cellSARA_11_io_in_r_data_3_data;
  wire                cellSARA_11_io_in_r_data_3_load_store;
  wire                cellSARA_11_io_in_r_data_3_df_is_ws;
  wire                cellSARA_11_io_in_r_data_3_stall;
  wire       [15:0]   cellSARA_11_io_in_r_bypass_0_0_data;
  wire                cellSARA_11_io_in_r_bypass_0_0_load_store;
  wire                cellSARA_11_io_in_r_bypass_0_0_df_is_ws;
  wire                cellSARA_11_io_in_r_bypass_0_0_stall;
  wire       [15:0]   cellSARA_11_io_in_r_bypass_0_1_data;
  wire                cellSARA_11_io_in_r_bypass_0_1_load_store;
  wire                cellSARA_11_io_in_r_bypass_0_1_df_is_ws;
  wire                cellSARA_11_io_in_r_bypass_0_1_stall;
  wire       [15:0]   cellSARA_11_io_in_r_bypass_0_2_data;
  wire                cellSARA_11_io_in_r_bypass_0_2_load_store;
  wire                cellSARA_11_io_in_r_bypass_0_2_df_is_ws;
  wire                cellSARA_11_io_in_r_bypass_0_2_stall;
  wire       [15:0]   cellSARA_11_io_in_r_bypass_0_3_data;
  wire                cellSARA_11_io_in_r_bypass_0_3_load_store;
  wire                cellSARA_11_io_in_r_bypass_0_3_df_is_ws;
  wire                cellSARA_11_io_in_r_bypass_0_3_stall;
  wire       [15:0]   cellSARA_11_io_in_r_bypass_1_0_data;
  wire                cellSARA_11_io_in_r_bypass_1_0_load_store;
  wire                cellSARA_11_io_in_r_bypass_1_0_df_is_ws;
  wire                cellSARA_11_io_in_r_bypass_1_0_stall;
  wire       [15:0]   cellSARA_11_io_in_r_bypass_1_1_data;
  wire                cellSARA_11_io_in_r_bypass_1_1_load_store;
  wire                cellSARA_11_io_in_r_bypass_1_1_df_is_ws;
  wire                cellSARA_11_io_in_r_bypass_1_1_stall;
  wire       [15:0]   cellSARA_11_io_in_r_bypass_1_2_data;
  wire                cellSARA_11_io_in_r_bypass_1_2_load_store;
  wire                cellSARA_11_io_in_r_bypass_1_2_df_is_ws;
  wire                cellSARA_11_io_in_r_bypass_1_2_stall;
  wire       [15:0]   cellSARA_11_io_in_r_bypass_1_3_data;
  wire                cellSARA_11_io_in_r_bypass_1_3_load_store;
  wire                cellSARA_11_io_in_r_bypass_1_3_df_is_ws;
  wire                cellSARA_11_io_in_r_bypass_1_3_stall;
  wire                cellSARA_11_io_in_r_input_from_bypass_0;
  wire                cellSARA_11_io_in_r_input_from_bypass_1;
  wire       [15:0]   cellSARA_11_io_in_c_data_0_data;
  wire                cellSARA_11_io_in_c_data_0_is_stationary;
  wire       [15:0]   cellSARA_11_io_in_c_data_1_data;
  wire                cellSARA_11_io_in_c_data_1_is_stationary;
  wire       [15:0]   cellSARA_11_io_in_c_data_2_data;
  wire                cellSARA_11_io_in_c_data_2_is_stationary;
  wire       [15:0]   cellSARA_11_io_in_c_data_3_data;
  wire                cellSARA_11_io_in_c_data_3_is_stationary;
  wire       [15:0]   cellSARA_11_io_in_c_bypass_0_0_data;
  wire                cellSARA_11_io_in_c_bypass_0_0_is_stationary;
  wire       [15:0]   cellSARA_11_io_in_c_bypass_0_1_data;
  wire                cellSARA_11_io_in_c_bypass_0_1_is_stationary;
  wire       [15:0]   cellSARA_11_io_in_c_bypass_0_2_data;
  wire                cellSARA_11_io_in_c_bypass_0_2_is_stationary;
  wire       [15:0]   cellSARA_11_io_in_c_bypass_0_3_data;
  wire                cellSARA_11_io_in_c_bypass_0_3_is_stationary;
  wire       [15:0]   cellSARA_11_io_in_c_bypass_1_0_data;
  wire                cellSARA_11_io_in_c_bypass_1_0_is_stationary;
  wire       [15:0]   cellSARA_11_io_in_c_bypass_1_1_data;
  wire                cellSARA_11_io_in_c_bypass_1_1_is_stationary;
  wire       [15:0]   cellSARA_11_io_in_c_bypass_1_2_data;
  wire                cellSARA_11_io_in_c_bypass_1_2_is_stationary;
  wire       [15:0]   cellSARA_11_io_in_c_bypass_1_3_data;
  wire                cellSARA_11_io_in_c_bypass_1_3_is_stationary;
  wire                cellSARA_11_io_in_c_input_from_bypass_0;
  wire                cellSARA_11_io_in_c_input_from_bypass_1;
  wire       [15:0]   pes_0_0_io_out_r_data_0_data;
  wire                pes_0_0_io_out_r_data_0_load_store;
  wire                pes_0_0_io_out_r_data_0_df_is_ws;
  wire                pes_0_0_io_out_r_data_0_stall;
  wire       [15:0]   pes_0_0_io_out_r_data_1_data;
  wire                pes_0_0_io_out_r_data_1_load_store;
  wire                pes_0_0_io_out_r_data_1_df_is_ws;
  wire                pes_0_0_io_out_r_data_1_stall;
  wire       [15:0]   pes_0_0_io_out_r_data_2_data;
  wire                pes_0_0_io_out_r_data_2_load_store;
  wire                pes_0_0_io_out_r_data_2_df_is_ws;
  wire                pes_0_0_io_out_r_data_2_stall;
  wire       [15:0]   pes_0_0_io_out_r_data_3_data;
  wire                pes_0_0_io_out_r_data_3_load_store;
  wire                pes_0_0_io_out_r_data_3_df_is_ws;
  wire                pes_0_0_io_out_r_data_3_stall;
  wire       [15:0]   pes_0_0_io_out_r_bypass_0_0_data;
  wire                pes_0_0_io_out_r_bypass_0_0_load_store;
  wire                pes_0_0_io_out_r_bypass_0_0_df_is_ws;
  wire                pes_0_0_io_out_r_bypass_0_0_stall;
  wire       [15:0]   pes_0_0_io_out_r_bypass_0_1_data;
  wire                pes_0_0_io_out_r_bypass_0_1_load_store;
  wire                pes_0_0_io_out_r_bypass_0_1_df_is_ws;
  wire                pes_0_0_io_out_r_bypass_0_1_stall;
  wire       [15:0]   pes_0_0_io_out_r_bypass_0_2_data;
  wire                pes_0_0_io_out_r_bypass_0_2_load_store;
  wire                pes_0_0_io_out_r_bypass_0_2_df_is_ws;
  wire                pes_0_0_io_out_r_bypass_0_2_stall;
  wire       [15:0]   pes_0_0_io_out_r_bypass_0_3_data;
  wire                pes_0_0_io_out_r_bypass_0_3_load_store;
  wire                pes_0_0_io_out_r_bypass_0_3_df_is_ws;
  wire                pes_0_0_io_out_r_bypass_0_3_stall;
  wire       [15:0]   pes_0_0_io_out_r_bypass_1_0_data;
  wire                pes_0_0_io_out_r_bypass_1_0_load_store;
  wire                pes_0_0_io_out_r_bypass_1_0_df_is_ws;
  wire                pes_0_0_io_out_r_bypass_1_0_stall;
  wire       [15:0]   pes_0_0_io_out_r_bypass_1_1_data;
  wire                pes_0_0_io_out_r_bypass_1_1_load_store;
  wire                pes_0_0_io_out_r_bypass_1_1_df_is_ws;
  wire                pes_0_0_io_out_r_bypass_1_1_stall;
  wire       [15:0]   pes_0_0_io_out_r_bypass_1_2_data;
  wire                pes_0_0_io_out_r_bypass_1_2_load_store;
  wire                pes_0_0_io_out_r_bypass_1_2_df_is_ws;
  wire                pes_0_0_io_out_r_bypass_1_2_stall;
  wire       [15:0]   pes_0_0_io_out_r_bypass_1_3_data;
  wire                pes_0_0_io_out_r_bypass_1_3_load_store;
  wire                pes_0_0_io_out_r_bypass_1_3_df_is_ws;
  wire                pes_0_0_io_out_r_bypass_1_3_stall;
  wire                pes_0_0_io_out_r_input_from_bypass_0;
  wire                pes_0_0_io_out_r_input_from_bypass_1;
  wire       [15:0]   pes_0_0_io_out_c_data_0_data;
  wire                pes_0_0_io_out_c_data_0_is_stationary;
  wire       [15:0]   pes_0_0_io_out_c_data_1_data;
  wire                pes_0_0_io_out_c_data_1_is_stationary;
  wire       [15:0]   pes_0_0_io_out_c_data_2_data;
  wire                pes_0_0_io_out_c_data_2_is_stationary;
  wire       [15:0]   pes_0_0_io_out_c_data_3_data;
  wire                pes_0_0_io_out_c_data_3_is_stationary;
  wire       [15:0]   pes_0_0_io_out_c_bypass_0_0_data;
  wire                pes_0_0_io_out_c_bypass_0_0_is_stationary;
  wire       [15:0]   pes_0_0_io_out_c_bypass_0_1_data;
  wire                pes_0_0_io_out_c_bypass_0_1_is_stationary;
  wire       [15:0]   pes_0_0_io_out_c_bypass_0_2_data;
  wire                pes_0_0_io_out_c_bypass_0_2_is_stationary;
  wire       [15:0]   pes_0_0_io_out_c_bypass_0_3_data;
  wire                pes_0_0_io_out_c_bypass_0_3_is_stationary;
  wire       [15:0]   pes_0_0_io_out_c_bypass_1_0_data;
  wire                pes_0_0_io_out_c_bypass_1_0_is_stationary;
  wire       [15:0]   pes_0_0_io_out_c_bypass_1_1_data;
  wire                pes_0_0_io_out_c_bypass_1_1_is_stationary;
  wire       [15:0]   pes_0_0_io_out_c_bypass_1_2_data;
  wire                pes_0_0_io_out_c_bypass_1_2_is_stationary;
  wire       [15:0]   pes_0_0_io_out_c_bypass_1_3_data;
  wire                pes_0_0_io_out_c_bypass_1_3_is_stationary;
  wire                pes_0_0_io_out_c_input_from_bypass_0;
  wire                pes_0_0_io_out_c_input_from_bypass_1;
  wire       [15:0]   pes_0_1_io_out_r_data_0_data;
  wire                pes_0_1_io_out_r_data_0_load_store;
  wire                pes_0_1_io_out_r_data_0_df_is_ws;
  wire                pes_0_1_io_out_r_data_0_stall;
  wire       [15:0]   pes_0_1_io_out_r_data_1_data;
  wire                pes_0_1_io_out_r_data_1_load_store;
  wire                pes_0_1_io_out_r_data_1_df_is_ws;
  wire                pes_0_1_io_out_r_data_1_stall;
  wire       [15:0]   pes_0_1_io_out_r_data_2_data;
  wire                pes_0_1_io_out_r_data_2_load_store;
  wire                pes_0_1_io_out_r_data_2_df_is_ws;
  wire                pes_0_1_io_out_r_data_2_stall;
  wire       [15:0]   pes_0_1_io_out_r_data_3_data;
  wire                pes_0_1_io_out_r_data_3_load_store;
  wire                pes_0_1_io_out_r_data_3_df_is_ws;
  wire                pes_0_1_io_out_r_data_3_stall;
  wire       [15:0]   pes_0_1_io_out_r_bypass_0_0_data;
  wire                pes_0_1_io_out_r_bypass_0_0_load_store;
  wire                pes_0_1_io_out_r_bypass_0_0_df_is_ws;
  wire                pes_0_1_io_out_r_bypass_0_0_stall;
  wire       [15:0]   pes_0_1_io_out_r_bypass_0_1_data;
  wire                pes_0_1_io_out_r_bypass_0_1_load_store;
  wire                pes_0_1_io_out_r_bypass_0_1_df_is_ws;
  wire                pes_0_1_io_out_r_bypass_0_1_stall;
  wire       [15:0]   pes_0_1_io_out_r_bypass_0_2_data;
  wire                pes_0_1_io_out_r_bypass_0_2_load_store;
  wire                pes_0_1_io_out_r_bypass_0_2_df_is_ws;
  wire                pes_0_1_io_out_r_bypass_0_2_stall;
  wire       [15:0]   pes_0_1_io_out_r_bypass_0_3_data;
  wire                pes_0_1_io_out_r_bypass_0_3_load_store;
  wire                pes_0_1_io_out_r_bypass_0_3_df_is_ws;
  wire                pes_0_1_io_out_r_bypass_0_3_stall;
  wire       [15:0]   pes_0_1_io_out_r_bypass_1_0_data;
  wire                pes_0_1_io_out_r_bypass_1_0_load_store;
  wire                pes_0_1_io_out_r_bypass_1_0_df_is_ws;
  wire                pes_0_1_io_out_r_bypass_1_0_stall;
  wire       [15:0]   pes_0_1_io_out_r_bypass_1_1_data;
  wire                pes_0_1_io_out_r_bypass_1_1_load_store;
  wire                pes_0_1_io_out_r_bypass_1_1_df_is_ws;
  wire                pes_0_1_io_out_r_bypass_1_1_stall;
  wire       [15:0]   pes_0_1_io_out_r_bypass_1_2_data;
  wire                pes_0_1_io_out_r_bypass_1_2_load_store;
  wire                pes_0_1_io_out_r_bypass_1_2_df_is_ws;
  wire                pes_0_1_io_out_r_bypass_1_2_stall;
  wire       [15:0]   pes_0_1_io_out_r_bypass_1_3_data;
  wire                pes_0_1_io_out_r_bypass_1_3_load_store;
  wire                pes_0_1_io_out_r_bypass_1_3_df_is_ws;
  wire                pes_0_1_io_out_r_bypass_1_3_stall;
  wire                pes_0_1_io_out_r_input_from_bypass_0;
  wire                pes_0_1_io_out_r_input_from_bypass_1;
  wire       [15:0]   pes_0_1_io_out_c_data_0_data;
  wire                pes_0_1_io_out_c_data_0_is_stationary;
  wire       [15:0]   pes_0_1_io_out_c_data_1_data;
  wire                pes_0_1_io_out_c_data_1_is_stationary;
  wire       [15:0]   pes_0_1_io_out_c_data_2_data;
  wire                pes_0_1_io_out_c_data_2_is_stationary;
  wire       [15:0]   pes_0_1_io_out_c_data_3_data;
  wire                pes_0_1_io_out_c_data_3_is_stationary;
  wire       [15:0]   pes_0_1_io_out_c_bypass_0_0_data;
  wire                pes_0_1_io_out_c_bypass_0_0_is_stationary;
  wire       [15:0]   pes_0_1_io_out_c_bypass_0_1_data;
  wire                pes_0_1_io_out_c_bypass_0_1_is_stationary;
  wire       [15:0]   pes_0_1_io_out_c_bypass_0_2_data;
  wire                pes_0_1_io_out_c_bypass_0_2_is_stationary;
  wire       [15:0]   pes_0_1_io_out_c_bypass_0_3_data;
  wire                pes_0_1_io_out_c_bypass_0_3_is_stationary;
  wire       [15:0]   pes_0_1_io_out_c_bypass_1_0_data;
  wire                pes_0_1_io_out_c_bypass_1_0_is_stationary;
  wire       [15:0]   pes_0_1_io_out_c_bypass_1_1_data;
  wire                pes_0_1_io_out_c_bypass_1_1_is_stationary;
  wire       [15:0]   pes_0_1_io_out_c_bypass_1_2_data;
  wire                pes_0_1_io_out_c_bypass_1_2_is_stationary;
  wire       [15:0]   pes_0_1_io_out_c_bypass_1_3_data;
  wire                pes_0_1_io_out_c_bypass_1_3_is_stationary;
  wire                pes_0_1_io_out_c_input_from_bypass_0;
  wire                pes_0_1_io_out_c_input_from_bypass_1;
  wire       [15:0]   pes_1_0_io_out_r_data_0_data;
  wire                pes_1_0_io_out_r_data_0_load_store;
  wire                pes_1_0_io_out_r_data_0_df_is_ws;
  wire                pes_1_0_io_out_r_data_0_stall;
  wire       [15:0]   pes_1_0_io_out_r_data_1_data;
  wire                pes_1_0_io_out_r_data_1_load_store;
  wire                pes_1_0_io_out_r_data_1_df_is_ws;
  wire                pes_1_0_io_out_r_data_1_stall;
  wire       [15:0]   pes_1_0_io_out_r_data_2_data;
  wire                pes_1_0_io_out_r_data_2_load_store;
  wire                pes_1_0_io_out_r_data_2_df_is_ws;
  wire                pes_1_0_io_out_r_data_2_stall;
  wire       [15:0]   pes_1_0_io_out_r_data_3_data;
  wire                pes_1_0_io_out_r_data_3_load_store;
  wire                pes_1_0_io_out_r_data_3_df_is_ws;
  wire                pes_1_0_io_out_r_data_3_stall;
  wire       [15:0]   pes_1_0_io_out_r_bypass_0_0_data;
  wire                pes_1_0_io_out_r_bypass_0_0_load_store;
  wire                pes_1_0_io_out_r_bypass_0_0_df_is_ws;
  wire                pes_1_0_io_out_r_bypass_0_0_stall;
  wire       [15:0]   pes_1_0_io_out_r_bypass_0_1_data;
  wire                pes_1_0_io_out_r_bypass_0_1_load_store;
  wire                pes_1_0_io_out_r_bypass_0_1_df_is_ws;
  wire                pes_1_0_io_out_r_bypass_0_1_stall;
  wire       [15:0]   pes_1_0_io_out_r_bypass_0_2_data;
  wire                pes_1_0_io_out_r_bypass_0_2_load_store;
  wire                pes_1_0_io_out_r_bypass_0_2_df_is_ws;
  wire                pes_1_0_io_out_r_bypass_0_2_stall;
  wire       [15:0]   pes_1_0_io_out_r_bypass_0_3_data;
  wire                pes_1_0_io_out_r_bypass_0_3_load_store;
  wire                pes_1_0_io_out_r_bypass_0_3_df_is_ws;
  wire                pes_1_0_io_out_r_bypass_0_3_stall;
  wire       [15:0]   pes_1_0_io_out_r_bypass_1_0_data;
  wire                pes_1_0_io_out_r_bypass_1_0_load_store;
  wire                pes_1_0_io_out_r_bypass_1_0_df_is_ws;
  wire                pes_1_0_io_out_r_bypass_1_0_stall;
  wire       [15:0]   pes_1_0_io_out_r_bypass_1_1_data;
  wire                pes_1_0_io_out_r_bypass_1_1_load_store;
  wire                pes_1_0_io_out_r_bypass_1_1_df_is_ws;
  wire                pes_1_0_io_out_r_bypass_1_1_stall;
  wire       [15:0]   pes_1_0_io_out_r_bypass_1_2_data;
  wire                pes_1_0_io_out_r_bypass_1_2_load_store;
  wire                pes_1_0_io_out_r_bypass_1_2_df_is_ws;
  wire                pes_1_0_io_out_r_bypass_1_2_stall;
  wire       [15:0]   pes_1_0_io_out_r_bypass_1_3_data;
  wire                pes_1_0_io_out_r_bypass_1_3_load_store;
  wire                pes_1_0_io_out_r_bypass_1_3_df_is_ws;
  wire                pes_1_0_io_out_r_bypass_1_3_stall;
  wire                pes_1_0_io_out_r_input_from_bypass_0;
  wire                pes_1_0_io_out_r_input_from_bypass_1;
  wire       [15:0]   pes_1_0_io_out_c_data_0_data;
  wire                pes_1_0_io_out_c_data_0_is_stationary;
  wire       [15:0]   pes_1_0_io_out_c_data_1_data;
  wire                pes_1_0_io_out_c_data_1_is_stationary;
  wire       [15:0]   pes_1_0_io_out_c_data_2_data;
  wire                pes_1_0_io_out_c_data_2_is_stationary;
  wire       [15:0]   pes_1_0_io_out_c_data_3_data;
  wire                pes_1_0_io_out_c_data_3_is_stationary;
  wire       [15:0]   pes_1_0_io_out_c_bypass_0_0_data;
  wire                pes_1_0_io_out_c_bypass_0_0_is_stationary;
  wire       [15:0]   pes_1_0_io_out_c_bypass_0_1_data;
  wire                pes_1_0_io_out_c_bypass_0_1_is_stationary;
  wire       [15:0]   pes_1_0_io_out_c_bypass_0_2_data;
  wire                pes_1_0_io_out_c_bypass_0_2_is_stationary;
  wire       [15:0]   pes_1_0_io_out_c_bypass_0_3_data;
  wire                pes_1_0_io_out_c_bypass_0_3_is_stationary;
  wire       [15:0]   pes_1_0_io_out_c_bypass_1_0_data;
  wire                pes_1_0_io_out_c_bypass_1_0_is_stationary;
  wire       [15:0]   pes_1_0_io_out_c_bypass_1_1_data;
  wire                pes_1_0_io_out_c_bypass_1_1_is_stationary;
  wire       [15:0]   pes_1_0_io_out_c_bypass_1_2_data;
  wire                pes_1_0_io_out_c_bypass_1_2_is_stationary;
  wire       [15:0]   pes_1_0_io_out_c_bypass_1_3_data;
  wire                pes_1_0_io_out_c_bypass_1_3_is_stationary;
  wire                pes_1_0_io_out_c_input_from_bypass_0;
  wire                pes_1_0_io_out_c_input_from_bypass_1;
  wire       [15:0]   pes_1_1_io_out_r_data_0_data;
  wire                pes_1_1_io_out_r_data_0_load_store;
  wire                pes_1_1_io_out_r_data_0_df_is_ws;
  wire                pes_1_1_io_out_r_data_0_stall;
  wire       [15:0]   pes_1_1_io_out_r_data_1_data;
  wire                pes_1_1_io_out_r_data_1_load_store;
  wire                pes_1_1_io_out_r_data_1_df_is_ws;
  wire                pes_1_1_io_out_r_data_1_stall;
  wire       [15:0]   pes_1_1_io_out_r_data_2_data;
  wire                pes_1_1_io_out_r_data_2_load_store;
  wire                pes_1_1_io_out_r_data_2_df_is_ws;
  wire                pes_1_1_io_out_r_data_2_stall;
  wire       [15:0]   pes_1_1_io_out_r_data_3_data;
  wire                pes_1_1_io_out_r_data_3_load_store;
  wire                pes_1_1_io_out_r_data_3_df_is_ws;
  wire                pes_1_1_io_out_r_data_3_stall;
  wire       [15:0]   pes_1_1_io_out_r_bypass_0_0_data;
  wire                pes_1_1_io_out_r_bypass_0_0_load_store;
  wire                pes_1_1_io_out_r_bypass_0_0_df_is_ws;
  wire                pes_1_1_io_out_r_bypass_0_0_stall;
  wire       [15:0]   pes_1_1_io_out_r_bypass_0_1_data;
  wire                pes_1_1_io_out_r_bypass_0_1_load_store;
  wire                pes_1_1_io_out_r_bypass_0_1_df_is_ws;
  wire                pes_1_1_io_out_r_bypass_0_1_stall;
  wire       [15:0]   pes_1_1_io_out_r_bypass_0_2_data;
  wire                pes_1_1_io_out_r_bypass_0_2_load_store;
  wire                pes_1_1_io_out_r_bypass_0_2_df_is_ws;
  wire                pes_1_1_io_out_r_bypass_0_2_stall;
  wire       [15:0]   pes_1_1_io_out_r_bypass_0_3_data;
  wire                pes_1_1_io_out_r_bypass_0_3_load_store;
  wire                pes_1_1_io_out_r_bypass_0_3_df_is_ws;
  wire                pes_1_1_io_out_r_bypass_0_3_stall;
  wire       [15:0]   pes_1_1_io_out_r_bypass_1_0_data;
  wire                pes_1_1_io_out_r_bypass_1_0_load_store;
  wire                pes_1_1_io_out_r_bypass_1_0_df_is_ws;
  wire                pes_1_1_io_out_r_bypass_1_0_stall;
  wire       [15:0]   pes_1_1_io_out_r_bypass_1_1_data;
  wire                pes_1_1_io_out_r_bypass_1_1_load_store;
  wire                pes_1_1_io_out_r_bypass_1_1_df_is_ws;
  wire                pes_1_1_io_out_r_bypass_1_1_stall;
  wire       [15:0]   pes_1_1_io_out_r_bypass_1_2_data;
  wire                pes_1_1_io_out_r_bypass_1_2_load_store;
  wire                pes_1_1_io_out_r_bypass_1_2_df_is_ws;
  wire                pes_1_1_io_out_r_bypass_1_2_stall;
  wire       [15:0]   pes_1_1_io_out_r_bypass_1_3_data;
  wire                pes_1_1_io_out_r_bypass_1_3_load_store;
  wire                pes_1_1_io_out_r_bypass_1_3_df_is_ws;
  wire                pes_1_1_io_out_r_bypass_1_3_stall;
  wire                pes_1_1_io_out_r_input_from_bypass_0;
  wire                pes_1_1_io_out_r_input_from_bypass_1;
  wire       [15:0]   pes_1_1_io_out_c_data_0_data;
  wire                pes_1_1_io_out_c_data_0_is_stationary;
  wire       [15:0]   pes_1_1_io_out_c_data_1_data;
  wire                pes_1_1_io_out_c_data_1_is_stationary;
  wire       [15:0]   pes_1_1_io_out_c_data_2_data;
  wire                pes_1_1_io_out_c_data_2_is_stationary;
  wire       [15:0]   pes_1_1_io_out_c_data_3_data;
  wire                pes_1_1_io_out_c_data_3_is_stationary;
  wire       [15:0]   pes_1_1_io_out_c_bypass_0_0_data;
  wire                pes_1_1_io_out_c_bypass_0_0_is_stationary;
  wire       [15:0]   pes_1_1_io_out_c_bypass_0_1_data;
  wire                pes_1_1_io_out_c_bypass_0_1_is_stationary;
  wire       [15:0]   pes_1_1_io_out_c_bypass_0_2_data;
  wire                pes_1_1_io_out_c_bypass_0_2_is_stationary;
  wire       [15:0]   pes_1_1_io_out_c_bypass_0_3_data;
  wire                pes_1_1_io_out_c_bypass_0_3_is_stationary;
  wire       [15:0]   pes_1_1_io_out_c_bypass_1_0_data;
  wire                pes_1_1_io_out_c_bypass_1_0_is_stationary;
  wire       [15:0]   pes_1_1_io_out_c_bypass_1_1_data;
  wire                pes_1_1_io_out_c_bypass_1_1_is_stationary;
  wire       [15:0]   pes_1_1_io_out_c_bypass_1_2_data;
  wire                pes_1_1_io_out_c_bypass_1_2_is_stationary;
  wire       [15:0]   pes_1_1_io_out_c_bypass_1_3_data;
  wire                pes_1_1_io_out_c_bypass_1_3_is_stationary;
  wire                pes_1_1_io_out_c_input_from_bypass_0;
  wire                pes_1_1_io_out_c_input_from_bypass_1;
  wire       [15:0]   cellSARA_8_io_out_r_data_0_data;
  wire                cellSARA_8_io_out_r_data_0_load_store;
  wire                cellSARA_8_io_out_r_data_0_df_is_ws;
  wire                cellSARA_8_io_out_r_data_0_stall;
  wire       [15:0]   cellSARA_8_io_out_r_data_1_data;
  wire                cellSARA_8_io_out_r_data_1_load_store;
  wire                cellSARA_8_io_out_r_data_1_df_is_ws;
  wire                cellSARA_8_io_out_r_data_1_stall;
  wire       [15:0]   cellSARA_8_io_out_r_data_2_data;
  wire                cellSARA_8_io_out_r_data_2_load_store;
  wire                cellSARA_8_io_out_r_data_2_df_is_ws;
  wire                cellSARA_8_io_out_r_data_2_stall;
  wire       [15:0]   cellSARA_8_io_out_r_data_3_data;
  wire                cellSARA_8_io_out_r_data_3_load_store;
  wire                cellSARA_8_io_out_r_data_3_df_is_ws;
  wire                cellSARA_8_io_out_r_data_3_stall;
  wire       [15:0]   cellSARA_8_io_out_r_bypass_0_0_data;
  wire                cellSARA_8_io_out_r_bypass_0_0_load_store;
  wire                cellSARA_8_io_out_r_bypass_0_0_df_is_ws;
  wire                cellSARA_8_io_out_r_bypass_0_0_stall;
  wire       [15:0]   cellSARA_8_io_out_r_bypass_0_1_data;
  wire                cellSARA_8_io_out_r_bypass_0_1_load_store;
  wire                cellSARA_8_io_out_r_bypass_0_1_df_is_ws;
  wire                cellSARA_8_io_out_r_bypass_0_1_stall;
  wire       [15:0]   cellSARA_8_io_out_r_bypass_0_2_data;
  wire                cellSARA_8_io_out_r_bypass_0_2_load_store;
  wire                cellSARA_8_io_out_r_bypass_0_2_df_is_ws;
  wire                cellSARA_8_io_out_r_bypass_0_2_stall;
  wire       [15:0]   cellSARA_8_io_out_r_bypass_0_3_data;
  wire                cellSARA_8_io_out_r_bypass_0_3_load_store;
  wire                cellSARA_8_io_out_r_bypass_0_3_df_is_ws;
  wire                cellSARA_8_io_out_r_bypass_0_3_stall;
  wire       [15:0]   cellSARA_8_io_out_r_bypass_1_0_data;
  wire                cellSARA_8_io_out_r_bypass_1_0_load_store;
  wire                cellSARA_8_io_out_r_bypass_1_0_df_is_ws;
  wire                cellSARA_8_io_out_r_bypass_1_0_stall;
  wire       [15:0]   cellSARA_8_io_out_r_bypass_1_1_data;
  wire                cellSARA_8_io_out_r_bypass_1_1_load_store;
  wire                cellSARA_8_io_out_r_bypass_1_1_df_is_ws;
  wire                cellSARA_8_io_out_r_bypass_1_1_stall;
  wire       [15:0]   cellSARA_8_io_out_r_bypass_1_2_data;
  wire                cellSARA_8_io_out_r_bypass_1_2_load_store;
  wire                cellSARA_8_io_out_r_bypass_1_2_df_is_ws;
  wire                cellSARA_8_io_out_r_bypass_1_2_stall;
  wire       [15:0]   cellSARA_8_io_out_r_bypass_1_3_data;
  wire                cellSARA_8_io_out_r_bypass_1_3_load_store;
  wire                cellSARA_8_io_out_r_bypass_1_3_df_is_ws;
  wire                cellSARA_8_io_out_r_bypass_1_3_stall;
  wire                cellSARA_8_io_out_r_input_from_bypass_0;
  wire                cellSARA_8_io_out_r_input_from_bypass_1;
  wire       [15:0]   cellSARA_8_io_out_c_data_0_data;
  wire                cellSARA_8_io_out_c_data_0_is_stationary;
  wire       [15:0]   cellSARA_8_io_out_c_data_1_data;
  wire                cellSARA_8_io_out_c_data_1_is_stationary;
  wire       [15:0]   cellSARA_8_io_out_c_data_2_data;
  wire                cellSARA_8_io_out_c_data_2_is_stationary;
  wire       [15:0]   cellSARA_8_io_out_c_data_3_data;
  wire                cellSARA_8_io_out_c_data_3_is_stationary;
  wire       [15:0]   cellSARA_8_io_out_c_bypass_0_0_data;
  wire                cellSARA_8_io_out_c_bypass_0_0_is_stationary;
  wire       [15:0]   cellSARA_8_io_out_c_bypass_0_1_data;
  wire                cellSARA_8_io_out_c_bypass_0_1_is_stationary;
  wire       [15:0]   cellSARA_8_io_out_c_bypass_0_2_data;
  wire                cellSARA_8_io_out_c_bypass_0_2_is_stationary;
  wire       [15:0]   cellSARA_8_io_out_c_bypass_0_3_data;
  wire                cellSARA_8_io_out_c_bypass_0_3_is_stationary;
  wire       [15:0]   cellSARA_8_io_out_c_bypass_1_0_data;
  wire                cellSARA_8_io_out_c_bypass_1_0_is_stationary;
  wire       [15:0]   cellSARA_8_io_out_c_bypass_1_1_data;
  wire                cellSARA_8_io_out_c_bypass_1_1_is_stationary;
  wire       [15:0]   cellSARA_8_io_out_c_bypass_1_2_data;
  wire                cellSARA_8_io_out_c_bypass_1_2_is_stationary;
  wire       [15:0]   cellSARA_8_io_out_c_bypass_1_3_data;
  wire                cellSARA_8_io_out_c_bypass_1_3_is_stationary;
  wire                cellSARA_8_io_out_c_input_from_bypass_0;
  wire                cellSARA_8_io_out_c_input_from_bypass_1;
  wire       [15:0]   cellSARA_9_io_out_r_data_0_data;
  wire                cellSARA_9_io_out_r_data_0_load_store;
  wire                cellSARA_9_io_out_r_data_0_df_is_ws;
  wire                cellSARA_9_io_out_r_data_0_stall;
  wire       [15:0]   cellSARA_9_io_out_r_data_1_data;
  wire                cellSARA_9_io_out_r_data_1_load_store;
  wire                cellSARA_9_io_out_r_data_1_df_is_ws;
  wire                cellSARA_9_io_out_r_data_1_stall;
  wire       [15:0]   cellSARA_9_io_out_r_data_2_data;
  wire                cellSARA_9_io_out_r_data_2_load_store;
  wire                cellSARA_9_io_out_r_data_2_df_is_ws;
  wire                cellSARA_9_io_out_r_data_2_stall;
  wire       [15:0]   cellSARA_9_io_out_r_data_3_data;
  wire                cellSARA_9_io_out_r_data_3_load_store;
  wire                cellSARA_9_io_out_r_data_3_df_is_ws;
  wire                cellSARA_9_io_out_r_data_3_stall;
  wire       [15:0]   cellSARA_9_io_out_r_bypass_0_0_data;
  wire                cellSARA_9_io_out_r_bypass_0_0_load_store;
  wire                cellSARA_9_io_out_r_bypass_0_0_df_is_ws;
  wire                cellSARA_9_io_out_r_bypass_0_0_stall;
  wire       [15:0]   cellSARA_9_io_out_r_bypass_0_1_data;
  wire                cellSARA_9_io_out_r_bypass_0_1_load_store;
  wire                cellSARA_9_io_out_r_bypass_0_1_df_is_ws;
  wire                cellSARA_9_io_out_r_bypass_0_1_stall;
  wire       [15:0]   cellSARA_9_io_out_r_bypass_0_2_data;
  wire                cellSARA_9_io_out_r_bypass_0_2_load_store;
  wire                cellSARA_9_io_out_r_bypass_0_2_df_is_ws;
  wire                cellSARA_9_io_out_r_bypass_0_2_stall;
  wire       [15:0]   cellSARA_9_io_out_r_bypass_0_3_data;
  wire                cellSARA_9_io_out_r_bypass_0_3_load_store;
  wire                cellSARA_9_io_out_r_bypass_0_3_df_is_ws;
  wire                cellSARA_9_io_out_r_bypass_0_3_stall;
  wire       [15:0]   cellSARA_9_io_out_r_bypass_1_0_data;
  wire                cellSARA_9_io_out_r_bypass_1_0_load_store;
  wire                cellSARA_9_io_out_r_bypass_1_0_df_is_ws;
  wire                cellSARA_9_io_out_r_bypass_1_0_stall;
  wire       [15:0]   cellSARA_9_io_out_r_bypass_1_1_data;
  wire                cellSARA_9_io_out_r_bypass_1_1_load_store;
  wire                cellSARA_9_io_out_r_bypass_1_1_df_is_ws;
  wire                cellSARA_9_io_out_r_bypass_1_1_stall;
  wire       [15:0]   cellSARA_9_io_out_r_bypass_1_2_data;
  wire                cellSARA_9_io_out_r_bypass_1_2_load_store;
  wire                cellSARA_9_io_out_r_bypass_1_2_df_is_ws;
  wire                cellSARA_9_io_out_r_bypass_1_2_stall;
  wire       [15:0]   cellSARA_9_io_out_r_bypass_1_3_data;
  wire                cellSARA_9_io_out_r_bypass_1_3_load_store;
  wire                cellSARA_9_io_out_r_bypass_1_3_df_is_ws;
  wire                cellSARA_9_io_out_r_bypass_1_3_stall;
  wire                cellSARA_9_io_out_r_input_from_bypass_0;
  wire                cellSARA_9_io_out_r_input_from_bypass_1;
  wire       [15:0]   cellSARA_9_io_out_c_data_0_data;
  wire                cellSARA_9_io_out_c_data_0_is_stationary;
  wire       [15:0]   cellSARA_9_io_out_c_data_1_data;
  wire                cellSARA_9_io_out_c_data_1_is_stationary;
  wire       [15:0]   cellSARA_9_io_out_c_data_2_data;
  wire                cellSARA_9_io_out_c_data_2_is_stationary;
  wire       [15:0]   cellSARA_9_io_out_c_data_3_data;
  wire                cellSARA_9_io_out_c_data_3_is_stationary;
  wire       [15:0]   cellSARA_9_io_out_c_bypass_0_0_data;
  wire                cellSARA_9_io_out_c_bypass_0_0_is_stationary;
  wire       [15:0]   cellSARA_9_io_out_c_bypass_0_1_data;
  wire                cellSARA_9_io_out_c_bypass_0_1_is_stationary;
  wire       [15:0]   cellSARA_9_io_out_c_bypass_0_2_data;
  wire                cellSARA_9_io_out_c_bypass_0_2_is_stationary;
  wire       [15:0]   cellSARA_9_io_out_c_bypass_0_3_data;
  wire                cellSARA_9_io_out_c_bypass_0_3_is_stationary;
  wire       [15:0]   cellSARA_9_io_out_c_bypass_1_0_data;
  wire                cellSARA_9_io_out_c_bypass_1_0_is_stationary;
  wire       [15:0]   cellSARA_9_io_out_c_bypass_1_1_data;
  wire                cellSARA_9_io_out_c_bypass_1_1_is_stationary;
  wire       [15:0]   cellSARA_9_io_out_c_bypass_1_2_data;
  wire                cellSARA_9_io_out_c_bypass_1_2_is_stationary;
  wire       [15:0]   cellSARA_9_io_out_c_bypass_1_3_data;
  wire                cellSARA_9_io_out_c_bypass_1_3_is_stationary;
  wire                cellSARA_9_io_out_c_input_from_bypass_0;
  wire                cellSARA_9_io_out_c_input_from_bypass_1;
  wire       [15:0]   cellSARA_10_io_out_r_data_0_data;
  wire                cellSARA_10_io_out_r_data_0_load_store;
  wire                cellSARA_10_io_out_r_data_0_df_is_ws;
  wire                cellSARA_10_io_out_r_data_0_stall;
  wire       [15:0]   cellSARA_10_io_out_r_data_1_data;
  wire                cellSARA_10_io_out_r_data_1_load_store;
  wire                cellSARA_10_io_out_r_data_1_df_is_ws;
  wire                cellSARA_10_io_out_r_data_1_stall;
  wire       [15:0]   cellSARA_10_io_out_r_data_2_data;
  wire                cellSARA_10_io_out_r_data_2_load_store;
  wire                cellSARA_10_io_out_r_data_2_df_is_ws;
  wire                cellSARA_10_io_out_r_data_2_stall;
  wire       [15:0]   cellSARA_10_io_out_r_data_3_data;
  wire                cellSARA_10_io_out_r_data_3_load_store;
  wire                cellSARA_10_io_out_r_data_3_df_is_ws;
  wire                cellSARA_10_io_out_r_data_3_stall;
  wire       [15:0]   cellSARA_10_io_out_r_bypass_0_0_data;
  wire                cellSARA_10_io_out_r_bypass_0_0_load_store;
  wire                cellSARA_10_io_out_r_bypass_0_0_df_is_ws;
  wire                cellSARA_10_io_out_r_bypass_0_0_stall;
  wire       [15:0]   cellSARA_10_io_out_r_bypass_0_1_data;
  wire                cellSARA_10_io_out_r_bypass_0_1_load_store;
  wire                cellSARA_10_io_out_r_bypass_0_1_df_is_ws;
  wire                cellSARA_10_io_out_r_bypass_0_1_stall;
  wire       [15:0]   cellSARA_10_io_out_r_bypass_0_2_data;
  wire                cellSARA_10_io_out_r_bypass_0_2_load_store;
  wire                cellSARA_10_io_out_r_bypass_0_2_df_is_ws;
  wire                cellSARA_10_io_out_r_bypass_0_2_stall;
  wire       [15:0]   cellSARA_10_io_out_r_bypass_0_3_data;
  wire                cellSARA_10_io_out_r_bypass_0_3_load_store;
  wire                cellSARA_10_io_out_r_bypass_0_3_df_is_ws;
  wire                cellSARA_10_io_out_r_bypass_0_3_stall;
  wire       [15:0]   cellSARA_10_io_out_r_bypass_1_0_data;
  wire                cellSARA_10_io_out_r_bypass_1_0_load_store;
  wire                cellSARA_10_io_out_r_bypass_1_0_df_is_ws;
  wire                cellSARA_10_io_out_r_bypass_1_0_stall;
  wire       [15:0]   cellSARA_10_io_out_r_bypass_1_1_data;
  wire                cellSARA_10_io_out_r_bypass_1_1_load_store;
  wire                cellSARA_10_io_out_r_bypass_1_1_df_is_ws;
  wire                cellSARA_10_io_out_r_bypass_1_1_stall;
  wire       [15:0]   cellSARA_10_io_out_r_bypass_1_2_data;
  wire                cellSARA_10_io_out_r_bypass_1_2_load_store;
  wire                cellSARA_10_io_out_r_bypass_1_2_df_is_ws;
  wire                cellSARA_10_io_out_r_bypass_1_2_stall;
  wire       [15:0]   cellSARA_10_io_out_r_bypass_1_3_data;
  wire                cellSARA_10_io_out_r_bypass_1_3_load_store;
  wire                cellSARA_10_io_out_r_bypass_1_3_df_is_ws;
  wire                cellSARA_10_io_out_r_bypass_1_3_stall;
  wire                cellSARA_10_io_out_r_input_from_bypass_0;
  wire                cellSARA_10_io_out_r_input_from_bypass_1;
  wire       [15:0]   cellSARA_10_io_out_c_data_0_data;
  wire                cellSARA_10_io_out_c_data_0_is_stationary;
  wire       [15:0]   cellSARA_10_io_out_c_data_1_data;
  wire                cellSARA_10_io_out_c_data_1_is_stationary;
  wire       [15:0]   cellSARA_10_io_out_c_data_2_data;
  wire                cellSARA_10_io_out_c_data_2_is_stationary;
  wire       [15:0]   cellSARA_10_io_out_c_data_3_data;
  wire                cellSARA_10_io_out_c_data_3_is_stationary;
  wire       [15:0]   cellSARA_10_io_out_c_bypass_0_0_data;
  wire                cellSARA_10_io_out_c_bypass_0_0_is_stationary;
  wire       [15:0]   cellSARA_10_io_out_c_bypass_0_1_data;
  wire                cellSARA_10_io_out_c_bypass_0_1_is_stationary;
  wire       [15:0]   cellSARA_10_io_out_c_bypass_0_2_data;
  wire                cellSARA_10_io_out_c_bypass_0_2_is_stationary;
  wire       [15:0]   cellSARA_10_io_out_c_bypass_0_3_data;
  wire                cellSARA_10_io_out_c_bypass_0_3_is_stationary;
  wire       [15:0]   cellSARA_10_io_out_c_bypass_1_0_data;
  wire                cellSARA_10_io_out_c_bypass_1_0_is_stationary;
  wire       [15:0]   cellSARA_10_io_out_c_bypass_1_1_data;
  wire                cellSARA_10_io_out_c_bypass_1_1_is_stationary;
  wire       [15:0]   cellSARA_10_io_out_c_bypass_1_2_data;
  wire                cellSARA_10_io_out_c_bypass_1_2_is_stationary;
  wire       [15:0]   cellSARA_10_io_out_c_bypass_1_3_data;
  wire                cellSARA_10_io_out_c_bypass_1_3_is_stationary;
  wire                cellSARA_10_io_out_c_input_from_bypass_0;
  wire                cellSARA_10_io_out_c_input_from_bypass_1;
  wire       [15:0]   cellSARA_11_io_out_r_data_0_data;
  wire                cellSARA_11_io_out_r_data_0_load_store;
  wire                cellSARA_11_io_out_r_data_0_df_is_ws;
  wire                cellSARA_11_io_out_r_data_0_stall;
  wire       [15:0]   cellSARA_11_io_out_r_data_1_data;
  wire                cellSARA_11_io_out_r_data_1_load_store;
  wire                cellSARA_11_io_out_r_data_1_df_is_ws;
  wire                cellSARA_11_io_out_r_data_1_stall;
  wire       [15:0]   cellSARA_11_io_out_r_data_2_data;
  wire                cellSARA_11_io_out_r_data_2_load_store;
  wire                cellSARA_11_io_out_r_data_2_df_is_ws;
  wire                cellSARA_11_io_out_r_data_2_stall;
  wire       [15:0]   cellSARA_11_io_out_r_data_3_data;
  wire                cellSARA_11_io_out_r_data_3_load_store;
  wire                cellSARA_11_io_out_r_data_3_df_is_ws;
  wire                cellSARA_11_io_out_r_data_3_stall;
  wire       [15:0]   cellSARA_11_io_out_r_bypass_0_0_data;
  wire                cellSARA_11_io_out_r_bypass_0_0_load_store;
  wire                cellSARA_11_io_out_r_bypass_0_0_df_is_ws;
  wire                cellSARA_11_io_out_r_bypass_0_0_stall;
  wire       [15:0]   cellSARA_11_io_out_r_bypass_0_1_data;
  wire                cellSARA_11_io_out_r_bypass_0_1_load_store;
  wire                cellSARA_11_io_out_r_bypass_0_1_df_is_ws;
  wire                cellSARA_11_io_out_r_bypass_0_1_stall;
  wire       [15:0]   cellSARA_11_io_out_r_bypass_0_2_data;
  wire                cellSARA_11_io_out_r_bypass_0_2_load_store;
  wire                cellSARA_11_io_out_r_bypass_0_2_df_is_ws;
  wire                cellSARA_11_io_out_r_bypass_0_2_stall;
  wire       [15:0]   cellSARA_11_io_out_r_bypass_0_3_data;
  wire                cellSARA_11_io_out_r_bypass_0_3_load_store;
  wire                cellSARA_11_io_out_r_bypass_0_3_df_is_ws;
  wire                cellSARA_11_io_out_r_bypass_0_3_stall;
  wire       [15:0]   cellSARA_11_io_out_r_bypass_1_0_data;
  wire                cellSARA_11_io_out_r_bypass_1_0_load_store;
  wire                cellSARA_11_io_out_r_bypass_1_0_df_is_ws;
  wire                cellSARA_11_io_out_r_bypass_1_0_stall;
  wire       [15:0]   cellSARA_11_io_out_r_bypass_1_1_data;
  wire                cellSARA_11_io_out_r_bypass_1_1_load_store;
  wire                cellSARA_11_io_out_r_bypass_1_1_df_is_ws;
  wire                cellSARA_11_io_out_r_bypass_1_1_stall;
  wire       [15:0]   cellSARA_11_io_out_r_bypass_1_2_data;
  wire                cellSARA_11_io_out_r_bypass_1_2_load_store;
  wire                cellSARA_11_io_out_r_bypass_1_2_df_is_ws;
  wire                cellSARA_11_io_out_r_bypass_1_2_stall;
  wire       [15:0]   cellSARA_11_io_out_r_bypass_1_3_data;
  wire                cellSARA_11_io_out_r_bypass_1_3_load_store;
  wire                cellSARA_11_io_out_r_bypass_1_3_df_is_ws;
  wire                cellSARA_11_io_out_r_bypass_1_3_stall;
  wire                cellSARA_11_io_out_r_input_from_bypass_0;
  wire                cellSARA_11_io_out_r_input_from_bypass_1;
  wire       [15:0]   cellSARA_11_io_out_c_data_0_data;
  wire                cellSARA_11_io_out_c_data_0_is_stationary;
  wire       [15:0]   cellSARA_11_io_out_c_data_1_data;
  wire                cellSARA_11_io_out_c_data_1_is_stationary;
  wire       [15:0]   cellSARA_11_io_out_c_data_2_data;
  wire                cellSARA_11_io_out_c_data_2_is_stationary;
  wire       [15:0]   cellSARA_11_io_out_c_data_3_data;
  wire                cellSARA_11_io_out_c_data_3_is_stationary;
  wire       [15:0]   cellSARA_11_io_out_c_bypass_0_0_data;
  wire                cellSARA_11_io_out_c_bypass_0_0_is_stationary;
  wire       [15:0]   cellSARA_11_io_out_c_bypass_0_1_data;
  wire                cellSARA_11_io_out_c_bypass_0_1_is_stationary;
  wire       [15:0]   cellSARA_11_io_out_c_bypass_0_2_data;
  wire                cellSARA_11_io_out_c_bypass_0_2_is_stationary;
  wire       [15:0]   cellSARA_11_io_out_c_bypass_0_3_data;
  wire                cellSARA_11_io_out_c_bypass_0_3_is_stationary;
  wire       [15:0]   cellSARA_11_io_out_c_bypass_1_0_data;
  wire                cellSARA_11_io_out_c_bypass_1_0_is_stationary;
  wire       [15:0]   cellSARA_11_io_out_c_bypass_1_1_data;
  wire                cellSARA_11_io_out_c_bypass_1_1_is_stationary;
  wire       [15:0]   cellSARA_11_io_out_c_bypass_1_2_data;
  wire                cellSARA_11_io_out_c_bypass_1_2_is_stationary;
  wire       [15:0]   cellSARA_11_io_out_c_bypass_1_3_data;
  wire                cellSARA_11_io_out_c_bypass_1_3_is_stationary;
  wire                cellSARA_11_io_out_c_input_from_bypass_0;
  wire                cellSARA_11_io_out_c_input_from_bypass_1;

  CellSARA_7 pes_0_0 (
    .io_in_r_data_0_data               (io_in_r_0_data_0_data[15:0]              ), //i
    .io_in_r_data_0_load_store         (io_in_r_0_data_0_load_store              ), //i
    .io_in_r_data_0_df_is_ws           (io_in_r_0_data_0_df_is_ws                ), //i
    .io_in_r_data_0_stall              (io_in_r_0_data_0_stall                   ), //i
    .io_in_r_data_1_data               (io_in_r_0_data_1_data[15:0]              ), //i
    .io_in_r_data_1_load_store         (io_in_r_0_data_1_load_store              ), //i
    .io_in_r_data_1_df_is_ws           (io_in_r_0_data_1_df_is_ws                ), //i
    .io_in_r_data_1_stall              (io_in_r_0_data_1_stall                   ), //i
    .io_in_r_data_2_data               (io_in_r_0_data_2_data[15:0]              ), //i
    .io_in_r_data_2_load_store         (io_in_r_0_data_2_load_store              ), //i
    .io_in_r_data_2_df_is_ws           (io_in_r_0_data_2_df_is_ws                ), //i
    .io_in_r_data_2_stall              (io_in_r_0_data_2_stall                   ), //i
    .io_in_r_data_3_data               (io_in_r_0_data_3_data[15:0]              ), //i
    .io_in_r_data_3_load_store         (io_in_r_0_data_3_load_store              ), //i
    .io_in_r_data_3_df_is_ws           (io_in_r_0_data_3_df_is_ws                ), //i
    .io_in_r_data_3_stall              (io_in_r_0_data_3_stall                   ), //i
    .io_in_r_bypass_0_0_data           (io_in_r_0_bypass_0_0_data[15:0]          ), //i
    .io_in_r_bypass_0_0_load_store     (io_in_r_0_bypass_0_0_load_store          ), //i
    .io_in_r_bypass_0_0_df_is_ws       (io_in_r_0_bypass_0_0_df_is_ws            ), //i
    .io_in_r_bypass_0_0_stall          (io_in_r_0_bypass_0_0_stall               ), //i
    .io_in_r_bypass_0_1_data           (io_in_r_0_bypass_0_1_data[15:0]          ), //i
    .io_in_r_bypass_0_1_load_store     (io_in_r_0_bypass_0_1_load_store          ), //i
    .io_in_r_bypass_0_1_df_is_ws       (io_in_r_0_bypass_0_1_df_is_ws            ), //i
    .io_in_r_bypass_0_1_stall          (io_in_r_0_bypass_0_1_stall               ), //i
    .io_in_r_bypass_0_2_data           (io_in_r_0_bypass_0_2_data[15:0]          ), //i
    .io_in_r_bypass_0_2_load_store     (io_in_r_0_bypass_0_2_load_store          ), //i
    .io_in_r_bypass_0_2_df_is_ws       (io_in_r_0_bypass_0_2_df_is_ws            ), //i
    .io_in_r_bypass_0_2_stall          (io_in_r_0_bypass_0_2_stall               ), //i
    .io_in_r_bypass_0_3_data           (io_in_r_0_bypass_0_3_data[15:0]          ), //i
    .io_in_r_bypass_0_3_load_store     (io_in_r_0_bypass_0_3_load_store          ), //i
    .io_in_r_bypass_0_3_df_is_ws       (io_in_r_0_bypass_0_3_df_is_ws            ), //i
    .io_in_r_bypass_0_3_stall          (io_in_r_0_bypass_0_3_stall               ), //i
    .io_in_r_bypass_1_0_data           (io_in_r_0_bypass_1_0_data[15:0]          ), //i
    .io_in_r_bypass_1_0_load_store     (io_in_r_0_bypass_1_0_load_store          ), //i
    .io_in_r_bypass_1_0_df_is_ws       (io_in_r_0_bypass_1_0_df_is_ws            ), //i
    .io_in_r_bypass_1_0_stall          (io_in_r_0_bypass_1_0_stall               ), //i
    .io_in_r_bypass_1_1_data           (io_in_r_0_bypass_1_1_data[15:0]          ), //i
    .io_in_r_bypass_1_1_load_store     (io_in_r_0_bypass_1_1_load_store          ), //i
    .io_in_r_bypass_1_1_df_is_ws       (io_in_r_0_bypass_1_1_df_is_ws            ), //i
    .io_in_r_bypass_1_1_stall          (io_in_r_0_bypass_1_1_stall               ), //i
    .io_in_r_bypass_1_2_data           (io_in_r_0_bypass_1_2_data[15:0]          ), //i
    .io_in_r_bypass_1_2_load_store     (io_in_r_0_bypass_1_2_load_store          ), //i
    .io_in_r_bypass_1_2_df_is_ws       (io_in_r_0_bypass_1_2_df_is_ws            ), //i
    .io_in_r_bypass_1_2_stall          (io_in_r_0_bypass_1_2_stall               ), //i
    .io_in_r_bypass_1_3_data           (io_in_r_0_bypass_1_3_data[15:0]          ), //i
    .io_in_r_bypass_1_3_load_store     (io_in_r_0_bypass_1_3_load_store          ), //i
    .io_in_r_bypass_1_3_df_is_ws       (io_in_r_0_bypass_1_3_df_is_ws            ), //i
    .io_in_r_bypass_1_3_stall          (io_in_r_0_bypass_1_3_stall               ), //i
    .io_in_r_input_from_bypass_0       (io_in_r_0_input_from_bypass_0            ), //i
    .io_in_r_input_from_bypass_1       (io_in_r_0_input_from_bypass_1            ), //i
    .io_out_r_data_0_data              (pes_0_0_io_out_r_data_0_data[15:0]       ), //o
    .io_out_r_data_0_load_store        (pes_0_0_io_out_r_data_0_load_store       ), //o
    .io_out_r_data_0_df_is_ws          (pes_0_0_io_out_r_data_0_df_is_ws         ), //o
    .io_out_r_data_0_stall             (pes_0_0_io_out_r_data_0_stall            ), //o
    .io_out_r_data_1_data              (pes_0_0_io_out_r_data_1_data[15:0]       ), //o
    .io_out_r_data_1_load_store        (pes_0_0_io_out_r_data_1_load_store       ), //o
    .io_out_r_data_1_df_is_ws          (pes_0_0_io_out_r_data_1_df_is_ws         ), //o
    .io_out_r_data_1_stall             (pes_0_0_io_out_r_data_1_stall            ), //o
    .io_out_r_data_2_data              (pes_0_0_io_out_r_data_2_data[15:0]       ), //o
    .io_out_r_data_2_load_store        (pes_0_0_io_out_r_data_2_load_store       ), //o
    .io_out_r_data_2_df_is_ws          (pes_0_0_io_out_r_data_2_df_is_ws         ), //o
    .io_out_r_data_2_stall             (pes_0_0_io_out_r_data_2_stall            ), //o
    .io_out_r_data_3_data              (pes_0_0_io_out_r_data_3_data[15:0]       ), //o
    .io_out_r_data_3_load_store        (pes_0_0_io_out_r_data_3_load_store       ), //o
    .io_out_r_data_3_df_is_ws          (pes_0_0_io_out_r_data_3_df_is_ws         ), //o
    .io_out_r_data_3_stall             (pes_0_0_io_out_r_data_3_stall            ), //o
    .io_out_r_bypass_0_0_data          (pes_0_0_io_out_r_bypass_0_0_data[15:0]   ), //o
    .io_out_r_bypass_0_0_load_store    (pes_0_0_io_out_r_bypass_0_0_load_store   ), //o
    .io_out_r_bypass_0_0_df_is_ws      (pes_0_0_io_out_r_bypass_0_0_df_is_ws     ), //o
    .io_out_r_bypass_0_0_stall         (pes_0_0_io_out_r_bypass_0_0_stall        ), //o
    .io_out_r_bypass_0_1_data          (pes_0_0_io_out_r_bypass_0_1_data[15:0]   ), //o
    .io_out_r_bypass_0_1_load_store    (pes_0_0_io_out_r_bypass_0_1_load_store   ), //o
    .io_out_r_bypass_0_1_df_is_ws      (pes_0_0_io_out_r_bypass_0_1_df_is_ws     ), //o
    .io_out_r_bypass_0_1_stall         (pes_0_0_io_out_r_bypass_0_1_stall        ), //o
    .io_out_r_bypass_0_2_data          (pes_0_0_io_out_r_bypass_0_2_data[15:0]   ), //o
    .io_out_r_bypass_0_2_load_store    (pes_0_0_io_out_r_bypass_0_2_load_store   ), //o
    .io_out_r_bypass_0_2_df_is_ws      (pes_0_0_io_out_r_bypass_0_2_df_is_ws     ), //o
    .io_out_r_bypass_0_2_stall         (pes_0_0_io_out_r_bypass_0_2_stall        ), //o
    .io_out_r_bypass_0_3_data          (pes_0_0_io_out_r_bypass_0_3_data[15:0]   ), //o
    .io_out_r_bypass_0_3_load_store    (pes_0_0_io_out_r_bypass_0_3_load_store   ), //o
    .io_out_r_bypass_0_3_df_is_ws      (pes_0_0_io_out_r_bypass_0_3_df_is_ws     ), //o
    .io_out_r_bypass_0_3_stall         (pes_0_0_io_out_r_bypass_0_3_stall        ), //o
    .io_out_r_bypass_1_0_data          (pes_0_0_io_out_r_bypass_1_0_data[15:0]   ), //o
    .io_out_r_bypass_1_0_load_store    (pes_0_0_io_out_r_bypass_1_0_load_store   ), //o
    .io_out_r_bypass_1_0_df_is_ws      (pes_0_0_io_out_r_bypass_1_0_df_is_ws     ), //o
    .io_out_r_bypass_1_0_stall         (pes_0_0_io_out_r_bypass_1_0_stall        ), //o
    .io_out_r_bypass_1_1_data          (pes_0_0_io_out_r_bypass_1_1_data[15:0]   ), //o
    .io_out_r_bypass_1_1_load_store    (pes_0_0_io_out_r_bypass_1_1_load_store   ), //o
    .io_out_r_bypass_1_1_df_is_ws      (pes_0_0_io_out_r_bypass_1_1_df_is_ws     ), //o
    .io_out_r_bypass_1_1_stall         (pes_0_0_io_out_r_bypass_1_1_stall        ), //o
    .io_out_r_bypass_1_2_data          (pes_0_0_io_out_r_bypass_1_2_data[15:0]   ), //o
    .io_out_r_bypass_1_2_load_store    (pes_0_0_io_out_r_bypass_1_2_load_store   ), //o
    .io_out_r_bypass_1_2_df_is_ws      (pes_0_0_io_out_r_bypass_1_2_df_is_ws     ), //o
    .io_out_r_bypass_1_2_stall         (pes_0_0_io_out_r_bypass_1_2_stall        ), //o
    .io_out_r_bypass_1_3_data          (pes_0_0_io_out_r_bypass_1_3_data[15:0]   ), //o
    .io_out_r_bypass_1_3_load_store    (pes_0_0_io_out_r_bypass_1_3_load_store   ), //o
    .io_out_r_bypass_1_3_df_is_ws      (pes_0_0_io_out_r_bypass_1_3_df_is_ws     ), //o
    .io_out_r_bypass_1_3_stall         (pes_0_0_io_out_r_bypass_1_3_stall        ), //o
    .io_out_r_input_from_bypass_0      (pes_0_0_io_out_r_input_from_bypass_0     ), //o
    .io_out_r_input_from_bypass_1      (pes_0_0_io_out_r_input_from_bypass_1     ), //o
    .io_in_c_data_0_data               (io_in_c_0_data_0_data[15:0]              ), //i
    .io_in_c_data_0_is_stationary      (io_in_c_0_data_0_is_stationary           ), //i
    .io_in_c_data_1_data               (io_in_c_0_data_1_data[15:0]              ), //i
    .io_in_c_data_1_is_stationary      (io_in_c_0_data_1_is_stationary           ), //i
    .io_in_c_data_2_data               (io_in_c_0_data_2_data[15:0]              ), //i
    .io_in_c_data_2_is_stationary      (io_in_c_0_data_2_is_stationary           ), //i
    .io_in_c_data_3_data               (io_in_c_0_data_3_data[15:0]              ), //i
    .io_in_c_data_3_is_stationary      (io_in_c_0_data_3_is_stationary           ), //i
    .io_in_c_bypass_0_0_data           (io_in_c_0_bypass_0_0_data[15:0]          ), //i
    .io_in_c_bypass_0_0_is_stationary  (io_in_c_0_bypass_0_0_is_stationary       ), //i
    .io_in_c_bypass_0_1_data           (io_in_c_0_bypass_0_1_data[15:0]          ), //i
    .io_in_c_bypass_0_1_is_stationary  (io_in_c_0_bypass_0_1_is_stationary       ), //i
    .io_in_c_bypass_0_2_data           (io_in_c_0_bypass_0_2_data[15:0]          ), //i
    .io_in_c_bypass_0_2_is_stationary  (io_in_c_0_bypass_0_2_is_stationary       ), //i
    .io_in_c_bypass_0_3_data           (io_in_c_0_bypass_0_3_data[15:0]          ), //i
    .io_in_c_bypass_0_3_is_stationary  (io_in_c_0_bypass_0_3_is_stationary       ), //i
    .io_in_c_bypass_1_0_data           (io_in_c_0_bypass_1_0_data[15:0]          ), //i
    .io_in_c_bypass_1_0_is_stationary  (io_in_c_0_bypass_1_0_is_stationary       ), //i
    .io_in_c_bypass_1_1_data           (io_in_c_0_bypass_1_1_data[15:0]          ), //i
    .io_in_c_bypass_1_1_is_stationary  (io_in_c_0_bypass_1_1_is_stationary       ), //i
    .io_in_c_bypass_1_2_data           (io_in_c_0_bypass_1_2_data[15:0]          ), //i
    .io_in_c_bypass_1_2_is_stationary  (io_in_c_0_bypass_1_2_is_stationary       ), //i
    .io_in_c_bypass_1_3_data           (io_in_c_0_bypass_1_3_data[15:0]          ), //i
    .io_in_c_bypass_1_3_is_stationary  (io_in_c_0_bypass_1_3_is_stationary       ), //i
    .io_in_c_input_from_bypass_0       (io_in_c_0_input_from_bypass_0            ), //i
    .io_in_c_input_from_bypass_1       (io_in_c_0_input_from_bypass_1            ), //i
    .io_out_c_data_0_data              (pes_0_0_io_out_c_data_0_data[15:0]       ), //o
    .io_out_c_data_0_is_stationary     (pes_0_0_io_out_c_data_0_is_stationary    ), //o
    .io_out_c_data_1_data              (pes_0_0_io_out_c_data_1_data[15:0]       ), //o
    .io_out_c_data_1_is_stationary     (pes_0_0_io_out_c_data_1_is_stationary    ), //o
    .io_out_c_data_2_data              (pes_0_0_io_out_c_data_2_data[15:0]       ), //o
    .io_out_c_data_2_is_stationary     (pes_0_0_io_out_c_data_2_is_stationary    ), //o
    .io_out_c_data_3_data              (pes_0_0_io_out_c_data_3_data[15:0]       ), //o
    .io_out_c_data_3_is_stationary     (pes_0_0_io_out_c_data_3_is_stationary    ), //o
    .io_out_c_bypass_0_0_data          (pes_0_0_io_out_c_bypass_0_0_data[15:0]   ), //o
    .io_out_c_bypass_0_0_is_stationary (pes_0_0_io_out_c_bypass_0_0_is_stationary), //o
    .io_out_c_bypass_0_1_data          (pes_0_0_io_out_c_bypass_0_1_data[15:0]   ), //o
    .io_out_c_bypass_0_1_is_stationary (pes_0_0_io_out_c_bypass_0_1_is_stationary), //o
    .io_out_c_bypass_0_2_data          (pes_0_0_io_out_c_bypass_0_2_data[15:0]   ), //o
    .io_out_c_bypass_0_2_is_stationary (pes_0_0_io_out_c_bypass_0_2_is_stationary), //o
    .io_out_c_bypass_0_3_data          (pes_0_0_io_out_c_bypass_0_3_data[15:0]   ), //o
    .io_out_c_bypass_0_3_is_stationary (pes_0_0_io_out_c_bypass_0_3_is_stationary), //o
    .io_out_c_bypass_1_0_data          (pes_0_0_io_out_c_bypass_1_0_data[15:0]   ), //o
    .io_out_c_bypass_1_0_is_stationary (pes_0_0_io_out_c_bypass_1_0_is_stationary), //o
    .io_out_c_bypass_1_1_data          (pes_0_0_io_out_c_bypass_1_1_data[15:0]   ), //o
    .io_out_c_bypass_1_1_is_stationary (pes_0_0_io_out_c_bypass_1_1_is_stationary), //o
    .io_out_c_bypass_1_2_data          (pes_0_0_io_out_c_bypass_1_2_data[15:0]   ), //o
    .io_out_c_bypass_1_2_is_stationary (pes_0_0_io_out_c_bypass_1_2_is_stationary), //o
    .io_out_c_bypass_1_3_data          (pes_0_0_io_out_c_bypass_1_3_data[15:0]   ), //o
    .io_out_c_bypass_1_3_is_stationary (pes_0_0_io_out_c_bypass_1_3_is_stationary), //o
    .io_out_c_input_from_bypass_0      (pes_0_0_io_out_c_input_from_bypass_0     ), //o
    .io_out_c_input_from_bypass_1      (pes_0_0_io_out_c_input_from_bypass_1     ), //o
    .clk                               (clk                                      ), //i
    .reset                             (reset                                    )  //i
  );
  CellSARA_7 pes_0_1 (
    .io_in_r_data_0_data               (pes_0_0_io_out_r_data_0_data[15:0]       ), //i
    .io_in_r_data_0_load_store         (pes_0_0_io_out_r_data_0_load_store       ), //i
    .io_in_r_data_0_df_is_ws           (pes_0_0_io_out_r_data_0_df_is_ws         ), //i
    .io_in_r_data_0_stall              (pes_0_0_io_out_r_data_0_stall            ), //i
    .io_in_r_data_1_data               (pes_0_0_io_out_r_data_1_data[15:0]       ), //i
    .io_in_r_data_1_load_store         (pes_0_0_io_out_r_data_1_load_store       ), //i
    .io_in_r_data_1_df_is_ws           (pes_0_0_io_out_r_data_1_df_is_ws         ), //i
    .io_in_r_data_1_stall              (pes_0_0_io_out_r_data_1_stall            ), //i
    .io_in_r_data_2_data               (pes_0_0_io_out_r_data_2_data[15:0]       ), //i
    .io_in_r_data_2_load_store         (pes_0_0_io_out_r_data_2_load_store       ), //i
    .io_in_r_data_2_df_is_ws           (pes_0_0_io_out_r_data_2_df_is_ws         ), //i
    .io_in_r_data_2_stall              (pes_0_0_io_out_r_data_2_stall            ), //i
    .io_in_r_data_3_data               (pes_0_0_io_out_r_data_3_data[15:0]       ), //i
    .io_in_r_data_3_load_store         (pes_0_0_io_out_r_data_3_load_store       ), //i
    .io_in_r_data_3_df_is_ws           (pes_0_0_io_out_r_data_3_df_is_ws         ), //i
    .io_in_r_data_3_stall              (pes_0_0_io_out_r_data_3_stall            ), //i
    .io_in_r_bypass_0_0_data           (pes_0_0_io_out_r_bypass_0_0_data[15:0]   ), //i
    .io_in_r_bypass_0_0_load_store     (pes_0_0_io_out_r_bypass_0_0_load_store   ), //i
    .io_in_r_bypass_0_0_df_is_ws       (pes_0_0_io_out_r_bypass_0_0_df_is_ws     ), //i
    .io_in_r_bypass_0_0_stall          (pes_0_0_io_out_r_bypass_0_0_stall        ), //i
    .io_in_r_bypass_0_1_data           (pes_0_0_io_out_r_bypass_0_1_data[15:0]   ), //i
    .io_in_r_bypass_0_1_load_store     (pes_0_0_io_out_r_bypass_0_1_load_store   ), //i
    .io_in_r_bypass_0_1_df_is_ws       (pes_0_0_io_out_r_bypass_0_1_df_is_ws     ), //i
    .io_in_r_bypass_0_1_stall          (pes_0_0_io_out_r_bypass_0_1_stall        ), //i
    .io_in_r_bypass_0_2_data           (pes_0_0_io_out_r_bypass_0_2_data[15:0]   ), //i
    .io_in_r_bypass_0_2_load_store     (pes_0_0_io_out_r_bypass_0_2_load_store   ), //i
    .io_in_r_bypass_0_2_df_is_ws       (pes_0_0_io_out_r_bypass_0_2_df_is_ws     ), //i
    .io_in_r_bypass_0_2_stall          (pes_0_0_io_out_r_bypass_0_2_stall        ), //i
    .io_in_r_bypass_0_3_data           (pes_0_0_io_out_r_bypass_0_3_data[15:0]   ), //i
    .io_in_r_bypass_0_3_load_store     (pes_0_0_io_out_r_bypass_0_3_load_store   ), //i
    .io_in_r_bypass_0_3_df_is_ws       (pes_0_0_io_out_r_bypass_0_3_df_is_ws     ), //i
    .io_in_r_bypass_0_3_stall          (pes_0_0_io_out_r_bypass_0_3_stall        ), //i
    .io_in_r_bypass_1_0_data           (pes_0_0_io_out_r_bypass_1_0_data[15:0]   ), //i
    .io_in_r_bypass_1_0_load_store     (pes_0_0_io_out_r_bypass_1_0_load_store   ), //i
    .io_in_r_bypass_1_0_df_is_ws       (pes_0_0_io_out_r_bypass_1_0_df_is_ws     ), //i
    .io_in_r_bypass_1_0_stall          (pes_0_0_io_out_r_bypass_1_0_stall        ), //i
    .io_in_r_bypass_1_1_data           (pes_0_0_io_out_r_bypass_1_1_data[15:0]   ), //i
    .io_in_r_bypass_1_1_load_store     (pes_0_0_io_out_r_bypass_1_1_load_store   ), //i
    .io_in_r_bypass_1_1_df_is_ws       (pes_0_0_io_out_r_bypass_1_1_df_is_ws     ), //i
    .io_in_r_bypass_1_1_stall          (pes_0_0_io_out_r_bypass_1_1_stall        ), //i
    .io_in_r_bypass_1_2_data           (pes_0_0_io_out_r_bypass_1_2_data[15:0]   ), //i
    .io_in_r_bypass_1_2_load_store     (pes_0_0_io_out_r_bypass_1_2_load_store   ), //i
    .io_in_r_bypass_1_2_df_is_ws       (pes_0_0_io_out_r_bypass_1_2_df_is_ws     ), //i
    .io_in_r_bypass_1_2_stall          (pes_0_0_io_out_r_bypass_1_2_stall        ), //i
    .io_in_r_bypass_1_3_data           (pes_0_0_io_out_r_bypass_1_3_data[15:0]   ), //i
    .io_in_r_bypass_1_3_load_store     (pes_0_0_io_out_r_bypass_1_3_load_store   ), //i
    .io_in_r_bypass_1_3_df_is_ws       (pes_0_0_io_out_r_bypass_1_3_df_is_ws     ), //i
    .io_in_r_bypass_1_3_stall          (pes_0_0_io_out_r_bypass_1_3_stall        ), //i
    .io_in_r_input_from_bypass_0       (pes_0_0_io_out_r_input_from_bypass_0     ), //i
    .io_in_r_input_from_bypass_1       (pes_0_0_io_out_r_input_from_bypass_1     ), //i
    .io_out_r_data_0_data              (pes_0_1_io_out_r_data_0_data[15:0]       ), //o
    .io_out_r_data_0_load_store        (pes_0_1_io_out_r_data_0_load_store       ), //o
    .io_out_r_data_0_df_is_ws          (pes_0_1_io_out_r_data_0_df_is_ws         ), //o
    .io_out_r_data_0_stall             (pes_0_1_io_out_r_data_0_stall            ), //o
    .io_out_r_data_1_data              (pes_0_1_io_out_r_data_1_data[15:0]       ), //o
    .io_out_r_data_1_load_store        (pes_0_1_io_out_r_data_1_load_store       ), //o
    .io_out_r_data_1_df_is_ws          (pes_0_1_io_out_r_data_1_df_is_ws         ), //o
    .io_out_r_data_1_stall             (pes_0_1_io_out_r_data_1_stall            ), //o
    .io_out_r_data_2_data              (pes_0_1_io_out_r_data_2_data[15:0]       ), //o
    .io_out_r_data_2_load_store        (pes_0_1_io_out_r_data_2_load_store       ), //o
    .io_out_r_data_2_df_is_ws          (pes_0_1_io_out_r_data_2_df_is_ws         ), //o
    .io_out_r_data_2_stall             (pes_0_1_io_out_r_data_2_stall            ), //o
    .io_out_r_data_3_data              (pes_0_1_io_out_r_data_3_data[15:0]       ), //o
    .io_out_r_data_3_load_store        (pes_0_1_io_out_r_data_3_load_store       ), //o
    .io_out_r_data_3_df_is_ws          (pes_0_1_io_out_r_data_3_df_is_ws         ), //o
    .io_out_r_data_3_stall             (pes_0_1_io_out_r_data_3_stall            ), //o
    .io_out_r_bypass_0_0_data          (pes_0_1_io_out_r_bypass_0_0_data[15:0]   ), //o
    .io_out_r_bypass_0_0_load_store    (pes_0_1_io_out_r_bypass_0_0_load_store   ), //o
    .io_out_r_bypass_0_0_df_is_ws      (pes_0_1_io_out_r_bypass_0_0_df_is_ws     ), //o
    .io_out_r_bypass_0_0_stall         (pes_0_1_io_out_r_bypass_0_0_stall        ), //o
    .io_out_r_bypass_0_1_data          (pes_0_1_io_out_r_bypass_0_1_data[15:0]   ), //o
    .io_out_r_bypass_0_1_load_store    (pes_0_1_io_out_r_bypass_0_1_load_store   ), //o
    .io_out_r_bypass_0_1_df_is_ws      (pes_0_1_io_out_r_bypass_0_1_df_is_ws     ), //o
    .io_out_r_bypass_0_1_stall         (pes_0_1_io_out_r_bypass_0_1_stall        ), //o
    .io_out_r_bypass_0_2_data          (pes_0_1_io_out_r_bypass_0_2_data[15:0]   ), //o
    .io_out_r_bypass_0_2_load_store    (pes_0_1_io_out_r_bypass_0_2_load_store   ), //o
    .io_out_r_bypass_0_2_df_is_ws      (pes_0_1_io_out_r_bypass_0_2_df_is_ws     ), //o
    .io_out_r_bypass_0_2_stall         (pes_0_1_io_out_r_bypass_0_2_stall        ), //o
    .io_out_r_bypass_0_3_data          (pes_0_1_io_out_r_bypass_0_3_data[15:0]   ), //o
    .io_out_r_bypass_0_3_load_store    (pes_0_1_io_out_r_bypass_0_3_load_store   ), //o
    .io_out_r_bypass_0_3_df_is_ws      (pes_0_1_io_out_r_bypass_0_3_df_is_ws     ), //o
    .io_out_r_bypass_0_3_stall         (pes_0_1_io_out_r_bypass_0_3_stall        ), //o
    .io_out_r_bypass_1_0_data          (pes_0_1_io_out_r_bypass_1_0_data[15:0]   ), //o
    .io_out_r_bypass_1_0_load_store    (pes_0_1_io_out_r_bypass_1_0_load_store   ), //o
    .io_out_r_bypass_1_0_df_is_ws      (pes_0_1_io_out_r_bypass_1_0_df_is_ws     ), //o
    .io_out_r_bypass_1_0_stall         (pes_0_1_io_out_r_bypass_1_0_stall        ), //o
    .io_out_r_bypass_1_1_data          (pes_0_1_io_out_r_bypass_1_1_data[15:0]   ), //o
    .io_out_r_bypass_1_1_load_store    (pes_0_1_io_out_r_bypass_1_1_load_store   ), //o
    .io_out_r_bypass_1_1_df_is_ws      (pes_0_1_io_out_r_bypass_1_1_df_is_ws     ), //o
    .io_out_r_bypass_1_1_stall         (pes_0_1_io_out_r_bypass_1_1_stall        ), //o
    .io_out_r_bypass_1_2_data          (pes_0_1_io_out_r_bypass_1_2_data[15:0]   ), //o
    .io_out_r_bypass_1_2_load_store    (pes_0_1_io_out_r_bypass_1_2_load_store   ), //o
    .io_out_r_bypass_1_2_df_is_ws      (pes_0_1_io_out_r_bypass_1_2_df_is_ws     ), //o
    .io_out_r_bypass_1_2_stall         (pes_0_1_io_out_r_bypass_1_2_stall        ), //o
    .io_out_r_bypass_1_3_data          (pes_0_1_io_out_r_bypass_1_3_data[15:0]   ), //o
    .io_out_r_bypass_1_3_load_store    (pes_0_1_io_out_r_bypass_1_3_load_store   ), //o
    .io_out_r_bypass_1_3_df_is_ws      (pes_0_1_io_out_r_bypass_1_3_df_is_ws     ), //o
    .io_out_r_bypass_1_3_stall         (pes_0_1_io_out_r_bypass_1_3_stall        ), //o
    .io_out_r_input_from_bypass_0      (pes_0_1_io_out_r_input_from_bypass_0     ), //o
    .io_out_r_input_from_bypass_1      (pes_0_1_io_out_r_input_from_bypass_1     ), //o
    .io_in_c_data_0_data               (io_in_c_1_data_0_data[15:0]              ), //i
    .io_in_c_data_0_is_stationary      (io_in_c_1_data_0_is_stationary           ), //i
    .io_in_c_data_1_data               (io_in_c_1_data_1_data[15:0]              ), //i
    .io_in_c_data_1_is_stationary      (io_in_c_1_data_1_is_stationary           ), //i
    .io_in_c_data_2_data               (io_in_c_1_data_2_data[15:0]              ), //i
    .io_in_c_data_2_is_stationary      (io_in_c_1_data_2_is_stationary           ), //i
    .io_in_c_data_3_data               (io_in_c_1_data_3_data[15:0]              ), //i
    .io_in_c_data_3_is_stationary      (io_in_c_1_data_3_is_stationary           ), //i
    .io_in_c_bypass_0_0_data           (io_in_c_1_bypass_0_0_data[15:0]          ), //i
    .io_in_c_bypass_0_0_is_stationary  (io_in_c_1_bypass_0_0_is_stationary       ), //i
    .io_in_c_bypass_0_1_data           (io_in_c_1_bypass_0_1_data[15:0]          ), //i
    .io_in_c_bypass_0_1_is_stationary  (io_in_c_1_bypass_0_1_is_stationary       ), //i
    .io_in_c_bypass_0_2_data           (io_in_c_1_bypass_0_2_data[15:0]          ), //i
    .io_in_c_bypass_0_2_is_stationary  (io_in_c_1_bypass_0_2_is_stationary       ), //i
    .io_in_c_bypass_0_3_data           (io_in_c_1_bypass_0_3_data[15:0]          ), //i
    .io_in_c_bypass_0_3_is_stationary  (io_in_c_1_bypass_0_3_is_stationary       ), //i
    .io_in_c_bypass_1_0_data           (io_in_c_1_bypass_1_0_data[15:0]          ), //i
    .io_in_c_bypass_1_0_is_stationary  (io_in_c_1_bypass_1_0_is_stationary       ), //i
    .io_in_c_bypass_1_1_data           (io_in_c_1_bypass_1_1_data[15:0]          ), //i
    .io_in_c_bypass_1_1_is_stationary  (io_in_c_1_bypass_1_1_is_stationary       ), //i
    .io_in_c_bypass_1_2_data           (io_in_c_1_bypass_1_2_data[15:0]          ), //i
    .io_in_c_bypass_1_2_is_stationary  (io_in_c_1_bypass_1_2_is_stationary       ), //i
    .io_in_c_bypass_1_3_data           (io_in_c_1_bypass_1_3_data[15:0]          ), //i
    .io_in_c_bypass_1_3_is_stationary  (io_in_c_1_bypass_1_3_is_stationary       ), //i
    .io_in_c_input_from_bypass_0       (io_in_c_1_input_from_bypass_0            ), //i
    .io_in_c_input_from_bypass_1       (io_in_c_1_input_from_bypass_1            ), //i
    .io_out_c_data_0_data              (pes_0_1_io_out_c_data_0_data[15:0]       ), //o
    .io_out_c_data_0_is_stationary     (pes_0_1_io_out_c_data_0_is_stationary    ), //o
    .io_out_c_data_1_data              (pes_0_1_io_out_c_data_1_data[15:0]       ), //o
    .io_out_c_data_1_is_stationary     (pes_0_1_io_out_c_data_1_is_stationary    ), //o
    .io_out_c_data_2_data              (pes_0_1_io_out_c_data_2_data[15:0]       ), //o
    .io_out_c_data_2_is_stationary     (pes_0_1_io_out_c_data_2_is_stationary    ), //o
    .io_out_c_data_3_data              (pes_0_1_io_out_c_data_3_data[15:0]       ), //o
    .io_out_c_data_3_is_stationary     (pes_0_1_io_out_c_data_3_is_stationary    ), //o
    .io_out_c_bypass_0_0_data          (pes_0_1_io_out_c_bypass_0_0_data[15:0]   ), //o
    .io_out_c_bypass_0_0_is_stationary (pes_0_1_io_out_c_bypass_0_0_is_stationary), //o
    .io_out_c_bypass_0_1_data          (pes_0_1_io_out_c_bypass_0_1_data[15:0]   ), //o
    .io_out_c_bypass_0_1_is_stationary (pes_0_1_io_out_c_bypass_0_1_is_stationary), //o
    .io_out_c_bypass_0_2_data          (pes_0_1_io_out_c_bypass_0_2_data[15:0]   ), //o
    .io_out_c_bypass_0_2_is_stationary (pes_0_1_io_out_c_bypass_0_2_is_stationary), //o
    .io_out_c_bypass_0_3_data          (pes_0_1_io_out_c_bypass_0_3_data[15:0]   ), //o
    .io_out_c_bypass_0_3_is_stationary (pes_0_1_io_out_c_bypass_0_3_is_stationary), //o
    .io_out_c_bypass_1_0_data          (pes_0_1_io_out_c_bypass_1_0_data[15:0]   ), //o
    .io_out_c_bypass_1_0_is_stationary (pes_0_1_io_out_c_bypass_1_0_is_stationary), //o
    .io_out_c_bypass_1_1_data          (pes_0_1_io_out_c_bypass_1_1_data[15:0]   ), //o
    .io_out_c_bypass_1_1_is_stationary (pes_0_1_io_out_c_bypass_1_1_is_stationary), //o
    .io_out_c_bypass_1_2_data          (pes_0_1_io_out_c_bypass_1_2_data[15:0]   ), //o
    .io_out_c_bypass_1_2_is_stationary (pes_0_1_io_out_c_bypass_1_2_is_stationary), //o
    .io_out_c_bypass_1_3_data          (pes_0_1_io_out_c_bypass_1_3_data[15:0]   ), //o
    .io_out_c_bypass_1_3_is_stationary (pes_0_1_io_out_c_bypass_1_3_is_stationary), //o
    .io_out_c_input_from_bypass_0      (pes_0_1_io_out_c_input_from_bypass_0     ), //o
    .io_out_c_input_from_bypass_1      (pes_0_1_io_out_c_input_from_bypass_1     ), //o
    .clk                               (clk                                      ), //i
    .reset                             (reset                                    )  //i
  );
  CellSARA_7 pes_1_0 (
    .io_in_r_data_0_data               (io_in_r_1_data_0_data[15:0]              ), //i
    .io_in_r_data_0_load_store         (io_in_r_1_data_0_load_store              ), //i
    .io_in_r_data_0_df_is_ws           (io_in_r_1_data_0_df_is_ws                ), //i
    .io_in_r_data_0_stall              (io_in_r_1_data_0_stall                   ), //i
    .io_in_r_data_1_data               (io_in_r_1_data_1_data[15:0]              ), //i
    .io_in_r_data_1_load_store         (io_in_r_1_data_1_load_store              ), //i
    .io_in_r_data_1_df_is_ws           (io_in_r_1_data_1_df_is_ws                ), //i
    .io_in_r_data_1_stall              (io_in_r_1_data_1_stall                   ), //i
    .io_in_r_data_2_data               (io_in_r_1_data_2_data[15:0]              ), //i
    .io_in_r_data_2_load_store         (io_in_r_1_data_2_load_store              ), //i
    .io_in_r_data_2_df_is_ws           (io_in_r_1_data_2_df_is_ws                ), //i
    .io_in_r_data_2_stall              (io_in_r_1_data_2_stall                   ), //i
    .io_in_r_data_3_data               (io_in_r_1_data_3_data[15:0]              ), //i
    .io_in_r_data_3_load_store         (io_in_r_1_data_3_load_store              ), //i
    .io_in_r_data_3_df_is_ws           (io_in_r_1_data_3_df_is_ws                ), //i
    .io_in_r_data_3_stall              (io_in_r_1_data_3_stall                   ), //i
    .io_in_r_bypass_0_0_data           (io_in_r_1_bypass_0_0_data[15:0]          ), //i
    .io_in_r_bypass_0_0_load_store     (io_in_r_1_bypass_0_0_load_store          ), //i
    .io_in_r_bypass_0_0_df_is_ws       (io_in_r_1_bypass_0_0_df_is_ws            ), //i
    .io_in_r_bypass_0_0_stall          (io_in_r_1_bypass_0_0_stall               ), //i
    .io_in_r_bypass_0_1_data           (io_in_r_1_bypass_0_1_data[15:0]          ), //i
    .io_in_r_bypass_0_1_load_store     (io_in_r_1_bypass_0_1_load_store          ), //i
    .io_in_r_bypass_0_1_df_is_ws       (io_in_r_1_bypass_0_1_df_is_ws            ), //i
    .io_in_r_bypass_0_1_stall          (io_in_r_1_bypass_0_1_stall               ), //i
    .io_in_r_bypass_0_2_data           (io_in_r_1_bypass_0_2_data[15:0]          ), //i
    .io_in_r_bypass_0_2_load_store     (io_in_r_1_bypass_0_2_load_store          ), //i
    .io_in_r_bypass_0_2_df_is_ws       (io_in_r_1_bypass_0_2_df_is_ws            ), //i
    .io_in_r_bypass_0_2_stall          (io_in_r_1_bypass_0_2_stall               ), //i
    .io_in_r_bypass_0_3_data           (io_in_r_1_bypass_0_3_data[15:0]          ), //i
    .io_in_r_bypass_0_3_load_store     (io_in_r_1_bypass_0_3_load_store          ), //i
    .io_in_r_bypass_0_3_df_is_ws       (io_in_r_1_bypass_0_3_df_is_ws            ), //i
    .io_in_r_bypass_0_3_stall          (io_in_r_1_bypass_0_3_stall               ), //i
    .io_in_r_bypass_1_0_data           (io_in_r_1_bypass_1_0_data[15:0]          ), //i
    .io_in_r_bypass_1_0_load_store     (io_in_r_1_bypass_1_0_load_store          ), //i
    .io_in_r_bypass_1_0_df_is_ws       (io_in_r_1_bypass_1_0_df_is_ws            ), //i
    .io_in_r_bypass_1_0_stall          (io_in_r_1_bypass_1_0_stall               ), //i
    .io_in_r_bypass_1_1_data           (io_in_r_1_bypass_1_1_data[15:0]          ), //i
    .io_in_r_bypass_1_1_load_store     (io_in_r_1_bypass_1_1_load_store          ), //i
    .io_in_r_bypass_1_1_df_is_ws       (io_in_r_1_bypass_1_1_df_is_ws            ), //i
    .io_in_r_bypass_1_1_stall          (io_in_r_1_bypass_1_1_stall               ), //i
    .io_in_r_bypass_1_2_data           (io_in_r_1_bypass_1_2_data[15:0]          ), //i
    .io_in_r_bypass_1_2_load_store     (io_in_r_1_bypass_1_2_load_store          ), //i
    .io_in_r_bypass_1_2_df_is_ws       (io_in_r_1_bypass_1_2_df_is_ws            ), //i
    .io_in_r_bypass_1_2_stall          (io_in_r_1_bypass_1_2_stall               ), //i
    .io_in_r_bypass_1_3_data           (io_in_r_1_bypass_1_3_data[15:0]          ), //i
    .io_in_r_bypass_1_3_load_store     (io_in_r_1_bypass_1_3_load_store          ), //i
    .io_in_r_bypass_1_3_df_is_ws       (io_in_r_1_bypass_1_3_df_is_ws            ), //i
    .io_in_r_bypass_1_3_stall          (io_in_r_1_bypass_1_3_stall               ), //i
    .io_in_r_input_from_bypass_0       (io_in_r_1_input_from_bypass_0            ), //i
    .io_in_r_input_from_bypass_1       (io_in_r_1_input_from_bypass_1            ), //i
    .io_out_r_data_0_data              (pes_1_0_io_out_r_data_0_data[15:0]       ), //o
    .io_out_r_data_0_load_store        (pes_1_0_io_out_r_data_0_load_store       ), //o
    .io_out_r_data_0_df_is_ws          (pes_1_0_io_out_r_data_0_df_is_ws         ), //o
    .io_out_r_data_0_stall             (pes_1_0_io_out_r_data_0_stall            ), //o
    .io_out_r_data_1_data              (pes_1_0_io_out_r_data_1_data[15:0]       ), //o
    .io_out_r_data_1_load_store        (pes_1_0_io_out_r_data_1_load_store       ), //o
    .io_out_r_data_1_df_is_ws          (pes_1_0_io_out_r_data_1_df_is_ws         ), //o
    .io_out_r_data_1_stall             (pes_1_0_io_out_r_data_1_stall            ), //o
    .io_out_r_data_2_data              (pes_1_0_io_out_r_data_2_data[15:0]       ), //o
    .io_out_r_data_2_load_store        (pes_1_0_io_out_r_data_2_load_store       ), //o
    .io_out_r_data_2_df_is_ws          (pes_1_0_io_out_r_data_2_df_is_ws         ), //o
    .io_out_r_data_2_stall             (pes_1_0_io_out_r_data_2_stall            ), //o
    .io_out_r_data_3_data              (pes_1_0_io_out_r_data_3_data[15:0]       ), //o
    .io_out_r_data_3_load_store        (pes_1_0_io_out_r_data_3_load_store       ), //o
    .io_out_r_data_3_df_is_ws          (pes_1_0_io_out_r_data_3_df_is_ws         ), //o
    .io_out_r_data_3_stall             (pes_1_0_io_out_r_data_3_stall            ), //o
    .io_out_r_bypass_0_0_data          (pes_1_0_io_out_r_bypass_0_0_data[15:0]   ), //o
    .io_out_r_bypass_0_0_load_store    (pes_1_0_io_out_r_bypass_0_0_load_store   ), //o
    .io_out_r_bypass_0_0_df_is_ws      (pes_1_0_io_out_r_bypass_0_0_df_is_ws     ), //o
    .io_out_r_bypass_0_0_stall         (pes_1_0_io_out_r_bypass_0_0_stall        ), //o
    .io_out_r_bypass_0_1_data          (pes_1_0_io_out_r_bypass_0_1_data[15:0]   ), //o
    .io_out_r_bypass_0_1_load_store    (pes_1_0_io_out_r_bypass_0_1_load_store   ), //o
    .io_out_r_bypass_0_1_df_is_ws      (pes_1_0_io_out_r_bypass_0_1_df_is_ws     ), //o
    .io_out_r_bypass_0_1_stall         (pes_1_0_io_out_r_bypass_0_1_stall        ), //o
    .io_out_r_bypass_0_2_data          (pes_1_0_io_out_r_bypass_0_2_data[15:0]   ), //o
    .io_out_r_bypass_0_2_load_store    (pes_1_0_io_out_r_bypass_0_2_load_store   ), //o
    .io_out_r_bypass_0_2_df_is_ws      (pes_1_0_io_out_r_bypass_0_2_df_is_ws     ), //o
    .io_out_r_bypass_0_2_stall         (pes_1_0_io_out_r_bypass_0_2_stall        ), //o
    .io_out_r_bypass_0_3_data          (pes_1_0_io_out_r_bypass_0_3_data[15:0]   ), //o
    .io_out_r_bypass_0_3_load_store    (pes_1_0_io_out_r_bypass_0_3_load_store   ), //o
    .io_out_r_bypass_0_3_df_is_ws      (pes_1_0_io_out_r_bypass_0_3_df_is_ws     ), //o
    .io_out_r_bypass_0_3_stall         (pes_1_0_io_out_r_bypass_0_3_stall        ), //o
    .io_out_r_bypass_1_0_data          (pes_1_0_io_out_r_bypass_1_0_data[15:0]   ), //o
    .io_out_r_bypass_1_0_load_store    (pes_1_0_io_out_r_bypass_1_0_load_store   ), //o
    .io_out_r_bypass_1_0_df_is_ws      (pes_1_0_io_out_r_bypass_1_0_df_is_ws     ), //o
    .io_out_r_bypass_1_0_stall         (pes_1_0_io_out_r_bypass_1_0_stall        ), //o
    .io_out_r_bypass_1_1_data          (pes_1_0_io_out_r_bypass_1_1_data[15:0]   ), //o
    .io_out_r_bypass_1_1_load_store    (pes_1_0_io_out_r_bypass_1_1_load_store   ), //o
    .io_out_r_bypass_1_1_df_is_ws      (pes_1_0_io_out_r_bypass_1_1_df_is_ws     ), //o
    .io_out_r_bypass_1_1_stall         (pes_1_0_io_out_r_bypass_1_1_stall        ), //o
    .io_out_r_bypass_1_2_data          (pes_1_0_io_out_r_bypass_1_2_data[15:0]   ), //o
    .io_out_r_bypass_1_2_load_store    (pes_1_0_io_out_r_bypass_1_2_load_store   ), //o
    .io_out_r_bypass_1_2_df_is_ws      (pes_1_0_io_out_r_bypass_1_2_df_is_ws     ), //o
    .io_out_r_bypass_1_2_stall         (pes_1_0_io_out_r_bypass_1_2_stall        ), //o
    .io_out_r_bypass_1_3_data          (pes_1_0_io_out_r_bypass_1_3_data[15:0]   ), //o
    .io_out_r_bypass_1_3_load_store    (pes_1_0_io_out_r_bypass_1_3_load_store   ), //o
    .io_out_r_bypass_1_3_df_is_ws      (pes_1_0_io_out_r_bypass_1_3_df_is_ws     ), //o
    .io_out_r_bypass_1_3_stall         (pes_1_0_io_out_r_bypass_1_3_stall        ), //o
    .io_out_r_input_from_bypass_0      (pes_1_0_io_out_r_input_from_bypass_0     ), //o
    .io_out_r_input_from_bypass_1      (pes_1_0_io_out_r_input_from_bypass_1     ), //o
    .io_in_c_data_0_data               (pes_0_0_io_out_c_data_0_data[15:0]       ), //i
    .io_in_c_data_0_is_stationary      (pes_0_0_io_out_c_data_0_is_stationary    ), //i
    .io_in_c_data_1_data               (pes_0_0_io_out_c_data_1_data[15:0]       ), //i
    .io_in_c_data_1_is_stationary      (pes_0_0_io_out_c_data_1_is_stationary    ), //i
    .io_in_c_data_2_data               (pes_0_0_io_out_c_data_2_data[15:0]       ), //i
    .io_in_c_data_2_is_stationary      (pes_0_0_io_out_c_data_2_is_stationary    ), //i
    .io_in_c_data_3_data               (pes_0_0_io_out_c_data_3_data[15:0]       ), //i
    .io_in_c_data_3_is_stationary      (pes_0_0_io_out_c_data_3_is_stationary    ), //i
    .io_in_c_bypass_0_0_data           (pes_0_0_io_out_c_bypass_0_0_data[15:0]   ), //i
    .io_in_c_bypass_0_0_is_stationary  (pes_0_0_io_out_c_bypass_0_0_is_stationary), //i
    .io_in_c_bypass_0_1_data           (pes_0_0_io_out_c_bypass_0_1_data[15:0]   ), //i
    .io_in_c_bypass_0_1_is_stationary  (pes_0_0_io_out_c_bypass_0_1_is_stationary), //i
    .io_in_c_bypass_0_2_data           (pes_0_0_io_out_c_bypass_0_2_data[15:0]   ), //i
    .io_in_c_bypass_0_2_is_stationary  (pes_0_0_io_out_c_bypass_0_2_is_stationary), //i
    .io_in_c_bypass_0_3_data           (pes_0_0_io_out_c_bypass_0_3_data[15:0]   ), //i
    .io_in_c_bypass_0_3_is_stationary  (pes_0_0_io_out_c_bypass_0_3_is_stationary), //i
    .io_in_c_bypass_1_0_data           (pes_0_0_io_out_c_bypass_1_0_data[15:0]   ), //i
    .io_in_c_bypass_1_0_is_stationary  (pes_0_0_io_out_c_bypass_1_0_is_stationary), //i
    .io_in_c_bypass_1_1_data           (pes_0_0_io_out_c_bypass_1_1_data[15:0]   ), //i
    .io_in_c_bypass_1_1_is_stationary  (pes_0_0_io_out_c_bypass_1_1_is_stationary), //i
    .io_in_c_bypass_1_2_data           (pes_0_0_io_out_c_bypass_1_2_data[15:0]   ), //i
    .io_in_c_bypass_1_2_is_stationary  (pes_0_0_io_out_c_bypass_1_2_is_stationary), //i
    .io_in_c_bypass_1_3_data           (pes_0_0_io_out_c_bypass_1_3_data[15:0]   ), //i
    .io_in_c_bypass_1_3_is_stationary  (pes_0_0_io_out_c_bypass_1_3_is_stationary), //i
    .io_in_c_input_from_bypass_0       (pes_0_0_io_out_c_input_from_bypass_0     ), //i
    .io_in_c_input_from_bypass_1       (pes_0_0_io_out_c_input_from_bypass_1     ), //i
    .io_out_c_data_0_data              (pes_1_0_io_out_c_data_0_data[15:0]       ), //o
    .io_out_c_data_0_is_stationary     (pes_1_0_io_out_c_data_0_is_stationary    ), //o
    .io_out_c_data_1_data              (pes_1_0_io_out_c_data_1_data[15:0]       ), //o
    .io_out_c_data_1_is_stationary     (pes_1_0_io_out_c_data_1_is_stationary    ), //o
    .io_out_c_data_2_data              (pes_1_0_io_out_c_data_2_data[15:0]       ), //o
    .io_out_c_data_2_is_stationary     (pes_1_0_io_out_c_data_2_is_stationary    ), //o
    .io_out_c_data_3_data              (pes_1_0_io_out_c_data_3_data[15:0]       ), //o
    .io_out_c_data_3_is_stationary     (pes_1_0_io_out_c_data_3_is_stationary    ), //o
    .io_out_c_bypass_0_0_data          (pes_1_0_io_out_c_bypass_0_0_data[15:0]   ), //o
    .io_out_c_bypass_0_0_is_stationary (pes_1_0_io_out_c_bypass_0_0_is_stationary), //o
    .io_out_c_bypass_0_1_data          (pes_1_0_io_out_c_bypass_0_1_data[15:0]   ), //o
    .io_out_c_bypass_0_1_is_stationary (pes_1_0_io_out_c_bypass_0_1_is_stationary), //o
    .io_out_c_bypass_0_2_data          (pes_1_0_io_out_c_bypass_0_2_data[15:0]   ), //o
    .io_out_c_bypass_0_2_is_stationary (pes_1_0_io_out_c_bypass_0_2_is_stationary), //o
    .io_out_c_bypass_0_3_data          (pes_1_0_io_out_c_bypass_0_3_data[15:0]   ), //o
    .io_out_c_bypass_0_3_is_stationary (pes_1_0_io_out_c_bypass_0_3_is_stationary), //o
    .io_out_c_bypass_1_0_data          (pes_1_0_io_out_c_bypass_1_0_data[15:0]   ), //o
    .io_out_c_bypass_1_0_is_stationary (pes_1_0_io_out_c_bypass_1_0_is_stationary), //o
    .io_out_c_bypass_1_1_data          (pes_1_0_io_out_c_bypass_1_1_data[15:0]   ), //o
    .io_out_c_bypass_1_1_is_stationary (pes_1_0_io_out_c_bypass_1_1_is_stationary), //o
    .io_out_c_bypass_1_2_data          (pes_1_0_io_out_c_bypass_1_2_data[15:0]   ), //o
    .io_out_c_bypass_1_2_is_stationary (pes_1_0_io_out_c_bypass_1_2_is_stationary), //o
    .io_out_c_bypass_1_3_data          (pes_1_0_io_out_c_bypass_1_3_data[15:0]   ), //o
    .io_out_c_bypass_1_3_is_stationary (pes_1_0_io_out_c_bypass_1_3_is_stationary), //o
    .io_out_c_input_from_bypass_0      (pes_1_0_io_out_c_input_from_bypass_0     ), //o
    .io_out_c_input_from_bypass_1      (pes_1_0_io_out_c_input_from_bypass_1     ), //o
    .clk                               (clk                                      ), //i
    .reset                             (reset                                    )  //i
  );
  CellSARA_7 pes_1_1 (
    .io_in_r_data_0_data               (pes_1_0_io_out_r_data_0_data[15:0]       ), //i
    .io_in_r_data_0_load_store         (pes_1_0_io_out_r_data_0_load_store       ), //i
    .io_in_r_data_0_df_is_ws           (pes_1_0_io_out_r_data_0_df_is_ws         ), //i
    .io_in_r_data_0_stall              (pes_1_0_io_out_r_data_0_stall            ), //i
    .io_in_r_data_1_data               (pes_1_0_io_out_r_data_1_data[15:0]       ), //i
    .io_in_r_data_1_load_store         (pes_1_0_io_out_r_data_1_load_store       ), //i
    .io_in_r_data_1_df_is_ws           (pes_1_0_io_out_r_data_1_df_is_ws         ), //i
    .io_in_r_data_1_stall              (pes_1_0_io_out_r_data_1_stall            ), //i
    .io_in_r_data_2_data               (pes_1_0_io_out_r_data_2_data[15:0]       ), //i
    .io_in_r_data_2_load_store         (pes_1_0_io_out_r_data_2_load_store       ), //i
    .io_in_r_data_2_df_is_ws           (pes_1_0_io_out_r_data_2_df_is_ws         ), //i
    .io_in_r_data_2_stall              (pes_1_0_io_out_r_data_2_stall            ), //i
    .io_in_r_data_3_data               (pes_1_0_io_out_r_data_3_data[15:0]       ), //i
    .io_in_r_data_3_load_store         (pes_1_0_io_out_r_data_3_load_store       ), //i
    .io_in_r_data_3_df_is_ws           (pes_1_0_io_out_r_data_3_df_is_ws         ), //i
    .io_in_r_data_3_stall              (pes_1_0_io_out_r_data_3_stall            ), //i
    .io_in_r_bypass_0_0_data           (pes_1_0_io_out_r_bypass_0_0_data[15:0]   ), //i
    .io_in_r_bypass_0_0_load_store     (pes_1_0_io_out_r_bypass_0_0_load_store   ), //i
    .io_in_r_bypass_0_0_df_is_ws       (pes_1_0_io_out_r_bypass_0_0_df_is_ws     ), //i
    .io_in_r_bypass_0_0_stall          (pes_1_0_io_out_r_bypass_0_0_stall        ), //i
    .io_in_r_bypass_0_1_data           (pes_1_0_io_out_r_bypass_0_1_data[15:0]   ), //i
    .io_in_r_bypass_0_1_load_store     (pes_1_0_io_out_r_bypass_0_1_load_store   ), //i
    .io_in_r_bypass_0_1_df_is_ws       (pes_1_0_io_out_r_bypass_0_1_df_is_ws     ), //i
    .io_in_r_bypass_0_1_stall          (pes_1_0_io_out_r_bypass_0_1_stall        ), //i
    .io_in_r_bypass_0_2_data           (pes_1_0_io_out_r_bypass_0_2_data[15:0]   ), //i
    .io_in_r_bypass_0_2_load_store     (pes_1_0_io_out_r_bypass_0_2_load_store   ), //i
    .io_in_r_bypass_0_2_df_is_ws       (pes_1_0_io_out_r_bypass_0_2_df_is_ws     ), //i
    .io_in_r_bypass_0_2_stall          (pes_1_0_io_out_r_bypass_0_2_stall        ), //i
    .io_in_r_bypass_0_3_data           (pes_1_0_io_out_r_bypass_0_3_data[15:0]   ), //i
    .io_in_r_bypass_0_3_load_store     (pes_1_0_io_out_r_bypass_0_3_load_store   ), //i
    .io_in_r_bypass_0_3_df_is_ws       (pes_1_0_io_out_r_bypass_0_3_df_is_ws     ), //i
    .io_in_r_bypass_0_3_stall          (pes_1_0_io_out_r_bypass_0_3_stall        ), //i
    .io_in_r_bypass_1_0_data           (pes_1_0_io_out_r_bypass_1_0_data[15:0]   ), //i
    .io_in_r_bypass_1_0_load_store     (pes_1_0_io_out_r_bypass_1_0_load_store   ), //i
    .io_in_r_bypass_1_0_df_is_ws       (pes_1_0_io_out_r_bypass_1_0_df_is_ws     ), //i
    .io_in_r_bypass_1_0_stall          (pes_1_0_io_out_r_bypass_1_0_stall        ), //i
    .io_in_r_bypass_1_1_data           (pes_1_0_io_out_r_bypass_1_1_data[15:0]   ), //i
    .io_in_r_bypass_1_1_load_store     (pes_1_0_io_out_r_bypass_1_1_load_store   ), //i
    .io_in_r_bypass_1_1_df_is_ws       (pes_1_0_io_out_r_bypass_1_1_df_is_ws     ), //i
    .io_in_r_bypass_1_1_stall          (pes_1_0_io_out_r_bypass_1_1_stall        ), //i
    .io_in_r_bypass_1_2_data           (pes_1_0_io_out_r_bypass_1_2_data[15:0]   ), //i
    .io_in_r_bypass_1_2_load_store     (pes_1_0_io_out_r_bypass_1_2_load_store   ), //i
    .io_in_r_bypass_1_2_df_is_ws       (pes_1_0_io_out_r_bypass_1_2_df_is_ws     ), //i
    .io_in_r_bypass_1_2_stall          (pes_1_0_io_out_r_bypass_1_2_stall        ), //i
    .io_in_r_bypass_1_3_data           (pes_1_0_io_out_r_bypass_1_3_data[15:0]   ), //i
    .io_in_r_bypass_1_3_load_store     (pes_1_0_io_out_r_bypass_1_3_load_store   ), //i
    .io_in_r_bypass_1_3_df_is_ws       (pes_1_0_io_out_r_bypass_1_3_df_is_ws     ), //i
    .io_in_r_bypass_1_3_stall          (pes_1_0_io_out_r_bypass_1_3_stall        ), //i
    .io_in_r_input_from_bypass_0       (pes_1_0_io_out_r_input_from_bypass_0     ), //i
    .io_in_r_input_from_bypass_1       (pes_1_0_io_out_r_input_from_bypass_1     ), //i
    .io_out_r_data_0_data              (pes_1_1_io_out_r_data_0_data[15:0]       ), //o
    .io_out_r_data_0_load_store        (pes_1_1_io_out_r_data_0_load_store       ), //o
    .io_out_r_data_0_df_is_ws          (pes_1_1_io_out_r_data_0_df_is_ws         ), //o
    .io_out_r_data_0_stall             (pes_1_1_io_out_r_data_0_stall            ), //o
    .io_out_r_data_1_data              (pes_1_1_io_out_r_data_1_data[15:0]       ), //o
    .io_out_r_data_1_load_store        (pes_1_1_io_out_r_data_1_load_store       ), //o
    .io_out_r_data_1_df_is_ws          (pes_1_1_io_out_r_data_1_df_is_ws         ), //o
    .io_out_r_data_1_stall             (pes_1_1_io_out_r_data_1_stall            ), //o
    .io_out_r_data_2_data              (pes_1_1_io_out_r_data_2_data[15:0]       ), //o
    .io_out_r_data_2_load_store        (pes_1_1_io_out_r_data_2_load_store       ), //o
    .io_out_r_data_2_df_is_ws          (pes_1_1_io_out_r_data_2_df_is_ws         ), //o
    .io_out_r_data_2_stall             (pes_1_1_io_out_r_data_2_stall            ), //o
    .io_out_r_data_3_data              (pes_1_1_io_out_r_data_3_data[15:0]       ), //o
    .io_out_r_data_3_load_store        (pes_1_1_io_out_r_data_3_load_store       ), //o
    .io_out_r_data_3_df_is_ws          (pes_1_1_io_out_r_data_3_df_is_ws         ), //o
    .io_out_r_data_3_stall             (pes_1_1_io_out_r_data_3_stall            ), //o
    .io_out_r_bypass_0_0_data          (pes_1_1_io_out_r_bypass_0_0_data[15:0]   ), //o
    .io_out_r_bypass_0_0_load_store    (pes_1_1_io_out_r_bypass_0_0_load_store   ), //o
    .io_out_r_bypass_0_0_df_is_ws      (pes_1_1_io_out_r_bypass_0_0_df_is_ws     ), //o
    .io_out_r_bypass_0_0_stall         (pes_1_1_io_out_r_bypass_0_0_stall        ), //o
    .io_out_r_bypass_0_1_data          (pes_1_1_io_out_r_bypass_0_1_data[15:0]   ), //o
    .io_out_r_bypass_0_1_load_store    (pes_1_1_io_out_r_bypass_0_1_load_store   ), //o
    .io_out_r_bypass_0_1_df_is_ws      (pes_1_1_io_out_r_bypass_0_1_df_is_ws     ), //o
    .io_out_r_bypass_0_1_stall         (pes_1_1_io_out_r_bypass_0_1_stall        ), //o
    .io_out_r_bypass_0_2_data          (pes_1_1_io_out_r_bypass_0_2_data[15:0]   ), //o
    .io_out_r_bypass_0_2_load_store    (pes_1_1_io_out_r_bypass_0_2_load_store   ), //o
    .io_out_r_bypass_0_2_df_is_ws      (pes_1_1_io_out_r_bypass_0_2_df_is_ws     ), //o
    .io_out_r_bypass_0_2_stall         (pes_1_1_io_out_r_bypass_0_2_stall        ), //o
    .io_out_r_bypass_0_3_data          (pes_1_1_io_out_r_bypass_0_3_data[15:0]   ), //o
    .io_out_r_bypass_0_3_load_store    (pes_1_1_io_out_r_bypass_0_3_load_store   ), //o
    .io_out_r_bypass_0_3_df_is_ws      (pes_1_1_io_out_r_bypass_0_3_df_is_ws     ), //o
    .io_out_r_bypass_0_3_stall         (pes_1_1_io_out_r_bypass_0_3_stall        ), //o
    .io_out_r_bypass_1_0_data          (pes_1_1_io_out_r_bypass_1_0_data[15:0]   ), //o
    .io_out_r_bypass_1_0_load_store    (pes_1_1_io_out_r_bypass_1_0_load_store   ), //o
    .io_out_r_bypass_1_0_df_is_ws      (pes_1_1_io_out_r_bypass_1_0_df_is_ws     ), //o
    .io_out_r_bypass_1_0_stall         (pes_1_1_io_out_r_bypass_1_0_stall        ), //o
    .io_out_r_bypass_1_1_data          (pes_1_1_io_out_r_bypass_1_1_data[15:0]   ), //o
    .io_out_r_bypass_1_1_load_store    (pes_1_1_io_out_r_bypass_1_1_load_store   ), //o
    .io_out_r_bypass_1_1_df_is_ws      (pes_1_1_io_out_r_bypass_1_1_df_is_ws     ), //o
    .io_out_r_bypass_1_1_stall         (pes_1_1_io_out_r_bypass_1_1_stall        ), //o
    .io_out_r_bypass_1_2_data          (pes_1_1_io_out_r_bypass_1_2_data[15:0]   ), //o
    .io_out_r_bypass_1_2_load_store    (pes_1_1_io_out_r_bypass_1_2_load_store   ), //o
    .io_out_r_bypass_1_2_df_is_ws      (pes_1_1_io_out_r_bypass_1_2_df_is_ws     ), //o
    .io_out_r_bypass_1_2_stall         (pes_1_1_io_out_r_bypass_1_2_stall        ), //o
    .io_out_r_bypass_1_3_data          (pes_1_1_io_out_r_bypass_1_3_data[15:0]   ), //o
    .io_out_r_bypass_1_3_load_store    (pes_1_1_io_out_r_bypass_1_3_load_store   ), //o
    .io_out_r_bypass_1_3_df_is_ws      (pes_1_1_io_out_r_bypass_1_3_df_is_ws     ), //o
    .io_out_r_bypass_1_3_stall         (pes_1_1_io_out_r_bypass_1_3_stall        ), //o
    .io_out_r_input_from_bypass_0      (pes_1_1_io_out_r_input_from_bypass_0     ), //o
    .io_out_r_input_from_bypass_1      (pes_1_1_io_out_r_input_from_bypass_1     ), //o
    .io_in_c_data_0_data               (pes_0_1_io_out_c_data_0_data[15:0]       ), //i
    .io_in_c_data_0_is_stationary      (pes_0_1_io_out_c_data_0_is_stationary    ), //i
    .io_in_c_data_1_data               (pes_0_1_io_out_c_data_1_data[15:0]       ), //i
    .io_in_c_data_1_is_stationary      (pes_0_1_io_out_c_data_1_is_stationary    ), //i
    .io_in_c_data_2_data               (pes_0_1_io_out_c_data_2_data[15:0]       ), //i
    .io_in_c_data_2_is_stationary      (pes_0_1_io_out_c_data_2_is_stationary    ), //i
    .io_in_c_data_3_data               (pes_0_1_io_out_c_data_3_data[15:0]       ), //i
    .io_in_c_data_3_is_stationary      (pes_0_1_io_out_c_data_3_is_stationary    ), //i
    .io_in_c_bypass_0_0_data           (pes_0_1_io_out_c_bypass_0_0_data[15:0]   ), //i
    .io_in_c_bypass_0_0_is_stationary  (pes_0_1_io_out_c_bypass_0_0_is_stationary), //i
    .io_in_c_bypass_0_1_data           (pes_0_1_io_out_c_bypass_0_1_data[15:0]   ), //i
    .io_in_c_bypass_0_1_is_stationary  (pes_0_1_io_out_c_bypass_0_1_is_stationary), //i
    .io_in_c_bypass_0_2_data           (pes_0_1_io_out_c_bypass_0_2_data[15:0]   ), //i
    .io_in_c_bypass_0_2_is_stationary  (pes_0_1_io_out_c_bypass_0_2_is_stationary), //i
    .io_in_c_bypass_0_3_data           (pes_0_1_io_out_c_bypass_0_3_data[15:0]   ), //i
    .io_in_c_bypass_0_3_is_stationary  (pes_0_1_io_out_c_bypass_0_3_is_stationary), //i
    .io_in_c_bypass_1_0_data           (pes_0_1_io_out_c_bypass_1_0_data[15:0]   ), //i
    .io_in_c_bypass_1_0_is_stationary  (pes_0_1_io_out_c_bypass_1_0_is_stationary), //i
    .io_in_c_bypass_1_1_data           (pes_0_1_io_out_c_bypass_1_1_data[15:0]   ), //i
    .io_in_c_bypass_1_1_is_stationary  (pes_0_1_io_out_c_bypass_1_1_is_stationary), //i
    .io_in_c_bypass_1_2_data           (pes_0_1_io_out_c_bypass_1_2_data[15:0]   ), //i
    .io_in_c_bypass_1_2_is_stationary  (pes_0_1_io_out_c_bypass_1_2_is_stationary), //i
    .io_in_c_bypass_1_3_data           (pes_0_1_io_out_c_bypass_1_3_data[15:0]   ), //i
    .io_in_c_bypass_1_3_is_stationary  (pes_0_1_io_out_c_bypass_1_3_is_stationary), //i
    .io_in_c_input_from_bypass_0       (pes_0_1_io_out_c_input_from_bypass_0     ), //i
    .io_in_c_input_from_bypass_1       (pes_0_1_io_out_c_input_from_bypass_1     ), //i
    .io_out_c_data_0_data              (pes_1_1_io_out_c_data_0_data[15:0]       ), //o
    .io_out_c_data_0_is_stationary     (pes_1_1_io_out_c_data_0_is_stationary    ), //o
    .io_out_c_data_1_data              (pes_1_1_io_out_c_data_1_data[15:0]       ), //o
    .io_out_c_data_1_is_stationary     (pes_1_1_io_out_c_data_1_is_stationary    ), //o
    .io_out_c_data_2_data              (pes_1_1_io_out_c_data_2_data[15:0]       ), //o
    .io_out_c_data_2_is_stationary     (pes_1_1_io_out_c_data_2_is_stationary    ), //o
    .io_out_c_data_3_data              (pes_1_1_io_out_c_data_3_data[15:0]       ), //o
    .io_out_c_data_3_is_stationary     (pes_1_1_io_out_c_data_3_is_stationary    ), //o
    .io_out_c_bypass_0_0_data          (pes_1_1_io_out_c_bypass_0_0_data[15:0]   ), //o
    .io_out_c_bypass_0_0_is_stationary (pes_1_1_io_out_c_bypass_0_0_is_stationary), //o
    .io_out_c_bypass_0_1_data          (pes_1_1_io_out_c_bypass_0_1_data[15:0]   ), //o
    .io_out_c_bypass_0_1_is_stationary (pes_1_1_io_out_c_bypass_0_1_is_stationary), //o
    .io_out_c_bypass_0_2_data          (pes_1_1_io_out_c_bypass_0_2_data[15:0]   ), //o
    .io_out_c_bypass_0_2_is_stationary (pes_1_1_io_out_c_bypass_0_2_is_stationary), //o
    .io_out_c_bypass_0_3_data          (pes_1_1_io_out_c_bypass_0_3_data[15:0]   ), //o
    .io_out_c_bypass_0_3_is_stationary (pes_1_1_io_out_c_bypass_0_3_is_stationary), //o
    .io_out_c_bypass_1_0_data          (pes_1_1_io_out_c_bypass_1_0_data[15:0]   ), //o
    .io_out_c_bypass_1_0_is_stationary (pes_1_1_io_out_c_bypass_1_0_is_stationary), //o
    .io_out_c_bypass_1_1_data          (pes_1_1_io_out_c_bypass_1_1_data[15:0]   ), //o
    .io_out_c_bypass_1_1_is_stationary (pes_1_1_io_out_c_bypass_1_1_is_stationary), //o
    .io_out_c_bypass_1_2_data          (pes_1_1_io_out_c_bypass_1_2_data[15:0]   ), //o
    .io_out_c_bypass_1_2_is_stationary (pes_1_1_io_out_c_bypass_1_2_is_stationary), //o
    .io_out_c_bypass_1_3_data          (pes_1_1_io_out_c_bypass_1_3_data[15:0]   ), //o
    .io_out_c_bypass_1_3_is_stationary (pes_1_1_io_out_c_bypass_1_3_is_stationary), //o
    .io_out_c_input_from_bypass_0      (pes_1_1_io_out_c_input_from_bypass_0     ), //o
    .io_out_c_input_from_bypass_1      (pes_1_1_io_out_c_input_from_bypass_1     ), //o
    .clk                               (clk                                      ), //i
    .reset                             (reset                                    )  //i
  );
  CellSARA_7 cellSARA_8 (
    .io_in_r_data_0_data               (cellSARA_8_io_in_r_data_0_data[15:0]        ), //i
    .io_in_r_data_0_load_store         (cellSARA_8_io_in_r_data_0_load_store        ), //i
    .io_in_r_data_0_df_is_ws           (cellSARA_8_io_in_r_data_0_df_is_ws          ), //i
    .io_in_r_data_0_stall              (cellSARA_8_io_in_r_data_0_stall             ), //i
    .io_in_r_data_1_data               (cellSARA_8_io_in_r_data_1_data[15:0]        ), //i
    .io_in_r_data_1_load_store         (cellSARA_8_io_in_r_data_1_load_store        ), //i
    .io_in_r_data_1_df_is_ws           (cellSARA_8_io_in_r_data_1_df_is_ws          ), //i
    .io_in_r_data_1_stall              (cellSARA_8_io_in_r_data_1_stall             ), //i
    .io_in_r_data_2_data               (cellSARA_8_io_in_r_data_2_data[15:0]        ), //i
    .io_in_r_data_2_load_store         (cellSARA_8_io_in_r_data_2_load_store        ), //i
    .io_in_r_data_2_df_is_ws           (cellSARA_8_io_in_r_data_2_df_is_ws          ), //i
    .io_in_r_data_2_stall              (cellSARA_8_io_in_r_data_2_stall             ), //i
    .io_in_r_data_3_data               (cellSARA_8_io_in_r_data_3_data[15:0]        ), //i
    .io_in_r_data_3_load_store         (cellSARA_8_io_in_r_data_3_load_store        ), //i
    .io_in_r_data_3_df_is_ws           (cellSARA_8_io_in_r_data_3_df_is_ws          ), //i
    .io_in_r_data_3_stall              (cellSARA_8_io_in_r_data_3_stall             ), //i
    .io_in_r_bypass_0_0_data           (cellSARA_8_io_in_r_bypass_0_0_data[15:0]    ), //i
    .io_in_r_bypass_0_0_load_store     (cellSARA_8_io_in_r_bypass_0_0_load_store    ), //i
    .io_in_r_bypass_0_0_df_is_ws       (cellSARA_8_io_in_r_bypass_0_0_df_is_ws      ), //i
    .io_in_r_bypass_0_0_stall          (cellSARA_8_io_in_r_bypass_0_0_stall         ), //i
    .io_in_r_bypass_0_1_data           (cellSARA_8_io_in_r_bypass_0_1_data[15:0]    ), //i
    .io_in_r_bypass_0_1_load_store     (cellSARA_8_io_in_r_bypass_0_1_load_store    ), //i
    .io_in_r_bypass_0_1_df_is_ws       (cellSARA_8_io_in_r_bypass_0_1_df_is_ws      ), //i
    .io_in_r_bypass_0_1_stall          (cellSARA_8_io_in_r_bypass_0_1_stall         ), //i
    .io_in_r_bypass_0_2_data           (cellSARA_8_io_in_r_bypass_0_2_data[15:0]    ), //i
    .io_in_r_bypass_0_2_load_store     (cellSARA_8_io_in_r_bypass_0_2_load_store    ), //i
    .io_in_r_bypass_0_2_df_is_ws       (cellSARA_8_io_in_r_bypass_0_2_df_is_ws      ), //i
    .io_in_r_bypass_0_2_stall          (cellSARA_8_io_in_r_bypass_0_2_stall         ), //i
    .io_in_r_bypass_0_3_data           (cellSARA_8_io_in_r_bypass_0_3_data[15:0]    ), //i
    .io_in_r_bypass_0_3_load_store     (cellSARA_8_io_in_r_bypass_0_3_load_store    ), //i
    .io_in_r_bypass_0_3_df_is_ws       (cellSARA_8_io_in_r_bypass_0_3_df_is_ws      ), //i
    .io_in_r_bypass_0_3_stall          (cellSARA_8_io_in_r_bypass_0_3_stall         ), //i
    .io_in_r_bypass_1_0_data           (cellSARA_8_io_in_r_bypass_1_0_data[15:0]    ), //i
    .io_in_r_bypass_1_0_load_store     (cellSARA_8_io_in_r_bypass_1_0_load_store    ), //i
    .io_in_r_bypass_1_0_df_is_ws       (cellSARA_8_io_in_r_bypass_1_0_df_is_ws      ), //i
    .io_in_r_bypass_1_0_stall          (cellSARA_8_io_in_r_bypass_1_0_stall         ), //i
    .io_in_r_bypass_1_1_data           (cellSARA_8_io_in_r_bypass_1_1_data[15:0]    ), //i
    .io_in_r_bypass_1_1_load_store     (cellSARA_8_io_in_r_bypass_1_1_load_store    ), //i
    .io_in_r_bypass_1_1_df_is_ws       (cellSARA_8_io_in_r_bypass_1_1_df_is_ws      ), //i
    .io_in_r_bypass_1_1_stall          (cellSARA_8_io_in_r_bypass_1_1_stall         ), //i
    .io_in_r_bypass_1_2_data           (cellSARA_8_io_in_r_bypass_1_2_data[15:0]    ), //i
    .io_in_r_bypass_1_2_load_store     (cellSARA_8_io_in_r_bypass_1_2_load_store    ), //i
    .io_in_r_bypass_1_2_df_is_ws       (cellSARA_8_io_in_r_bypass_1_2_df_is_ws      ), //i
    .io_in_r_bypass_1_2_stall          (cellSARA_8_io_in_r_bypass_1_2_stall         ), //i
    .io_in_r_bypass_1_3_data           (cellSARA_8_io_in_r_bypass_1_3_data[15:0]    ), //i
    .io_in_r_bypass_1_3_load_store     (cellSARA_8_io_in_r_bypass_1_3_load_store    ), //i
    .io_in_r_bypass_1_3_df_is_ws       (cellSARA_8_io_in_r_bypass_1_3_df_is_ws      ), //i
    .io_in_r_bypass_1_3_stall          (cellSARA_8_io_in_r_bypass_1_3_stall         ), //i
    .io_in_r_input_from_bypass_0       (cellSARA_8_io_in_r_input_from_bypass_0      ), //i
    .io_in_r_input_from_bypass_1       (cellSARA_8_io_in_r_input_from_bypass_1      ), //i
    .io_out_r_data_0_data              (cellSARA_8_io_out_r_data_0_data[15:0]       ), //o
    .io_out_r_data_0_load_store        (cellSARA_8_io_out_r_data_0_load_store       ), //o
    .io_out_r_data_0_df_is_ws          (cellSARA_8_io_out_r_data_0_df_is_ws         ), //o
    .io_out_r_data_0_stall             (cellSARA_8_io_out_r_data_0_stall            ), //o
    .io_out_r_data_1_data              (cellSARA_8_io_out_r_data_1_data[15:0]       ), //o
    .io_out_r_data_1_load_store        (cellSARA_8_io_out_r_data_1_load_store       ), //o
    .io_out_r_data_1_df_is_ws          (cellSARA_8_io_out_r_data_1_df_is_ws         ), //o
    .io_out_r_data_1_stall             (cellSARA_8_io_out_r_data_1_stall            ), //o
    .io_out_r_data_2_data              (cellSARA_8_io_out_r_data_2_data[15:0]       ), //o
    .io_out_r_data_2_load_store        (cellSARA_8_io_out_r_data_2_load_store       ), //o
    .io_out_r_data_2_df_is_ws          (cellSARA_8_io_out_r_data_2_df_is_ws         ), //o
    .io_out_r_data_2_stall             (cellSARA_8_io_out_r_data_2_stall            ), //o
    .io_out_r_data_3_data              (cellSARA_8_io_out_r_data_3_data[15:0]       ), //o
    .io_out_r_data_3_load_store        (cellSARA_8_io_out_r_data_3_load_store       ), //o
    .io_out_r_data_3_df_is_ws          (cellSARA_8_io_out_r_data_3_df_is_ws         ), //o
    .io_out_r_data_3_stall             (cellSARA_8_io_out_r_data_3_stall            ), //o
    .io_out_r_bypass_0_0_data          (cellSARA_8_io_out_r_bypass_0_0_data[15:0]   ), //o
    .io_out_r_bypass_0_0_load_store    (cellSARA_8_io_out_r_bypass_0_0_load_store   ), //o
    .io_out_r_bypass_0_0_df_is_ws      (cellSARA_8_io_out_r_bypass_0_0_df_is_ws     ), //o
    .io_out_r_bypass_0_0_stall         (cellSARA_8_io_out_r_bypass_0_0_stall        ), //o
    .io_out_r_bypass_0_1_data          (cellSARA_8_io_out_r_bypass_0_1_data[15:0]   ), //o
    .io_out_r_bypass_0_1_load_store    (cellSARA_8_io_out_r_bypass_0_1_load_store   ), //o
    .io_out_r_bypass_0_1_df_is_ws      (cellSARA_8_io_out_r_bypass_0_1_df_is_ws     ), //o
    .io_out_r_bypass_0_1_stall         (cellSARA_8_io_out_r_bypass_0_1_stall        ), //o
    .io_out_r_bypass_0_2_data          (cellSARA_8_io_out_r_bypass_0_2_data[15:0]   ), //o
    .io_out_r_bypass_0_2_load_store    (cellSARA_8_io_out_r_bypass_0_2_load_store   ), //o
    .io_out_r_bypass_0_2_df_is_ws      (cellSARA_8_io_out_r_bypass_0_2_df_is_ws     ), //o
    .io_out_r_bypass_0_2_stall         (cellSARA_8_io_out_r_bypass_0_2_stall        ), //o
    .io_out_r_bypass_0_3_data          (cellSARA_8_io_out_r_bypass_0_3_data[15:0]   ), //o
    .io_out_r_bypass_0_3_load_store    (cellSARA_8_io_out_r_bypass_0_3_load_store   ), //o
    .io_out_r_bypass_0_3_df_is_ws      (cellSARA_8_io_out_r_bypass_0_3_df_is_ws     ), //o
    .io_out_r_bypass_0_3_stall         (cellSARA_8_io_out_r_bypass_0_3_stall        ), //o
    .io_out_r_bypass_1_0_data          (cellSARA_8_io_out_r_bypass_1_0_data[15:0]   ), //o
    .io_out_r_bypass_1_0_load_store    (cellSARA_8_io_out_r_bypass_1_0_load_store   ), //o
    .io_out_r_bypass_1_0_df_is_ws      (cellSARA_8_io_out_r_bypass_1_0_df_is_ws     ), //o
    .io_out_r_bypass_1_0_stall         (cellSARA_8_io_out_r_bypass_1_0_stall        ), //o
    .io_out_r_bypass_1_1_data          (cellSARA_8_io_out_r_bypass_1_1_data[15:0]   ), //o
    .io_out_r_bypass_1_1_load_store    (cellSARA_8_io_out_r_bypass_1_1_load_store   ), //o
    .io_out_r_bypass_1_1_df_is_ws      (cellSARA_8_io_out_r_bypass_1_1_df_is_ws     ), //o
    .io_out_r_bypass_1_1_stall         (cellSARA_8_io_out_r_bypass_1_1_stall        ), //o
    .io_out_r_bypass_1_2_data          (cellSARA_8_io_out_r_bypass_1_2_data[15:0]   ), //o
    .io_out_r_bypass_1_2_load_store    (cellSARA_8_io_out_r_bypass_1_2_load_store   ), //o
    .io_out_r_bypass_1_2_df_is_ws      (cellSARA_8_io_out_r_bypass_1_2_df_is_ws     ), //o
    .io_out_r_bypass_1_2_stall         (cellSARA_8_io_out_r_bypass_1_2_stall        ), //o
    .io_out_r_bypass_1_3_data          (cellSARA_8_io_out_r_bypass_1_3_data[15:0]   ), //o
    .io_out_r_bypass_1_3_load_store    (cellSARA_8_io_out_r_bypass_1_3_load_store   ), //o
    .io_out_r_bypass_1_3_df_is_ws      (cellSARA_8_io_out_r_bypass_1_3_df_is_ws     ), //o
    .io_out_r_bypass_1_3_stall         (cellSARA_8_io_out_r_bypass_1_3_stall        ), //o
    .io_out_r_input_from_bypass_0      (cellSARA_8_io_out_r_input_from_bypass_0     ), //o
    .io_out_r_input_from_bypass_1      (cellSARA_8_io_out_r_input_from_bypass_1     ), //o
    .io_in_c_data_0_data               (cellSARA_8_io_in_c_data_0_data[15:0]        ), //i
    .io_in_c_data_0_is_stationary      (cellSARA_8_io_in_c_data_0_is_stationary     ), //i
    .io_in_c_data_1_data               (cellSARA_8_io_in_c_data_1_data[15:0]        ), //i
    .io_in_c_data_1_is_stationary      (cellSARA_8_io_in_c_data_1_is_stationary     ), //i
    .io_in_c_data_2_data               (cellSARA_8_io_in_c_data_2_data[15:0]        ), //i
    .io_in_c_data_2_is_stationary      (cellSARA_8_io_in_c_data_2_is_stationary     ), //i
    .io_in_c_data_3_data               (cellSARA_8_io_in_c_data_3_data[15:0]        ), //i
    .io_in_c_data_3_is_stationary      (cellSARA_8_io_in_c_data_3_is_stationary     ), //i
    .io_in_c_bypass_0_0_data           (cellSARA_8_io_in_c_bypass_0_0_data[15:0]    ), //i
    .io_in_c_bypass_0_0_is_stationary  (cellSARA_8_io_in_c_bypass_0_0_is_stationary ), //i
    .io_in_c_bypass_0_1_data           (cellSARA_8_io_in_c_bypass_0_1_data[15:0]    ), //i
    .io_in_c_bypass_0_1_is_stationary  (cellSARA_8_io_in_c_bypass_0_1_is_stationary ), //i
    .io_in_c_bypass_0_2_data           (cellSARA_8_io_in_c_bypass_0_2_data[15:0]    ), //i
    .io_in_c_bypass_0_2_is_stationary  (cellSARA_8_io_in_c_bypass_0_2_is_stationary ), //i
    .io_in_c_bypass_0_3_data           (cellSARA_8_io_in_c_bypass_0_3_data[15:0]    ), //i
    .io_in_c_bypass_0_3_is_stationary  (cellSARA_8_io_in_c_bypass_0_3_is_stationary ), //i
    .io_in_c_bypass_1_0_data           (cellSARA_8_io_in_c_bypass_1_0_data[15:0]    ), //i
    .io_in_c_bypass_1_0_is_stationary  (cellSARA_8_io_in_c_bypass_1_0_is_stationary ), //i
    .io_in_c_bypass_1_1_data           (cellSARA_8_io_in_c_bypass_1_1_data[15:0]    ), //i
    .io_in_c_bypass_1_1_is_stationary  (cellSARA_8_io_in_c_bypass_1_1_is_stationary ), //i
    .io_in_c_bypass_1_2_data           (cellSARA_8_io_in_c_bypass_1_2_data[15:0]    ), //i
    .io_in_c_bypass_1_2_is_stationary  (cellSARA_8_io_in_c_bypass_1_2_is_stationary ), //i
    .io_in_c_bypass_1_3_data           (cellSARA_8_io_in_c_bypass_1_3_data[15:0]    ), //i
    .io_in_c_bypass_1_3_is_stationary  (cellSARA_8_io_in_c_bypass_1_3_is_stationary ), //i
    .io_in_c_input_from_bypass_0       (cellSARA_8_io_in_c_input_from_bypass_0      ), //i
    .io_in_c_input_from_bypass_1       (cellSARA_8_io_in_c_input_from_bypass_1      ), //i
    .io_out_c_data_0_data              (cellSARA_8_io_out_c_data_0_data[15:0]       ), //o
    .io_out_c_data_0_is_stationary     (cellSARA_8_io_out_c_data_0_is_stationary    ), //o
    .io_out_c_data_1_data              (cellSARA_8_io_out_c_data_1_data[15:0]       ), //o
    .io_out_c_data_1_is_stationary     (cellSARA_8_io_out_c_data_1_is_stationary    ), //o
    .io_out_c_data_2_data              (cellSARA_8_io_out_c_data_2_data[15:0]       ), //o
    .io_out_c_data_2_is_stationary     (cellSARA_8_io_out_c_data_2_is_stationary    ), //o
    .io_out_c_data_3_data              (cellSARA_8_io_out_c_data_3_data[15:0]       ), //o
    .io_out_c_data_3_is_stationary     (cellSARA_8_io_out_c_data_3_is_stationary    ), //o
    .io_out_c_bypass_0_0_data          (cellSARA_8_io_out_c_bypass_0_0_data[15:0]   ), //o
    .io_out_c_bypass_0_0_is_stationary (cellSARA_8_io_out_c_bypass_0_0_is_stationary), //o
    .io_out_c_bypass_0_1_data          (cellSARA_8_io_out_c_bypass_0_1_data[15:0]   ), //o
    .io_out_c_bypass_0_1_is_stationary (cellSARA_8_io_out_c_bypass_0_1_is_stationary), //o
    .io_out_c_bypass_0_2_data          (cellSARA_8_io_out_c_bypass_0_2_data[15:0]   ), //o
    .io_out_c_bypass_0_2_is_stationary (cellSARA_8_io_out_c_bypass_0_2_is_stationary), //o
    .io_out_c_bypass_0_3_data          (cellSARA_8_io_out_c_bypass_0_3_data[15:0]   ), //o
    .io_out_c_bypass_0_3_is_stationary (cellSARA_8_io_out_c_bypass_0_3_is_stationary), //o
    .io_out_c_bypass_1_0_data          (cellSARA_8_io_out_c_bypass_1_0_data[15:0]   ), //o
    .io_out_c_bypass_1_0_is_stationary (cellSARA_8_io_out_c_bypass_1_0_is_stationary), //o
    .io_out_c_bypass_1_1_data          (cellSARA_8_io_out_c_bypass_1_1_data[15:0]   ), //o
    .io_out_c_bypass_1_1_is_stationary (cellSARA_8_io_out_c_bypass_1_1_is_stationary), //o
    .io_out_c_bypass_1_2_data          (cellSARA_8_io_out_c_bypass_1_2_data[15:0]   ), //o
    .io_out_c_bypass_1_2_is_stationary (cellSARA_8_io_out_c_bypass_1_2_is_stationary), //o
    .io_out_c_bypass_1_3_data          (cellSARA_8_io_out_c_bypass_1_3_data[15:0]   ), //o
    .io_out_c_bypass_1_3_is_stationary (cellSARA_8_io_out_c_bypass_1_3_is_stationary), //o
    .io_out_c_input_from_bypass_0      (cellSARA_8_io_out_c_input_from_bypass_0     ), //o
    .io_out_c_input_from_bypass_1      (cellSARA_8_io_out_c_input_from_bypass_1     ), //o
    .clk                               (clk                                         ), //i
    .reset                             (reset                                       )  //i
  );
  CellSARA_2 cellSARA_9 (
    .io_in_r_data_0_data               (cellSARA_9_io_in_r_data_0_data[15:0]        ), //i
    .io_in_r_data_0_load_store         (cellSARA_9_io_in_r_data_0_load_store        ), //i
    .io_in_r_data_0_df_is_ws           (cellSARA_9_io_in_r_data_0_df_is_ws          ), //i
    .io_in_r_data_0_stall              (cellSARA_9_io_in_r_data_0_stall             ), //i
    .io_in_r_data_1_data               (cellSARA_9_io_in_r_data_1_data[15:0]        ), //i
    .io_in_r_data_1_load_store         (cellSARA_9_io_in_r_data_1_load_store        ), //i
    .io_in_r_data_1_df_is_ws           (cellSARA_9_io_in_r_data_1_df_is_ws          ), //i
    .io_in_r_data_1_stall              (cellSARA_9_io_in_r_data_1_stall             ), //i
    .io_in_r_data_2_data               (cellSARA_9_io_in_r_data_2_data[15:0]        ), //i
    .io_in_r_data_2_load_store         (cellSARA_9_io_in_r_data_2_load_store        ), //i
    .io_in_r_data_2_df_is_ws           (cellSARA_9_io_in_r_data_2_df_is_ws          ), //i
    .io_in_r_data_2_stall              (cellSARA_9_io_in_r_data_2_stall             ), //i
    .io_in_r_data_3_data               (cellSARA_9_io_in_r_data_3_data[15:0]        ), //i
    .io_in_r_data_3_load_store         (cellSARA_9_io_in_r_data_3_load_store        ), //i
    .io_in_r_data_3_df_is_ws           (cellSARA_9_io_in_r_data_3_df_is_ws          ), //i
    .io_in_r_data_3_stall              (cellSARA_9_io_in_r_data_3_stall             ), //i
    .io_in_r_bypass_0_0_data           (cellSARA_9_io_in_r_bypass_0_0_data[15:0]    ), //i
    .io_in_r_bypass_0_0_load_store     (cellSARA_9_io_in_r_bypass_0_0_load_store    ), //i
    .io_in_r_bypass_0_0_df_is_ws       (cellSARA_9_io_in_r_bypass_0_0_df_is_ws      ), //i
    .io_in_r_bypass_0_0_stall          (cellSARA_9_io_in_r_bypass_0_0_stall         ), //i
    .io_in_r_bypass_0_1_data           (cellSARA_9_io_in_r_bypass_0_1_data[15:0]    ), //i
    .io_in_r_bypass_0_1_load_store     (cellSARA_9_io_in_r_bypass_0_1_load_store    ), //i
    .io_in_r_bypass_0_1_df_is_ws       (cellSARA_9_io_in_r_bypass_0_1_df_is_ws      ), //i
    .io_in_r_bypass_0_1_stall          (cellSARA_9_io_in_r_bypass_0_1_stall         ), //i
    .io_in_r_bypass_0_2_data           (cellSARA_9_io_in_r_bypass_0_2_data[15:0]    ), //i
    .io_in_r_bypass_0_2_load_store     (cellSARA_9_io_in_r_bypass_0_2_load_store    ), //i
    .io_in_r_bypass_0_2_df_is_ws       (cellSARA_9_io_in_r_bypass_0_2_df_is_ws      ), //i
    .io_in_r_bypass_0_2_stall          (cellSARA_9_io_in_r_bypass_0_2_stall         ), //i
    .io_in_r_bypass_0_3_data           (cellSARA_9_io_in_r_bypass_0_3_data[15:0]    ), //i
    .io_in_r_bypass_0_3_load_store     (cellSARA_9_io_in_r_bypass_0_3_load_store    ), //i
    .io_in_r_bypass_0_3_df_is_ws       (cellSARA_9_io_in_r_bypass_0_3_df_is_ws      ), //i
    .io_in_r_bypass_0_3_stall          (cellSARA_9_io_in_r_bypass_0_3_stall         ), //i
    .io_in_r_bypass_1_0_data           (cellSARA_9_io_in_r_bypass_1_0_data[15:0]    ), //i
    .io_in_r_bypass_1_0_load_store     (cellSARA_9_io_in_r_bypass_1_0_load_store    ), //i
    .io_in_r_bypass_1_0_df_is_ws       (cellSARA_9_io_in_r_bypass_1_0_df_is_ws      ), //i
    .io_in_r_bypass_1_0_stall          (cellSARA_9_io_in_r_bypass_1_0_stall         ), //i
    .io_in_r_bypass_1_1_data           (cellSARA_9_io_in_r_bypass_1_1_data[15:0]    ), //i
    .io_in_r_bypass_1_1_load_store     (cellSARA_9_io_in_r_bypass_1_1_load_store    ), //i
    .io_in_r_bypass_1_1_df_is_ws       (cellSARA_9_io_in_r_bypass_1_1_df_is_ws      ), //i
    .io_in_r_bypass_1_1_stall          (cellSARA_9_io_in_r_bypass_1_1_stall         ), //i
    .io_in_r_bypass_1_2_data           (cellSARA_9_io_in_r_bypass_1_2_data[15:0]    ), //i
    .io_in_r_bypass_1_2_load_store     (cellSARA_9_io_in_r_bypass_1_2_load_store    ), //i
    .io_in_r_bypass_1_2_df_is_ws       (cellSARA_9_io_in_r_bypass_1_2_df_is_ws      ), //i
    .io_in_r_bypass_1_2_stall          (cellSARA_9_io_in_r_bypass_1_2_stall         ), //i
    .io_in_r_bypass_1_3_data           (cellSARA_9_io_in_r_bypass_1_3_data[15:0]    ), //i
    .io_in_r_bypass_1_3_load_store     (cellSARA_9_io_in_r_bypass_1_3_load_store    ), //i
    .io_in_r_bypass_1_3_df_is_ws       (cellSARA_9_io_in_r_bypass_1_3_df_is_ws      ), //i
    .io_in_r_bypass_1_3_stall          (cellSARA_9_io_in_r_bypass_1_3_stall         ), //i
    .io_in_r_input_from_bypass_0       (cellSARA_9_io_in_r_input_from_bypass_0      ), //i
    .io_in_r_input_from_bypass_1       (cellSARA_9_io_in_r_input_from_bypass_1      ), //i
    .io_out_r_data_0_data              (cellSARA_9_io_out_r_data_0_data[15:0]       ), //o
    .io_out_r_data_0_load_store        (cellSARA_9_io_out_r_data_0_load_store       ), //o
    .io_out_r_data_0_df_is_ws          (cellSARA_9_io_out_r_data_0_df_is_ws         ), //o
    .io_out_r_data_0_stall             (cellSARA_9_io_out_r_data_0_stall            ), //o
    .io_out_r_data_1_data              (cellSARA_9_io_out_r_data_1_data[15:0]       ), //o
    .io_out_r_data_1_load_store        (cellSARA_9_io_out_r_data_1_load_store       ), //o
    .io_out_r_data_1_df_is_ws          (cellSARA_9_io_out_r_data_1_df_is_ws         ), //o
    .io_out_r_data_1_stall             (cellSARA_9_io_out_r_data_1_stall            ), //o
    .io_out_r_data_2_data              (cellSARA_9_io_out_r_data_2_data[15:0]       ), //o
    .io_out_r_data_2_load_store        (cellSARA_9_io_out_r_data_2_load_store       ), //o
    .io_out_r_data_2_df_is_ws          (cellSARA_9_io_out_r_data_2_df_is_ws         ), //o
    .io_out_r_data_2_stall             (cellSARA_9_io_out_r_data_2_stall            ), //o
    .io_out_r_data_3_data              (cellSARA_9_io_out_r_data_3_data[15:0]       ), //o
    .io_out_r_data_3_load_store        (cellSARA_9_io_out_r_data_3_load_store       ), //o
    .io_out_r_data_3_df_is_ws          (cellSARA_9_io_out_r_data_3_df_is_ws         ), //o
    .io_out_r_data_3_stall             (cellSARA_9_io_out_r_data_3_stall            ), //o
    .io_out_r_bypass_0_0_data          (cellSARA_9_io_out_r_bypass_0_0_data[15:0]   ), //o
    .io_out_r_bypass_0_0_load_store    (cellSARA_9_io_out_r_bypass_0_0_load_store   ), //o
    .io_out_r_bypass_0_0_df_is_ws      (cellSARA_9_io_out_r_bypass_0_0_df_is_ws     ), //o
    .io_out_r_bypass_0_0_stall         (cellSARA_9_io_out_r_bypass_0_0_stall        ), //o
    .io_out_r_bypass_0_1_data          (cellSARA_9_io_out_r_bypass_0_1_data[15:0]   ), //o
    .io_out_r_bypass_0_1_load_store    (cellSARA_9_io_out_r_bypass_0_1_load_store   ), //o
    .io_out_r_bypass_0_1_df_is_ws      (cellSARA_9_io_out_r_bypass_0_1_df_is_ws     ), //o
    .io_out_r_bypass_0_1_stall         (cellSARA_9_io_out_r_bypass_0_1_stall        ), //o
    .io_out_r_bypass_0_2_data          (cellSARA_9_io_out_r_bypass_0_2_data[15:0]   ), //o
    .io_out_r_bypass_0_2_load_store    (cellSARA_9_io_out_r_bypass_0_2_load_store   ), //o
    .io_out_r_bypass_0_2_df_is_ws      (cellSARA_9_io_out_r_bypass_0_2_df_is_ws     ), //o
    .io_out_r_bypass_0_2_stall         (cellSARA_9_io_out_r_bypass_0_2_stall        ), //o
    .io_out_r_bypass_0_3_data          (cellSARA_9_io_out_r_bypass_0_3_data[15:0]   ), //o
    .io_out_r_bypass_0_3_load_store    (cellSARA_9_io_out_r_bypass_0_3_load_store   ), //o
    .io_out_r_bypass_0_3_df_is_ws      (cellSARA_9_io_out_r_bypass_0_3_df_is_ws     ), //o
    .io_out_r_bypass_0_3_stall         (cellSARA_9_io_out_r_bypass_0_3_stall        ), //o
    .io_out_r_bypass_1_0_data          (cellSARA_9_io_out_r_bypass_1_0_data[15:0]   ), //o
    .io_out_r_bypass_1_0_load_store    (cellSARA_9_io_out_r_bypass_1_0_load_store   ), //o
    .io_out_r_bypass_1_0_df_is_ws      (cellSARA_9_io_out_r_bypass_1_0_df_is_ws     ), //o
    .io_out_r_bypass_1_0_stall         (cellSARA_9_io_out_r_bypass_1_0_stall        ), //o
    .io_out_r_bypass_1_1_data          (cellSARA_9_io_out_r_bypass_1_1_data[15:0]   ), //o
    .io_out_r_bypass_1_1_load_store    (cellSARA_9_io_out_r_bypass_1_1_load_store   ), //o
    .io_out_r_bypass_1_1_df_is_ws      (cellSARA_9_io_out_r_bypass_1_1_df_is_ws     ), //o
    .io_out_r_bypass_1_1_stall         (cellSARA_9_io_out_r_bypass_1_1_stall        ), //o
    .io_out_r_bypass_1_2_data          (cellSARA_9_io_out_r_bypass_1_2_data[15:0]   ), //o
    .io_out_r_bypass_1_2_load_store    (cellSARA_9_io_out_r_bypass_1_2_load_store   ), //o
    .io_out_r_bypass_1_2_df_is_ws      (cellSARA_9_io_out_r_bypass_1_2_df_is_ws     ), //o
    .io_out_r_bypass_1_2_stall         (cellSARA_9_io_out_r_bypass_1_2_stall        ), //o
    .io_out_r_bypass_1_3_data          (cellSARA_9_io_out_r_bypass_1_3_data[15:0]   ), //o
    .io_out_r_bypass_1_3_load_store    (cellSARA_9_io_out_r_bypass_1_3_load_store   ), //o
    .io_out_r_bypass_1_3_df_is_ws      (cellSARA_9_io_out_r_bypass_1_3_df_is_ws     ), //o
    .io_out_r_bypass_1_3_stall         (cellSARA_9_io_out_r_bypass_1_3_stall        ), //o
    .io_out_r_input_from_bypass_0      (cellSARA_9_io_out_r_input_from_bypass_0     ), //o
    .io_out_r_input_from_bypass_1      (cellSARA_9_io_out_r_input_from_bypass_1     ), //o
    .io_in_c_data_0_data               (cellSARA_9_io_in_c_data_0_data[15:0]        ), //i
    .io_in_c_data_0_is_stationary      (cellSARA_9_io_in_c_data_0_is_stationary     ), //i
    .io_in_c_data_1_data               (cellSARA_9_io_in_c_data_1_data[15:0]        ), //i
    .io_in_c_data_1_is_stationary      (cellSARA_9_io_in_c_data_1_is_stationary     ), //i
    .io_in_c_data_2_data               (cellSARA_9_io_in_c_data_2_data[15:0]        ), //i
    .io_in_c_data_2_is_stationary      (cellSARA_9_io_in_c_data_2_is_stationary     ), //i
    .io_in_c_data_3_data               (cellSARA_9_io_in_c_data_3_data[15:0]        ), //i
    .io_in_c_data_3_is_stationary      (cellSARA_9_io_in_c_data_3_is_stationary     ), //i
    .io_in_c_bypass_0_0_data           (cellSARA_9_io_in_c_bypass_0_0_data[15:0]    ), //i
    .io_in_c_bypass_0_0_is_stationary  (cellSARA_9_io_in_c_bypass_0_0_is_stationary ), //i
    .io_in_c_bypass_0_1_data           (cellSARA_9_io_in_c_bypass_0_1_data[15:0]    ), //i
    .io_in_c_bypass_0_1_is_stationary  (cellSARA_9_io_in_c_bypass_0_1_is_stationary ), //i
    .io_in_c_bypass_0_2_data           (cellSARA_9_io_in_c_bypass_0_2_data[15:0]    ), //i
    .io_in_c_bypass_0_2_is_stationary  (cellSARA_9_io_in_c_bypass_0_2_is_stationary ), //i
    .io_in_c_bypass_0_3_data           (cellSARA_9_io_in_c_bypass_0_3_data[15:0]    ), //i
    .io_in_c_bypass_0_3_is_stationary  (cellSARA_9_io_in_c_bypass_0_3_is_stationary ), //i
    .io_in_c_bypass_1_0_data           (cellSARA_9_io_in_c_bypass_1_0_data[15:0]    ), //i
    .io_in_c_bypass_1_0_is_stationary  (cellSARA_9_io_in_c_bypass_1_0_is_stationary ), //i
    .io_in_c_bypass_1_1_data           (cellSARA_9_io_in_c_bypass_1_1_data[15:0]    ), //i
    .io_in_c_bypass_1_1_is_stationary  (cellSARA_9_io_in_c_bypass_1_1_is_stationary ), //i
    .io_in_c_bypass_1_2_data           (cellSARA_9_io_in_c_bypass_1_2_data[15:0]    ), //i
    .io_in_c_bypass_1_2_is_stationary  (cellSARA_9_io_in_c_bypass_1_2_is_stationary ), //i
    .io_in_c_bypass_1_3_data           (cellSARA_9_io_in_c_bypass_1_3_data[15:0]    ), //i
    .io_in_c_bypass_1_3_is_stationary  (cellSARA_9_io_in_c_bypass_1_3_is_stationary ), //i
    .io_in_c_input_from_bypass_0       (cellSARA_9_io_in_c_input_from_bypass_0      ), //i
    .io_in_c_input_from_bypass_1       (cellSARA_9_io_in_c_input_from_bypass_1      ), //i
    .io_out_c_data_0_data              (cellSARA_9_io_out_c_data_0_data[15:0]       ), //o
    .io_out_c_data_0_is_stationary     (cellSARA_9_io_out_c_data_0_is_stationary    ), //o
    .io_out_c_data_1_data              (cellSARA_9_io_out_c_data_1_data[15:0]       ), //o
    .io_out_c_data_1_is_stationary     (cellSARA_9_io_out_c_data_1_is_stationary    ), //o
    .io_out_c_data_2_data              (cellSARA_9_io_out_c_data_2_data[15:0]       ), //o
    .io_out_c_data_2_is_stationary     (cellSARA_9_io_out_c_data_2_is_stationary    ), //o
    .io_out_c_data_3_data              (cellSARA_9_io_out_c_data_3_data[15:0]       ), //o
    .io_out_c_data_3_is_stationary     (cellSARA_9_io_out_c_data_3_is_stationary    ), //o
    .io_out_c_bypass_0_0_data          (cellSARA_9_io_out_c_bypass_0_0_data[15:0]   ), //o
    .io_out_c_bypass_0_0_is_stationary (cellSARA_9_io_out_c_bypass_0_0_is_stationary), //o
    .io_out_c_bypass_0_1_data          (cellSARA_9_io_out_c_bypass_0_1_data[15:0]   ), //o
    .io_out_c_bypass_0_1_is_stationary (cellSARA_9_io_out_c_bypass_0_1_is_stationary), //o
    .io_out_c_bypass_0_2_data          (cellSARA_9_io_out_c_bypass_0_2_data[15:0]   ), //o
    .io_out_c_bypass_0_2_is_stationary (cellSARA_9_io_out_c_bypass_0_2_is_stationary), //o
    .io_out_c_bypass_0_3_data          (cellSARA_9_io_out_c_bypass_0_3_data[15:0]   ), //o
    .io_out_c_bypass_0_3_is_stationary (cellSARA_9_io_out_c_bypass_0_3_is_stationary), //o
    .io_out_c_bypass_1_0_data          (cellSARA_9_io_out_c_bypass_1_0_data[15:0]   ), //o
    .io_out_c_bypass_1_0_is_stationary (cellSARA_9_io_out_c_bypass_1_0_is_stationary), //o
    .io_out_c_bypass_1_1_data          (cellSARA_9_io_out_c_bypass_1_1_data[15:0]   ), //o
    .io_out_c_bypass_1_1_is_stationary (cellSARA_9_io_out_c_bypass_1_1_is_stationary), //o
    .io_out_c_bypass_1_2_data          (cellSARA_9_io_out_c_bypass_1_2_data[15:0]   ), //o
    .io_out_c_bypass_1_2_is_stationary (cellSARA_9_io_out_c_bypass_1_2_is_stationary), //o
    .io_out_c_bypass_1_3_data          (cellSARA_9_io_out_c_bypass_1_3_data[15:0]   ), //o
    .io_out_c_bypass_1_3_is_stationary (cellSARA_9_io_out_c_bypass_1_3_is_stationary), //o
    .io_out_c_input_from_bypass_0      (cellSARA_9_io_out_c_input_from_bypass_0     ), //o
    .io_out_c_input_from_bypass_1      (cellSARA_9_io_out_c_input_from_bypass_1     ), //o
    .clk                               (clk                                         ), //i
    .reset                             (reset                                       )  //i
  );
  CellSARA_1 cellSARA_10 (
    .io_in_r_data_0_data               (cellSARA_10_io_in_r_data_0_data[15:0]        ), //i
    .io_in_r_data_0_load_store         (cellSARA_10_io_in_r_data_0_load_store        ), //i
    .io_in_r_data_0_df_is_ws           (cellSARA_10_io_in_r_data_0_df_is_ws          ), //i
    .io_in_r_data_0_stall              (cellSARA_10_io_in_r_data_0_stall             ), //i
    .io_in_r_data_1_data               (cellSARA_10_io_in_r_data_1_data[15:0]        ), //i
    .io_in_r_data_1_load_store         (cellSARA_10_io_in_r_data_1_load_store        ), //i
    .io_in_r_data_1_df_is_ws           (cellSARA_10_io_in_r_data_1_df_is_ws          ), //i
    .io_in_r_data_1_stall              (cellSARA_10_io_in_r_data_1_stall             ), //i
    .io_in_r_data_2_data               (cellSARA_10_io_in_r_data_2_data[15:0]        ), //i
    .io_in_r_data_2_load_store         (cellSARA_10_io_in_r_data_2_load_store        ), //i
    .io_in_r_data_2_df_is_ws           (cellSARA_10_io_in_r_data_2_df_is_ws          ), //i
    .io_in_r_data_2_stall              (cellSARA_10_io_in_r_data_2_stall             ), //i
    .io_in_r_data_3_data               (cellSARA_10_io_in_r_data_3_data[15:0]        ), //i
    .io_in_r_data_3_load_store         (cellSARA_10_io_in_r_data_3_load_store        ), //i
    .io_in_r_data_3_df_is_ws           (cellSARA_10_io_in_r_data_3_df_is_ws          ), //i
    .io_in_r_data_3_stall              (cellSARA_10_io_in_r_data_3_stall             ), //i
    .io_in_r_bypass_0_0_data           (cellSARA_10_io_in_r_bypass_0_0_data[15:0]    ), //i
    .io_in_r_bypass_0_0_load_store     (cellSARA_10_io_in_r_bypass_0_0_load_store    ), //i
    .io_in_r_bypass_0_0_df_is_ws       (cellSARA_10_io_in_r_bypass_0_0_df_is_ws      ), //i
    .io_in_r_bypass_0_0_stall          (cellSARA_10_io_in_r_bypass_0_0_stall         ), //i
    .io_in_r_bypass_0_1_data           (cellSARA_10_io_in_r_bypass_0_1_data[15:0]    ), //i
    .io_in_r_bypass_0_1_load_store     (cellSARA_10_io_in_r_bypass_0_1_load_store    ), //i
    .io_in_r_bypass_0_1_df_is_ws       (cellSARA_10_io_in_r_bypass_0_1_df_is_ws      ), //i
    .io_in_r_bypass_0_1_stall          (cellSARA_10_io_in_r_bypass_0_1_stall         ), //i
    .io_in_r_bypass_0_2_data           (cellSARA_10_io_in_r_bypass_0_2_data[15:0]    ), //i
    .io_in_r_bypass_0_2_load_store     (cellSARA_10_io_in_r_bypass_0_2_load_store    ), //i
    .io_in_r_bypass_0_2_df_is_ws       (cellSARA_10_io_in_r_bypass_0_2_df_is_ws      ), //i
    .io_in_r_bypass_0_2_stall          (cellSARA_10_io_in_r_bypass_0_2_stall         ), //i
    .io_in_r_bypass_0_3_data           (cellSARA_10_io_in_r_bypass_0_3_data[15:0]    ), //i
    .io_in_r_bypass_0_3_load_store     (cellSARA_10_io_in_r_bypass_0_3_load_store    ), //i
    .io_in_r_bypass_0_3_df_is_ws       (cellSARA_10_io_in_r_bypass_0_3_df_is_ws      ), //i
    .io_in_r_bypass_0_3_stall          (cellSARA_10_io_in_r_bypass_0_3_stall         ), //i
    .io_in_r_bypass_1_0_data           (cellSARA_10_io_in_r_bypass_1_0_data[15:0]    ), //i
    .io_in_r_bypass_1_0_load_store     (cellSARA_10_io_in_r_bypass_1_0_load_store    ), //i
    .io_in_r_bypass_1_0_df_is_ws       (cellSARA_10_io_in_r_bypass_1_0_df_is_ws      ), //i
    .io_in_r_bypass_1_0_stall          (cellSARA_10_io_in_r_bypass_1_0_stall         ), //i
    .io_in_r_bypass_1_1_data           (cellSARA_10_io_in_r_bypass_1_1_data[15:0]    ), //i
    .io_in_r_bypass_1_1_load_store     (cellSARA_10_io_in_r_bypass_1_1_load_store    ), //i
    .io_in_r_bypass_1_1_df_is_ws       (cellSARA_10_io_in_r_bypass_1_1_df_is_ws      ), //i
    .io_in_r_bypass_1_1_stall          (cellSARA_10_io_in_r_bypass_1_1_stall         ), //i
    .io_in_r_bypass_1_2_data           (cellSARA_10_io_in_r_bypass_1_2_data[15:0]    ), //i
    .io_in_r_bypass_1_2_load_store     (cellSARA_10_io_in_r_bypass_1_2_load_store    ), //i
    .io_in_r_bypass_1_2_df_is_ws       (cellSARA_10_io_in_r_bypass_1_2_df_is_ws      ), //i
    .io_in_r_bypass_1_2_stall          (cellSARA_10_io_in_r_bypass_1_2_stall         ), //i
    .io_in_r_bypass_1_3_data           (cellSARA_10_io_in_r_bypass_1_3_data[15:0]    ), //i
    .io_in_r_bypass_1_3_load_store     (cellSARA_10_io_in_r_bypass_1_3_load_store    ), //i
    .io_in_r_bypass_1_3_df_is_ws       (cellSARA_10_io_in_r_bypass_1_3_df_is_ws      ), //i
    .io_in_r_bypass_1_3_stall          (cellSARA_10_io_in_r_bypass_1_3_stall         ), //i
    .io_in_r_input_from_bypass_0       (cellSARA_10_io_in_r_input_from_bypass_0      ), //i
    .io_in_r_input_from_bypass_1       (cellSARA_10_io_in_r_input_from_bypass_1      ), //i
    .io_out_r_data_0_data              (cellSARA_10_io_out_r_data_0_data[15:0]       ), //o
    .io_out_r_data_0_load_store        (cellSARA_10_io_out_r_data_0_load_store       ), //o
    .io_out_r_data_0_df_is_ws          (cellSARA_10_io_out_r_data_0_df_is_ws         ), //o
    .io_out_r_data_0_stall             (cellSARA_10_io_out_r_data_0_stall            ), //o
    .io_out_r_data_1_data              (cellSARA_10_io_out_r_data_1_data[15:0]       ), //o
    .io_out_r_data_1_load_store        (cellSARA_10_io_out_r_data_1_load_store       ), //o
    .io_out_r_data_1_df_is_ws          (cellSARA_10_io_out_r_data_1_df_is_ws         ), //o
    .io_out_r_data_1_stall             (cellSARA_10_io_out_r_data_1_stall            ), //o
    .io_out_r_data_2_data              (cellSARA_10_io_out_r_data_2_data[15:0]       ), //o
    .io_out_r_data_2_load_store        (cellSARA_10_io_out_r_data_2_load_store       ), //o
    .io_out_r_data_2_df_is_ws          (cellSARA_10_io_out_r_data_2_df_is_ws         ), //o
    .io_out_r_data_2_stall             (cellSARA_10_io_out_r_data_2_stall            ), //o
    .io_out_r_data_3_data              (cellSARA_10_io_out_r_data_3_data[15:0]       ), //o
    .io_out_r_data_3_load_store        (cellSARA_10_io_out_r_data_3_load_store       ), //o
    .io_out_r_data_3_df_is_ws          (cellSARA_10_io_out_r_data_3_df_is_ws         ), //o
    .io_out_r_data_3_stall             (cellSARA_10_io_out_r_data_3_stall            ), //o
    .io_out_r_bypass_0_0_data          (cellSARA_10_io_out_r_bypass_0_0_data[15:0]   ), //o
    .io_out_r_bypass_0_0_load_store    (cellSARA_10_io_out_r_bypass_0_0_load_store   ), //o
    .io_out_r_bypass_0_0_df_is_ws      (cellSARA_10_io_out_r_bypass_0_0_df_is_ws     ), //o
    .io_out_r_bypass_0_0_stall         (cellSARA_10_io_out_r_bypass_0_0_stall        ), //o
    .io_out_r_bypass_0_1_data          (cellSARA_10_io_out_r_bypass_0_1_data[15:0]   ), //o
    .io_out_r_bypass_0_1_load_store    (cellSARA_10_io_out_r_bypass_0_1_load_store   ), //o
    .io_out_r_bypass_0_1_df_is_ws      (cellSARA_10_io_out_r_bypass_0_1_df_is_ws     ), //o
    .io_out_r_bypass_0_1_stall         (cellSARA_10_io_out_r_bypass_0_1_stall        ), //o
    .io_out_r_bypass_0_2_data          (cellSARA_10_io_out_r_bypass_0_2_data[15:0]   ), //o
    .io_out_r_bypass_0_2_load_store    (cellSARA_10_io_out_r_bypass_0_2_load_store   ), //o
    .io_out_r_bypass_0_2_df_is_ws      (cellSARA_10_io_out_r_bypass_0_2_df_is_ws     ), //o
    .io_out_r_bypass_0_2_stall         (cellSARA_10_io_out_r_bypass_0_2_stall        ), //o
    .io_out_r_bypass_0_3_data          (cellSARA_10_io_out_r_bypass_0_3_data[15:0]   ), //o
    .io_out_r_bypass_0_3_load_store    (cellSARA_10_io_out_r_bypass_0_3_load_store   ), //o
    .io_out_r_bypass_0_3_df_is_ws      (cellSARA_10_io_out_r_bypass_0_3_df_is_ws     ), //o
    .io_out_r_bypass_0_3_stall         (cellSARA_10_io_out_r_bypass_0_3_stall        ), //o
    .io_out_r_bypass_1_0_data          (cellSARA_10_io_out_r_bypass_1_0_data[15:0]   ), //o
    .io_out_r_bypass_1_0_load_store    (cellSARA_10_io_out_r_bypass_1_0_load_store   ), //o
    .io_out_r_bypass_1_0_df_is_ws      (cellSARA_10_io_out_r_bypass_1_0_df_is_ws     ), //o
    .io_out_r_bypass_1_0_stall         (cellSARA_10_io_out_r_bypass_1_0_stall        ), //o
    .io_out_r_bypass_1_1_data          (cellSARA_10_io_out_r_bypass_1_1_data[15:0]   ), //o
    .io_out_r_bypass_1_1_load_store    (cellSARA_10_io_out_r_bypass_1_1_load_store   ), //o
    .io_out_r_bypass_1_1_df_is_ws      (cellSARA_10_io_out_r_bypass_1_1_df_is_ws     ), //o
    .io_out_r_bypass_1_1_stall         (cellSARA_10_io_out_r_bypass_1_1_stall        ), //o
    .io_out_r_bypass_1_2_data          (cellSARA_10_io_out_r_bypass_1_2_data[15:0]   ), //o
    .io_out_r_bypass_1_2_load_store    (cellSARA_10_io_out_r_bypass_1_2_load_store   ), //o
    .io_out_r_bypass_1_2_df_is_ws      (cellSARA_10_io_out_r_bypass_1_2_df_is_ws     ), //o
    .io_out_r_bypass_1_2_stall         (cellSARA_10_io_out_r_bypass_1_2_stall        ), //o
    .io_out_r_bypass_1_3_data          (cellSARA_10_io_out_r_bypass_1_3_data[15:0]   ), //o
    .io_out_r_bypass_1_3_load_store    (cellSARA_10_io_out_r_bypass_1_3_load_store   ), //o
    .io_out_r_bypass_1_3_df_is_ws      (cellSARA_10_io_out_r_bypass_1_3_df_is_ws     ), //o
    .io_out_r_bypass_1_3_stall         (cellSARA_10_io_out_r_bypass_1_3_stall        ), //o
    .io_out_r_input_from_bypass_0      (cellSARA_10_io_out_r_input_from_bypass_0     ), //o
    .io_out_r_input_from_bypass_1      (cellSARA_10_io_out_r_input_from_bypass_1     ), //o
    .io_in_c_data_0_data               (cellSARA_10_io_in_c_data_0_data[15:0]        ), //i
    .io_in_c_data_0_is_stationary      (cellSARA_10_io_in_c_data_0_is_stationary     ), //i
    .io_in_c_data_1_data               (cellSARA_10_io_in_c_data_1_data[15:0]        ), //i
    .io_in_c_data_1_is_stationary      (cellSARA_10_io_in_c_data_1_is_stationary     ), //i
    .io_in_c_data_2_data               (cellSARA_10_io_in_c_data_2_data[15:0]        ), //i
    .io_in_c_data_2_is_stationary      (cellSARA_10_io_in_c_data_2_is_stationary     ), //i
    .io_in_c_data_3_data               (cellSARA_10_io_in_c_data_3_data[15:0]        ), //i
    .io_in_c_data_3_is_stationary      (cellSARA_10_io_in_c_data_3_is_stationary     ), //i
    .io_in_c_bypass_0_0_data           (cellSARA_10_io_in_c_bypass_0_0_data[15:0]    ), //i
    .io_in_c_bypass_0_0_is_stationary  (cellSARA_10_io_in_c_bypass_0_0_is_stationary ), //i
    .io_in_c_bypass_0_1_data           (cellSARA_10_io_in_c_bypass_0_1_data[15:0]    ), //i
    .io_in_c_bypass_0_1_is_stationary  (cellSARA_10_io_in_c_bypass_0_1_is_stationary ), //i
    .io_in_c_bypass_0_2_data           (cellSARA_10_io_in_c_bypass_0_2_data[15:0]    ), //i
    .io_in_c_bypass_0_2_is_stationary  (cellSARA_10_io_in_c_bypass_0_2_is_stationary ), //i
    .io_in_c_bypass_0_3_data           (cellSARA_10_io_in_c_bypass_0_3_data[15:0]    ), //i
    .io_in_c_bypass_0_3_is_stationary  (cellSARA_10_io_in_c_bypass_0_3_is_stationary ), //i
    .io_in_c_bypass_1_0_data           (cellSARA_10_io_in_c_bypass_1_0_data[15:0]    ), //i
    .io_in_c_bypass_1_0_is_stationary  (cellSARA_10_io_in_c_bypass_1_0_is_stationary ), //i
    .io_in_c_bypass_1_1_data           (cellSARA_10_io_in_c_bypass_1_1_data[15:0]    ), //i
    .io_in_c_bypass_1_1_is_stationary  (cellSARA_10_io_in_c_bypass_1_1_is_stationary ), //i
    .io_in_c_bypass_1_2_data           (cellSARA_10_io_in_c_bypass_1_2_data[15:0]    ), //i
    .io_in_c_bypass_1_2_is_stationary  (cellSARA_10_io_in_c_bypass_1_2_is_stationary ), //i
    .io_in_c_bypass_1_3_data           (cellSARA_10_io_in_c_bypass_1_3_data[15:0]    ), //i
    .io_in_c_bypass_1_3_is_stationary  (cellSARA_10_io_in_c_bypass_1_3_is_stationary ), //i
    .io_in_c_input_from_bypass_0       (cellSARA_10_io_in_c_input_from_bypass_0      ), //i
    .io_in_c_input_from_bypass_1       (cellSARA_10_io_in_c_input_from_bypass_1      ), //i
    .io_out_c_data_0_data              (cellSARA_10_io_out_c_data_0_data[15:0]       ), //o
    .io_out_c_data_0_is_stationary     (cellSARA_10_io_out_c_data_0_is_stationary    ), //o
    .io_out_c_data_1_data              (cellSARA_10_io_out_c_data_1_data[15:0]       ), //o
    .io_out_c_data_1_is_stationary     (cellSARA_10_io_out_c_data_1_is_stationary    ), //o
    .io_out_c_data_2_data              (cellSARA_10_io_out_c_data_2_data[15:0]       ), //o
    .io_out_c_data_2_is_stationary     (cellSARA_10_io_out_c_data_2_is_stationary    ), //o
    .io_out_c_data_3_data              (cellSARA_10_io_out_c_data_3_data[15:0]       ), //o
    .io_out_c_data_3_is_stationary     (cellSARA_10_io_out_c_data_3_is_stationary    ), //o
    .io_out_c_bypass_0_0_data          (cellSARA_10_io_out_c_bypass_0_0_data[15:0]   ), //o
    .io_out_c_bypass_0_0_is_stationary (cellSARA_10_io_out_c_bypass_0_0_is_stationary), //o
    .io_out_c_bypass_0_1_data          (cellSARA_10_io_out_c_bypass_0_1_data[15:0]   ), //o
    .io_out_c_bypass_0_1_is_stationary (cellSARA_10_io_out_c_bypass_0_1_is_stationary), //o
    .io_out_c_bypass_0_2_data          (cellSARA_10_io_out_c_bypass_0_2_data[15:0]   ), //o
    .io_out_c_bypass_0_2_is_stationary (cellSARA_10_io_out_c_bypass_0_2_is_stationary), //o
    .io_out_c_bypass_0_3_data          (cellSARA_10_io_out_c_bypass_0_3_data[15:0]   ), //o
    .io_out_c_bypass_0_3_is_stationary (cellSARA_10_io_out_c_bypass_0_3_is_stationary), //o
    .io_out_c_bypass_1_0_data          (cellSARA_10_io_out_c_bypass_1_0_data[15:0]   ), //o
    .io_out_c_bypass_1_0_is_stationary (cellSARA_10_io_out_c_bypass_1_0_is_stationary), //o
    .io_out_c_bypass_1_1_data          (cellSARA_10_io_out_c_bypass_1_1_data[15:0]   ), //o
    .io_out_c_bypass_1_1_is_stationary (cellSARA_10_io_out_c_bypass_1_1_is_stationary), //o
    .io_out_c_bypass_1_2_data          (cellSARA_10_io_out_c_bypass_1_2_data[15:0]   ), //o
    .io_out_c_bypass_1_2_is_stationary (cellSARA_10_io_out_c_bypass_1_2_is_stationary), //o
    .io_out_c_bypass_1_3_data          (cellSARA_10_io_out_c_bypass_1_3_data[15:0]   ), //o
    .io_out_c_bypass_1_3_is_stationary (cellSARA_10_io_out_c_bypass_1_3_is_stationary), //o
    .io_out_c_input_from_bypass_0      (cellSARA_10_io_out_c_input_from_bypass_0     ), //o
    .io_out_c_input_from_bypass_1      (cellSARA_10_io_out_c_input_from_bypass_1     ), //o
    .clk                               (clk                                          ), //i
    .reset                             (reset                                        )  //i
  );
  CellSARA cellSARA_11 (
    .io_in_r_data_0_data               (cellSARA_11_io_in_r_data_0_data[15:0]        ), //i
    .io_in_r_data_0_load_store         (cellSARA_11_io_in_r_data_0_load_store        ), //i
    .io_in_r_data_0_df_is_ws           (cellSARA_11_io_in_r_data_0_df_is_ws          ), //i
    .io_in_r_data_0_stall              (cellSARA_11_io_in_r_data_0_stall             ), //i
    .io_in_r_data_1_data               (cellSARA_11_io_in_r_data_1_data[15:0]        ), //i
    .io_in_r_data_1_load_store         (cellSARA_11_io_in_r_data_1_load_store        ), //i
    .io_in_r_data_1_df_is_ws           (cellSARA_11_io_in_r_data_1_df_is_ws          ), //i
    .io_in_r_data_1_stall              (cellSARA_11_io_in_r_data_1_stall             ), //i
    .io_in_r_data_2_data               (cellSARA_11_io_in_r_data_2_data[15:0]        ), //i
    .io_in_r_data_2_load_store         (cellSARA_11_io_in_r_data_2_load_store        ), //i
    .io_in_r_data_2_df_is_ws           (cellSARA_11_io_in_r_data_2_df_is_ws          ), //i
    .io_in_r_data_2_stall              (cellSARA_11_io_in_r_data_2_stall             ), //i
    .io_in_r_data_3_data               (cellSARA_11_io_in_r_data_3_data[15:0]        ), //i
    .io_in_r_data_3_load_store         (cellSARA_11_io_in_r_data_3_load_store        ), //i
    .io_in_r_data_3_df_is_ws           (cellSARA_11_io_in_r_data_3_df_is_ws          ), //i
    .io_in_r_data_3_stall              (cellSARA_11_io_in_r_data_3_stall             ), //i
    .io_in_r_bypass_0_0_data           (cellSARA_11_io_in_r_bypass_0_0_data[15:0]    ), //i
    .io_in_r_bypass_0_0_load_store     (cellSARA_11_io_in_r_bypass_0_0_load_store    ), //i
    .io_in_r_bypass_0_0_df_is_ws       (cellSARA_11_io_in_r_bypass_0_0_df_is_ws      ), //i
    .io_in_r_bypass_0_0_stall          (cellSARA_11_io_in_r_bypass_0_0_stall         ), //i
    .io_in_r_bypass_0_1_data           (cellSARA_11_io_in_r_bypass_0_1_data[15:0]    ), //i
    .io_in_r_bypass_0_1_load_store     (cellSARA_11_io_in_r_bypass_0_1_load_store    ), //i
    .io_in_r_bypass_0_1_df_is_ws       (cellSARA_11_io_in_r_bypass_0_1_df_is_ws      ), //i
    .io_in_r_bypass_0_1_stall          (cellSARA_11_io_in_r_bypass_0_1_stall         ), //i
    .io_in_r_bypass_0_2_data           (cellSARA_11_io_in_r_bypass_0_2_data[15:0]    ), //i
    .io_in_r_bypass_0_2_load_store     (cellSARA_11_io_in_r_bypass_0_2_load_store    ), //i
    .io_in_r_bypass_0_2_df_is_ws       (cellSARA_11_io_in_r_bypass_0_2_df_is_ws      ), //i
    .io_in_r_bypass_0_2_stall          (cellSARA_11_io_in_r_bypass_0_2_stall         ), //i
    .io_in_r_bypass_0_3_data           (cellSARA_11_io_in_r_bypass_0_3_data[15:0]    ), //i
    .io_in_r_bypass_0_3_load_store     (cellSARA_11_io_in_r_bypass_0_3_load_store    ), //i
    .io_in_r_bypass_0_3_df_is_ws       (cellSARA_11_io_in_r_bypass_0_3_df_is_ws      ), //i
    .io_in_r_bypass_0_3_stall          (cellSARA_11_io_in_r_bypass_0_3_stall         ), //i
    .io_in_r_bypass_1_0_data           (cellSARA_11_io_in_r_bypass_1_0_data[15:0]    ), //i
    .io_in_r_bypass_1_0_load_store     (cellSARA_11_io_in_r_bypass_1_0_load_store    ), //i
    .io_in_r_bypass_1_0_df_is_ws       (cellSARA_11_io_in_r_bypass_1_0_df_is_ws      ), //i
    .io_in_r_bypass_1_0_stall          (cellSARA_11_io_in_r_bypass_1_0_stall         ), //i
    .io_in_r_bypass_1_1_data           (cellSARA_11_io_in_r_bypass_1_1_data[15:0]    ), //i
    .io_in_r_bypass_1_1_load_store     (cellSARA_11_io_in_r_bypass_1_1_load_store    ), //i
    .io_in_r_bypass_1_1_df_is_ws       (cellSARA_11_io_in_r_bypass_1_1_df_is_ws      ), //i
    .io_in_r_bypass_1_1_stall          (cellSARA_11_io_in_r_bypass_1_1_stall         ), //i
    .io_in_r_bypass_1_2_data           (cellSARA_11_io_in_r_bypass_1_2_data[15:0]    ), //i
    .io_in_r_bypass_1_2_load_store     (cellSARA_11_io_in_r_bypass_1_2_load_store    ), //i
    .io_in_r_bypass_1_2_df_is_ws       (cellSARA_11_io_in_r_bypass_1_2_df_is_ws      ), //i
    .io_in_r_bypass_1_2_stall          (cellSARA_11_io_in_r_bypass_1_2_stall         ), //i
    .io_in_r_bypass_1_3_data           (cellSARA_11_io_in_r_bypass_1_3_data[15:0]    ), //i
    .io_in_r_bypass_1_3_load_store     (cellSARA_11_io_in_r_bypass_1_3_load_store    ), //i
    .io_in_r_bypass_1_3_df_is_ws       (cellSARA_11_io_in_r_bypass_1_3_df_is_ws      ), //i
    .io_in_r_bypass_1_3_stall          (cellSARA_11_io_in_r_bypass_1_3_stall         ), //i
    .io_in_r_input_from_bypass_0       (cellSARA_11_io_in_r_input_from_bypass_0      ), //i
    .io_in_r_input_from_bypass_1       (cellSARA_11_io_in_r_input_from_bypass_1      ), //i
    .io_out_r_data_0_data              (cellSARA_11_io_out_r_data_0_data[15:0]       ), //o
    .io_out_r_data_0_load_store        (cellSARA_11_io_out_r_data_0_load_store       ), //o
    .io_out_r_data_0_df_is_ws          (cellSARA_11_io_out_r_data_0_df_is_ws         ), //o
    .io_out_r_data_0_stall             (cellSARA_11_io_out_r_data_0_stall            ), //o
    .io_out_r_data_1_data              (cellSARA_11_io_out_r_data_1_data[15:0]       ), //o
    .io_out_r_data_1_load_store        (cellSARA_11_io_out_r_data_1_load_store       ), //o
    .io_out_r_data_1_df_is_ws          (cellSARA_11_io_out_r_data_1_df_is_ws         ), //o
    .io_out_r_data_1_stall             (cellSARA_11_io_out_r_data_1_stall            ), //o
    .io_out_r_data_2_data              (cellSARA_11_io_out_r_data_2_data[15:0]       ), //o
    .io_out_r_data_2_load_store        (cellSARA_11_io_out_r_data_2_load_store       ), //o
    .io_out_r_data_2_df_is_ws          (cellSARA_11_io_out_r_data_2_df_is_ws         ), //o
    .io_out_r_data_2_stall             (cellSARA_11_io_out_r_data_2_stall            ), //o
    .io_out_r_data_3_data              (cellSARA_11_io_out_r_data_3_data[15:0]       ), //o
    .io_out_r_data_3_load_store        (cellSARA_11_io_out_r_data_3_load_store       ), //o
    .io_out_r_data_3_df_is_ws          (cellSARA_11_io_out_r_data_3_df_is_ws         ), //o
    .io_out_r_data_3_stall             (cellSARA_11_io_out_r_data_3_stall            ), //o
    .io_out_r_bypass_0_0_data          (cellSARA_11_io_out_r_bypass_0_0_data[15:0]   ), //o
    .io_out_r_bypass_0_0_load_store    (cellSARA_11_io_out_r_bypass_0_0_load_store   ), //o
    .io_out_r_bypass_0_0_df_is_ws      (cellSARA_11_io_out_r_bypass_0_0_df_is_ws     ), //o
    .io_out_r_bypass_0_0_stall         (cellSARA_11_io_out_r_bypass_0_0_stall        ), //o
    .io_out_r_bypass_0_1_data          (cellSARA_11_io_out_r_bypass_0_1_data[15:0]   ), //o
    .io_out_r_bypass_0_1_load_store    (cellSARA_11_io_out_r_bypass_0_1_load_store   ), //o
    .io_out_r_bypass_0_1_df_is_ws      (cellSARA_11_io_out_r_bypass_0_1_df_is_ws     ), //o
    .io_out_r_bypass_0_1_stall         (cellSARA_11_io_out_r_bypass_0_1_stall        ), //o
    .io_out_r_bypass_0_2_data          (cellSARA_11_io_out_r_bypass_0_2_data[15:0]   ), //o
    .io_out_r_bypass_0_2_load_store    (cellSARA_11_io_out_r_bypass_0_2_load_store   ), //o
    .io_out_r_bypass_0_2_df_is_ws      (cellSARA_11_io_out_r_bypass_0_2_df_is_ws     ), //o
    .io_out_r_bypass_0_2_stall         (cellSARA_11_io_out_r_bypass_0_2_stall        ), //o
    .io_out_r_bypass_0_3_data          (cellSARA_11_io_out_r_bypass_0_3_data[15:0]   ), //o
    .io_out_r_bypass_0_3_load_store    (cellSARA_11_io_out_r_bypass_0_3_load_store   ), //o
    .io_out_r_bypass_0_3_df_is_ws      (cellSARA_11_io_out_r_bypass_0_3_df_is_ws     ), //o
    .io_out_r_bypass_0_3_stall         (cellSARA_11_io_out_r_bypass_0_3_stall        ), //o
    .io_out_r_bypass_1_0_data          (cellSARA_11_io_out_r_bypass_1_0_data[15:0]   ), //o
    .io_out_r_bypass_1_0_load_store    (cellSARA_11_io_out_r_bypass_1_0_load_store   ), //o
    .io_out_r_bypass_1_0_df_is_ws      (cellSARA_11_io_out_r_bypass_1_0_df_is_ws     ), //o
    .io_out_r_bypass_1_0_stall         (cellSARA_11_io_out_r_bypass_1_0_stall        ), //o
    .io_out_r_bypass_1_1_data          (cellSARA_11_io_out_r_bypass_1_1_data[15:0]   ), //o
    .io_out_r_bypass_1_1_load_store    (cellSARA_11_io_out_r_bypass_1_1_load_store   ), //o
    .io_out_r_bypass_1_1_df_is_ws      (cellSARA_11_io_out_r_bypass_1_1_df_is_ws     ), //o
    .io_out_r_bypass_1_1_stall         (cellSARA_11_io_out_r_bypass_1_1_stall        ), //o
    .io_out_r_bypass_1_2_data          (cellSARA_11_io_out_r_bypass_1_2_data[15:0]   ), //o
    .io_out_r_bypass_1_2_load_store    (cellSARA_11_io_out_r_bypass_1_2_load_store   ), //o
    .io_out_r_bypass_1_2_df_is_ws      (cellSARA_11_io_out_r_bypass_1_2_df_is_ws     ), //o
    .io_out_r_bypass_1_2_stall         (cellSARA_11_io_out_r_bypass_1_2_stall        ), //o
    .io_out_r_bypass_1_3_data          (cellSARA_11_io_out_r_bypass_1_3_data[15:0]   ), //o
    .io_out_r_bypass_1_3_load_store    (cellSARA_11_io_out_r_bypass_1_3_load_store   ), //o
    .io_out_r_bypass_1_3_df_is_ws      (cellSARA_11_io_out_r_bypass_1_3_df_is_ws     ), //o
    .io_out_r_bypass_1_3_stall         (cellSARA_11_io_out_r_bypass_1_3_stall        ), //o
    .io_out_r_input_from_bypass_0      (cellSARA_11_io_out_r_input_from_bypass_0     ), //o
    .io_out_r_input_from_bypass_1      (cellSARA_11_io_out_r_input_from_bypass_1     ), //o
    .io_in_c_data_0_data               (cellSARA_11_io_in_c_data_0_data[15:0]        ), //i
    .io_in_c_data_0_is_stationary      (cellSARA_11_io_in_c_data_0_is_stationary     ), //i
    .io_in_c_data_1_data               (cellSARA_11_io_in_c_data_1_data[15:0]        ), //i
    .io_in_c_data_1_is_stationary      (cellSARA_11_io_in_c_data_1_is_stationary     ), //i
    .io_in_c_data_2_data               (cellSARA_11_io_in_c_data_2_data[15:0]        ), //i
    .io_in_c_data_2_is_stationary      (cellSARA_11_io_in_c_data_2_is_stationary     ), //i
    .io_in_c_data_3_data               (cellSARA_11_io_in_c_data_3_data[15:0]        ), //i
    .io_in_c_data_3_is_stationary      (cellSARA_11_io_in_c_data_3_is_stationary     ), //i
    .io_in_c_bypass_0_0_data           (cellSARA_11_io_in_c_bypass_0_0_data[15:0]    ), //i
    .io_in_c_bypass_0_0_is_stationary  (cellSARA_11_io_in_c_bypass_0_0_is_stationary ), //i
    .io_in_c_bypass_0_1_data           (cellSARA_11_io_in_c_bypass_0_1_data[15:0]    ), //i
    .io_in_c_bypass_0_1_is_stationary  (cellSARA_11_io_in_c_bypass_0_1_is_stationary ), //i
    .io_in_c_bypass_0_2_data           (cellSARA_11_io_in_c_bypass_0_2_data[15:0]    ), //i
    .io_in_c_bypass_0_2_is_stationary  (cellSARA_11_io_in_c_bypass_0_2_is_stationary ), //i
    .io_in_c_bypass_0_3_data           (cellSARA_11_io_in_c_bypass_0_3_data[15:0]    ), //i
    .io_in_c_bypass_0_3_is_stationary  (cellSARA_11_io_in_c_bypass_0_3_is_stationary ), //i
    .io_in_c_bypass_1_0_data           (cellSARA_11_io_in_c_bypass_1_0_data[15:0]    ), //i
    .io_in_c_bypass_1_0_is_stationary  (cellSARA_11_io_in_c_bypass_1_0_is_stationary ), //i
    .io_in_c_bypass_1_1_data           (cellSARA_11_io_in_c_bypass_1_1_data[15:0]    ), //i
    .io_in_c_bypass_1_1_is_stationary  (cellSARA_11_io_in_c_bypass_1_1_is_stationary ), //i
    .io_in_c_bypass_1_2_data           (cellSARA_11_io_in_c_bypass_1_2_data[15:0]    ), //i
    .io_in_c_bypass_1_2_is_stationary  (cellSARA_11_io_in_c_bypass_1_2_is_stationary ), //i
    .io_in_c_bypass_1_3_data           (cellSARA_11_io_in_c_bypass_1_3_data[15:0]    ), //i
    .io_in_c_bypass_1_3_is_stationary  (cellSARA_11_io_in_c_bypass_1_3_is_stationary ), //i
    .io_in_c_input_from_bypass_0       (cellSARA_11_io_in_c_input_from_bypass_0      ), //i
    .io_in_c_input_from_bypass_1       (cellSARA_11_io_in_c_input_from_bypass_1      ), //i
    .io_out_c_data_0_data              (cellSARA_11_io_out_c_data_0_data[15:0]       ), //o
    .io_out_c_data_0_is_stationary     (cellSARA_11_io_out_c_data_0_is_stationary    ), //o
    .io_out_c_data_1_data              (cellSARA_11_io_out_c_data_1_data[15:0]       ), //o
    .io_out_c_data_1_is_stationary     (cellSARA_11_io_out_c_data_1_is_stationary    ), //o
    .io_out_c_data_2_data              (cellSARA_11_io_out_c_data_2_data[15:0]       ), //o
    .io_out_c_data_2_is_stationary     (cellSARA_11_io_out_c_data_2_is_stationary    ), //o
    .io_out_c_data_3_data              (cellSARA_11_io_out_c_data_3_data[15:0]       ), //o
    .io_out_c_data_3_is_stationary     (cellSARA_11_io_out_c_data_3_is_stationary    ), //o
    .io_out_c_bypass_0_0_data          (cellSARA_11_io_out_c_bypass_0_0_data[15:0]   ), //o
    .io_out_c_bypass_0_0_is_stationary (cellSARA_11_io_out_c_bypass_0_0_is_stationary), //o
    .io_out_c_bypass_0_1_data          (cellSARA_11_io_out_c_bypass_0_1_data[15:0]   ), //o
    .io_out_c_bypass_0_1_is_stationary (cellSARA_11_io_out_c_bypass_0_1_is_stationary), //o
    .io_out_c_bypass_0_2_data          (cellSARA_11_io_out_c_bypass_0_2_data[15:0]   ), //o
    .io_out_c_bypass_0_2_is_stationary (cellSARA_11_io_out_c_bypass_0_2_is_stationary), //o
    .io_out_c_bypass_0_3_data          (cellSARA_11_io_out_c_bypass_0_3_data[15:0]   ), //o
    .io_out_c_bypass_0_3_is_stationary (cellSARA_11_io_out_c_bypass_0_3_is_stationary), //o
    .io_out_c_bypass_1_0_data          (cellSARA_11_io_out_c_bypass_1_0_data[15:0]   ), //o
    .io_out_c_bypass_1_0_is_stationary (cellSARA_11_io_out_c_bypass_1_0_is_stationary), //o
    .io_out_c_bypass_1_1_data          (cellSARA_11_io_out_c_bypass_1_1_data[15:0]   ), //o
    .io_out_c_bypass_1_1_is_stationary (cellSARA_11_io_out_c_bypass_1_1_is_stationary), //o
    .io_out_c_bypass_1_2_data          (cellSARA_11_io_out_c_bypass_1_2_data[15:0]   ), //o
    .io_out_c_bypass_1_2_is_stationary (cellSARA_11_io_out_c_bypass_1_2_is_stationary), //o
    .io_out_c_bypass_1_3_data          (cellSARA_11_io_out_c_bypass_1_3_data[15:0]   ), //o
    .io_out_c_bypass_1_3_is_stationary (cellSARA_11_io_out_c_bypass_1_3_is_stationary), //o
    .io_out_c_input_from_bypass_0      (cellSARA_11_io_out_c_input_from_bypass_0     ), //o
    .io_out_c_input_from_bypass_1      (cellSARA_11_io_out_c_input_from_bypass_1     ), //o
    .clk                               (clk                                          ), //i
    .reset                             (reset                                        )  //i
  );
  assign io_out_r_0_data_0_data = pes_0_1_io_out_r_data_0_data; // @[SystolicConnect.scala 50:16]
  assign io_out_r_0_data_0_load_store = pes_0_1_io_out_r_data_0_load_store; // @[SystolicConnect.scala 50:16]
  assign io_out_r_0_data_0_df_is_ws = pes_0_1_io_out_r_data_0_df_is_ws; // @[SystolicConnect.scala 50:16]
  assign io_out_r_0_data_0_stall = pes_0_1_io_out_r_data_0_stall; // @[SystolicConnect.scala 50:16]
  assign io_out_r_0_data_1_data = pes_0_1_io_out_r_data_1_data; // @[SystolicConnect.scala 50:16]
  assign io_out_r_0_data_1_load_store = pes_0_1_io_out_r_data_1_load_store; // @[SystolicConnect.scala 50:16]
  assign io_out_r_0_data_1_df_is_ws = pes_0_1_io_out_r_data_1_df_is_ws; // @[SystolicConnect.scala 50:16]
  assign io_out_r_0_data_1_stall = pes_0_1_io_out_r_data_1_stall; // @[SystolicConnect.scala 50:16]
  assign io_out_r_0_data_2_data = pes_0_1_io_out_r_data_2_data; // @[SystolicConnect.scala 50:16]
  assign io_out_r_0_data_2_load_store = pes_0_1_io_out_r_data_2_load_store; // @[SystolicConnect.scala 50:16]
  assign io_out_r_0_data_2_df_is_ws = pes_0_1_io_out_r_data_2_df_is_ws; // @[SystolicConnect.scala 50:16]
  assign io_out_r_0_data_2_stall = pes_0_1_io_out_r_data_2_stall; // @[SystolicConnect.scala 50:16]
  assign io_out_r_0_data_3_data = pes_0_1_io_out_r_data_3_data; // @[SystolicConnect.scala 50:16]
  assign io_out_r_0_data_3_load_store = pes_0_1_io_out_r_data_3_load_store; // @[SystolicConnect.scala 50:16]
  assign io_out_r_0_data_3_df_is_ws = pes_0_1_io_out_r_data_3_df_is_ws; // @[SystolicConnect.scala 50:16]
  assign io_out_r_0_data_3_stall = pes_0_1_io_out_r_data_3_stall; // @[SystolicConnect.scala 50:16]
  assign io_out_r_0_bypass_0_0_data = pes_0_1_io_out_r_bypass_0_0_data; // @[SystolicConnect.scala 50:16]
  assign io_out_r_0_bypass_0_0_load_store = pes_0_1_io_out_r_bypass_0_0_load_store; // @[SystolicConnect.scala 50:16]
  assign io_out_r_0_bypass_0_0_df_is_ws = pes_0_1_io_out_r_bypass_0_0_df_is_ws; // @[SystolicConnect.scala 50:16]
  assign io_out_r_0_bypass_0_0_stall = pes_0_1_io_out_r_bypass_0_0_stall; // @[SystolicConnect.scala 50:16]
  assign io_out_r_0_bypass_0_1_data = pes_0_1_io_out_r_bypass_0_1_data; // @[SystolicConnect.scala 50:16]
  assign io_out_r_0_bypass_0_1_load_store = pes_0_1_io_out_r_bypass_0_1_load_store; // @[SystolicConnect.scala 50:16]
  assign io_out_r_0_bypass_0_1_df_is_ws = pes_0_1_io_out_r_bypass_0_1_df_is_ws; // @[SystolicConnect.scala 50:16]
  assign io_out_r_0_bypass_0_1_stall = pes_0_1_io_out_r_bypass_0_1_stall; // @[SystolicConnect.scala 50:16]
  assign io_out_r_0_bypass_0_2_data = pes_0_1_io_out_r_bypass_0_2_data; // @[SystolicConnect.scala 50:16]
  assign io_out_r_0_bypass_0_2_load_store = pes_0_1_io_out_r_bypass_0_2_load_store; // @[SystolicConnect.scala 50:16]
  assign io_out_r_0_bypass_0_2_df_is_ws = pes_0_1_io_out_r_bypass_0_2_df_is_ws; // @[SystolicConnect.scala 50:16]
  assign io_out_r_0_bypass_0_2_stall = pes_0_1_io_out_r_bypass_0_2_stall; // @[SystolicConnect.scala 50:16]
  assign io_out_r_0_bypass_0_3_data = pes_0_1_io_out_r_bypass_0_3_data; // @[SystolicConnect.scala 50:16]
  assign io_out_r_0_bypass_0_3_load_store = pes_0_1_io_out_r_bypass_0_3_load_store; // @[SystolicConnect.scala 50:16]
  assign io_out_r_0_bypass_0_3_df_is_ws = pes_0_1_io_out_r_bypass_0_3_df_is_ws; // @[SystolicConnect.scala 50:16]
  assign io_out_r_0_bypass_0_3_stall = pes_0_1_io_out_r_bypass_0_3_stall; // @[SystolicConnect.scala 50:16]
  assign io_out_r_0_bypass_1_0_data = pes_0_1_io_out_r_bypass_1_0_data; // @[SystolicConnect.scala 50:16]
  assign io_out_r_0_bypass_1_0_load_store = pes_0_1_io_out_r_bypass_1_0_load_store; // @[SystolicConnect.scala 50:16]
  assign io_out_r_0_bypass_1_0_df_is_ws = pes_0_1_io_out_r_bypass_1_0_df_is_ws; // @[SystolicConnect.scala 50:16]
  assign io_out_r_0_bypass_1_0_stall = pes_0_1_io_out_r_bypass_1_0_stall; // @[SystolicConnect.scala 50:16]
  assign io_out_r_0_bypass_1_1_data = pes_0_1_io_out_r_bypass_1_1_data; // @[SystolicConnect.scala 50:16]
  assign io_out_r_0_bypass_1_1_load_store = pes_0_1_io_out_r_bypass_1_1_load_store; // @[SystolicConnect.scala 50:16]
  assign io_out_r_0_bypass_1_1_df_is_ws = pes_0_1_io_out_r_bypass_1_1_df_is_ws; // @[SystolicConnect.scala 50:16]
  assign io_out_r_0_bypass_1_1_stall = pes_0_1_io_out_r_bypass_1_1_stall; // @[SystolicConnect.scala 50:16]
  assign io_out_r_0_bypass_1_2_data = pes_0_1_io_out_r_bypass_1_2_data; // @[SystolicConnect.scala 50:16]
  assign io_out_r_0_bypass_1_2_load_store = pes_0_1_io_out_r_bypass_1_2_load_store; // @[SystolicConnect.scala 50:16]
  assign io_out_r_0_bypass_1_2_df_is_ws = pes_0_1_io_out_r_bypass_1_2_df_is_ws; // @[SystolicConnect.scala 50:16]
  assign io_out_r_0_bypass_1_2_stall = pes_0_1_io_out_r_bypass_1_2_stall; // @[SystolicConnect.scala 50:16]
  assign io_out_r_0_bypass_1_3_data = pes_0_1_io_out_r_bypass_1_3_data; // @[SystolicConnect.scala 50:16]
  assign io_out_r_0_bypass_1_3_load_store = pes_0_1_io_out_r_bypass_1_3_load_store; // @[SystolicConnect.scala 50:16]
  assign io_out_r_0_bypass_1_3_df_is_ws = pes_0_1_io_out_r_bypass_1_3_df_is_ws; // @[SystolicConnect.scala 50:16]
  assign io_out_r_0_bypass_1_3_stall = pes_0_1_io_out_r_bypass_1_3_stall; // @[SystolicConnect.scala 50:16]
  assign io_out_r_0_input_from_bypass_0 = pes_0_1_io_out_r_input_from_bypass_0; // @[SystolicConnect.scala 50:16]
  assign io_out_r_0_input_from_bypass_1 = pes_0_1_io_out_r_input_from_bypass_1; // @[SystolicConnect.scala 50:16]
  assign io_out_r_1_data_0_data = pes_1_1_io_out_r_data_0_data; // @[SystolicConnect.scala 50:16]
  assign io_out_r_1_data_0_load_store = pes_1_1_io_out_r_data_0_load_store; // @[SystolicConnect.scala 50:16]
  assign io_out_r_1_data_0_df_is_ws = pes_1_1_io_out_r_data_0_df_is_ws; // @[SystolicConnect.scala 50:16]
  assign io_out_r_1_data_0_stall = pes_1_1_io_out_r_data_0_stall; // @[SystolicConnect.scala 50:16]
  assign io_out_r_1_data_1_data = pes_1_1_io_out_r_data_1_data; // @[SystolicConnect.scala 50:16]
  assign io_out_r_1_data_1_load_store = pes_1_1_io_out_r_data_1_load_store; // @[SystolicConnect.scala 50:16]
  assign io_out_r_1_data_1_df_is_ws = pes_1_1_io_out_r_data_1_df_is_ws; // @[SystolicConnect.scala 50:16]
  assign io_out_r_1_data_1_stall = pes_1_1_io_out_r_data_1_stall; // @[SystolicConnect.scala 50:16]
  assign io_out_r_1_data_2_data = pes_1_1_io_out_r_data_2_data; // @[SystolicConnect.scala 50:16]
  assign io_out_r_1_data_2_load_store = pes_1_1_io_out_r_data_2_load_store; // @[SystolicConnect.scala 50:16]
  assign io_out_r_1_data_2_df_is_ws = pes_1_1_io_out_r_data_2_df_is_ws; // @[SystolicConnect.scala 50:16]
  assign io_out_r_1_data_2_stall = pes_1_1_io_out_r_data_2_stall; // @[SystolicConnect.scala 50:16]
  assign io_out_r_1_data_3_data = pes_1_1_io_out_r_data_3_data; // @[SystolicConnect.scala 50:16]
  assign io_out_r_1_data_3_load_store = pes_1_1_io_out_r_data_3_load_store; // @[SystolicConnect.scala 50:16]
  assign io_out_r_1_data_3_df_is_ws = pes_1_1_io_out_r_data_3_df_is_ws; // @[SystolicConnect.scala 50:16]
  assign io_out_r_1_data_3_stall = pes_1_1_io_out_r_data_3_stall; // @[SystolicConnect.scala 50:16]
  assign io_out_r_1_bypass_0_0_data = pes_1_1_io_out_r_bypass_0_0_data; // @[SystolicConnect.scala 50:16]
  assign io_out_r_1_bypass_0_0_load_store = pes_1_1_io_out_r_bypass_0_0_load_store; // @[SystolicConnect.scala 50:16]
  assign io_out_r_1_bypass_0_0_df_is_ws = pes_1_1_io_out_r_bypass_0_0_df_is_ws; // @[SystolicConnect.scala 50:16]
  assign io_out_r_1_bypass_0_0_stall = pes_1_1_io_out_r_bypass_0_0_stall; // @[SystolicConnect.scala 50:16]
  assign io_out_r_1_bypass_0_1_data = pes_1_1_io_out_r_bypass_0_1_data; // @[SystolicConnect.scala 50:16]
  assign io_out_r_1_bypass_0_1_load_store = pes_1_1_io_out_r_bypass_0_1_load_store; // @[SystolicConnect.scala 50:16]
  assign io_out_r_1_bypass_0_1_df_is_ws = pes_1_1_io_out_r_bypass_0_1_df_is_ws; // @[SystolicConnect.scala 50:16]
  assign io_out_r_1_bypass_0_1_stall = pes_1_1_io_out_r_bypass_0_1_stall; // @[SystolicConnect.scala 50:16]
  assign io_out_r_1_bypass_0_2_data = pes_1_1_io_out_r_bypass_0_2_data; // @[SystolicConnect.scala 50:16]
  assign io_out_r_1_bypass_0_2_load_store = pes_1_1_io_out_r_bypass_0_2_load_store; // @[SystolicConnect.scala 50:16]
  assign io_out_r_1_bypass_0_2_df_is_ws = pes_1_1_io_out_r_bypass_0_2_df_is_ws; // @[SystolicConnect.scala 50:16]
  assign io_out_r_1_bypass_0_2_stall = pes_1_1_io_out_r_bypass_0_2_stall; // @[SystolicConnect.scala 50:16]
  assign io_out_r_1_bypass_0_3_data = pes_1_1_io_out_r_bypass_0_3_data; // @[SystolicConnect.scala 50:16]
  assign io_out_r_1_bypass_0_3_load_store = pes_1_1_io_out_r_bypass_0_3_load_store; // @[SystolicConnect.scala 50:16]
  assign io_out_r_1_bypass_0_3_df_is_ws = pes_1_1_io_out_r_bypass_0_3_df_is_ws; // @[SystolicConnect.scala 50:16]
  assign io_out_r_1_bypass_0_3_stall = pes_1_1_io_out_r_bypass_0_3_stall; // @[SystolicConnect.scala 50:16]
  assign io_out_r_1_bypass_1_0_data = pes_1_1_io_out_r_bypass_1_0_data; // @[SystolicConnect.scala 50:16]
  assign io_out_r_1_bypass_1_0_load_store = pes_1_1_io_out_r_bypass_1_0_load_store; // @[SystolicConnect.scala 50:16]
  assign io_out_r_1_bypass_1_0_df_is_ws = pes_1_1_io_out_r_bypass_1_0_df_is_ws; // @[SystolicConnect.scala 50:16]
  assign io_out_r_1_bypass_1_0_stall = pes_1_1_io_out_r_bypass_1_0_stall; // @[SystolicConnect.scala 50:16]
  assign io_out_r_1_bypass_1_1_data = pes_1_1_io_out_r_bypass_1_1_data; // @[SystolicConnect.scala 50:16]
  assign io_out_r_1_bypass_1_1_load_store = pes_1_1_io_out_r_bypass_1_1_load_store; // @[SystolicConnect.scala 50:16]
  assign io_out_r_1_bypass_1_1_df_is_ws = pes_1_1_io_out_r_bypass_1_1_df_is_ws; // @[SystolicConnect.scala 50:16]
  assign io_out_r_1_bypass_1_1_stall = pes_1_1_io_out_r_bypass_1_1_stall; // @[SystolicConnect.scala 50:16]
  assign io_out_r_1_bypass_1_2_data = pes_1_1_io_out_r_bypass_1_2_data; // @[SystolicConnect.scala 50:16]
  assign io_out_r_1_bypass_1_2_load_store = pes_1_1_io_out_r_bypass_1_2_load_store; // @[SystolicConnect.scala 50:16]
  assign io_out_r_1_bypass_1_2_df_is_ws = pes_1_1_io_out_r_bypass_1_2_df_is_ws; // @[SystolicConnect.scala 50:16]
  assign io_out_r_1_bypass_1_2_stall = pes_1_1_io_out_r_bypass_1_2_stall; // @[SystolicConnect.scala 50:16]
  assign io_out_r_1_bypass_1_3_data = pes_1_1_io_out_r_bypass_1_3_data; // @[SystolicConnect.scala 50:16]
  assign io_out_r_1_bypass_1_3_load_store = pes_1_1_io_out_r_bypass_1_3_load_store; // @[SystolicConnect.scala 50:16]
  assign io_out_r_1_bypass_1_3_df_is_ws = pes_1_1_io_out_r_bypass_1_3_df_is_ws; // @[SystolicConnect.scala 50:16]
  assign io_out_r_1_bypass_1_3_stall = pes_1_1_io_out_r_bypass_1_3_stall; // @[SystolicConnect.scala 50:16]
  assign io_out_r_1_input_from_bypass_0 = pes_1_1_io_out_r_input_from_bypass_0; // @[SystolicConnect.scala 50:16]
  assign io_out_r_1_input_from_bypass_1 = pes_1_1_io_out_r_input_from_bypass_1; // @[SystolicConnect.scala 50:16]
  assign io_out_c_0_data_0_data = pes_1_0_io_out_c_data_0_data; // @[SystolicConnect.scala 56:16]
  assign io_out_c_0_data_0_is_stationary = pes_1_0_io_out_c_data_0_is_stationary; // @[SystolicConnect.scala 56:16]
  assign io_out_c_0_data_1_data = pes_1_0_io_out_c_data_1_data; // @[SystolicConnect.scala 56:16]
  assign io_out_c_0_data_1_is_stationary = pes_1_0_io_out_c_data_1_is_stationary; // @[SystolicConnect.scala 56:16]
  assign io_out_c_0_data_2_data = pes_1_0_io_out_c_data_2_data; // @[SystolicConnect.scala 56:16]
  assign io_out_c_0_data_2_is_stationary = pes_1_0_io_out_c_data_2_is_stationary; // @[SystolicConnect.scala 56:16]
  assign io_out_c_0_data_3_data = pes_1_0_io_out_c_data_3_data; // @[SystolicConnect.scala 56:16]
  assign io_out_c_0_data_3_is_stationary = pes_1_0_io_out_c_data_3_is_stationary; // @[SystolicConnect.scala 56:16]
  assign io_out_c_0_bypass_0_0_data = pes_1_0_io_out_c_bypass_0_0_data; // @[SystolicConnect.scala 56:16]
  assign io_out_c_0_bypass_0_0_is_stationary = pes_1_0_io_out_c_bypass_0_0_is_stationary; // @[SystolicConnect.scala 56:16]
  assign io_out_c_0_bypass_0_1_data = pes_1_0_io_out_c_bypass_0_1_data; // @[SystolicConnect.scala 56:16]
  assign io_out_c_0_bypass_0_1_is_stationary = pes_1_0_io_out_c_bypass_0_1_is_stationary; // @[SystolicConnect.scala 56:16]
  assign io_out_c_0_bypass_0_2_data = pes_1_0_io_out_c_bypass_0_2_data; // @[SystolicConnect.scala 56:16]
  assign io_out_c_0_bypass_0_2_is_stationary = pes_1_0_io_out_c_bypass_0_2_is_stationary; // @[SystolicConnect.scala 56:16]
  assign io_out_c_0_bypass_0_3_data = pes_1_0_io_out_c_bypass_0_3_data; // @[SystolicConnect.scala 56:16]
  assign io_out_c_0_bypass_0_3_is_stationary = pes_1_0_io_out_c_bypass_0_3_is_stationary; // @[SystolicConnect.scala 56:16]
  assign io_out_c_0_bypass_1_0_data = pes_1_0_io_out_c_bypass_1_0_data; // @[SystolicConnect.scala 56:16]
  assign io_out_c_0_bypass_1_0_is_stationary = pes_1_0_io_out_c_bypass_1_0_is_stationary; // @[SystolicConnect.scala 56:16]
  assign io_out_c_0_bypass_1_1_data = pes_1_0_io_out_c_bypass_1_1_data; // @[SystolicConnect.scala 56:16]
  assign io_out_c_0_bypass_1_1_is_stationary = pes_1_0_io_out_c_bypass_1_1_is_stationary; // @[SystolicConnect.scala 56:16]
  assign io_out_c_0_bypass_1_2_data = pes_1_0_io_out_c_bypass_1_2_data; // @[SystolicConnect.scala 56:16]
  assign io_out_c_0_bypass_1_2_is_stationary = pes_1_0_io_out_c_bypass_1_2_is_stationary; // @[SystolicConnect.scala 56:16]
  assign io_out_c_0_bypass_1_3_data = pes_1_0_io_out_c_bypass_1_3_data; // @[SystolicConnect.scala 56:16]
  assign io_out_c_0_bypass_1_3_is_stationary = pes_1_0_io_out_c_bypass_1_3_is_stationary; // @[SystolicConnect.scala 56:16]
  assign io_out_c_0_input_from_bypass_0 = pes_1_0_io_out_c_input_from_bypass_0; // @[SystolicConnect.scala 56:16]
  assign io_out_c_0_input_from_bypass_1 = pes_1_0_io_out_c_input_from_bypass_1; // @[SystolicConnect.scala 56:16]
  assign io_out_c_1_data_0_data = pes_1_1_io_out_c_data_0_data; // @[SystolicConnect.scala 56:16]
  assign io_out_c_1_data_0_is_stationary = pes_1_1_io_out_c_data_0_is_stationary; // @[SystolicConnect.scala 56:16]
  assign io_out_c_1_data_1_data = pes_1_1_io_out_c_data_1_data; // @[SystolicConnect.scala 56:16]
  assign io_out_c_1_data_1_is_stationary = pes_1_1_io_out_c_data_1_is_stationary; // @[SystolicConnect.scala 56:16]
  assign io_out_c_1_data_2_data = pes_1_1_io_out_c_data_2_data; // @[SystolicConnect.scala 56:16]
  assign io_out_c_1_data_2_is_stationary = pes_1_1_io_out_c_data_2_is_stationary; // @[SystolicConnect.scala 56:16]
  assign io_out_c_1_data_3_data = pes_1_1_io_out_c_data_3_data; // @[SystolicConnect.scala 56:16]
  assign io_out_c_1_data_3_is_stationary = pes_1_1_io_out_c_data_3_is_stationary; // @[SystolicConnect.scala 56:16]
  assign io_out_c_1_bypass_0_0_data = pes_1_1_io_out_c_bypass_0_0_data; // @[SystolicConnect.scala 56:16]
  assign io_out_c_1_bypass_0_0_is_stationary = pes_1_1_io_out_c_bypass_0_0_is_stationary; // @[SystolicConnect.scala 56:16]
  assign io_out_c_1_bypass_0_1_data = pes_1_1_io_out_c_bypass_0_1_data; // @[SystolicConnect.scala 56:16]
  assign io_out_c_1_bypass_0_1_is_stationary = pes_1_1_io_out_c_bypass_0_1_is_stationary; // @[SystolicConnect.scala 56:16]
  assign io_out_c_1_bypass_0_2_data = pes_1_1_io_out_c_bypass_0_2_data; // @[SystolicConnect.scala 56:16]
  assign io_out_c_1_bypass_0_2_is_stationary = pes_1_1_io_out_c_bypass_0_2_is_stationary; // @[SystolicConnect.scala 56:16]
  assign io_out_c_1_bypass_0_3_data = pes_1_1_io_out_c_bypass_0_3_data; // @[SystolicConnect.scala 56:16]
  assign io_out_c_1_bypass_0_3_is_stationary = pes_1_1_io_out_c_bypass_0_3_is_stationary; // @[SystolicConnect.scala 56:16]
  assign io_out_c_1_bypass_1_0_data = pes_1_1_io_out_c_bypass_1_0_data; // @[SystolicConnect.scala 56:16]
  assign io_out_c_1_bypass_1_0_is_stationary = pes_1_1_io_out_c_bypass_1_0_is_stationary; // @[SystolicConnect.scala 56:16]
  assign io_out_c_1_bypass_1_1_data = pes_1_1_io_out_c_bypass_1_1_data; // @[SystolicConnect.scala 56:16]
  assign io_out_c_1_bypass_1_1_is_stationary = pes_1_1_io_out_c_bypass_1_1_is_stationary; // @[SystolicConnect.scala 56:16]
  assign io_out_c_1_bypass_1_2_data = pes_1_1_io_out_c_bypass_1_2_data; // @[SystolicConnect.scala 56:16]
  assign io_out_c_1_bypass_1_2_is_stationary = pes_1_1_io_out_c_bypass_1_2_is_stationary; // @[SystolicConnect.scala 56:16]
  assign io_out_c_1_bypass_1_3_data = pes_1_1_io_out_c_bypass_1_3_data; // @[SystolicConnect.scala 56:16]
  assign io_out_c_1_bypass_1_3_is_stationary = pes_1_1_io_out_c_bypass_1_3_is_stationary; // @[SystolicConnect.scala 56:16]
  assign io_out_c_1_input_from_bypass_0 = pes_1_1_io_out_c_input_from_bypass_0; // @[SystolicConnect.scala 56:16]
  assign io_out_c_1_input_from_bypass_1 = pes_1_1_io_out_c_input_from_bypass_1; // @[SystolicConnect.scala 56:16]

endmodule

module CellSARA (
  input      [15:0]   io_in_r_data_0_data,
  input               io_in_r_data_0_load_store,
  input               io_in_r_data_0_df_is_ws,
  input               io_in_r_data_0_stall,
  input      [15:0]   io_in_r_data_1_data,
  input               io_in_r_data_1_load_store,
  input               io_in_r_data_1_df_is_ws,
  input               io_in_r_data_1_stall,
  input      [15:0]   io_in_r_data_2_data,
  input               io_in_r_data_2_load_store,
  input               io_in_r_data_2_df_is_ws,
  input               io_in_r_data_2_stall,
  input      [15:0]   io_in_r_data_3_data,
  input               io_in_r_data_3_load_store,
  input               io_in_r_data_3_df_is_ws,
  input               io_in_r_data_3_stall,
  input      [15:0]   io_in_r_bypass_0_0_data,
  input               io_in_r_bypass_0_0_load_store,
  input               io_in_r_bypass_0_0_df_is_ws,
  input               io_in_r_bypass_0_0_stall,
  input      [15:0]   io_in_r_bypass_0_1_data,
  input               io_in_r_bypass_0_1_load_store,
  input               io_in_r_bypass_0_1_df_is_ws,
  input               io_in_r_bypass_0_1_stall,
  input      [15:0]   io_in_r_bypass_0_2_data,
  input               io_in_r_bypass_0_2_load_store,
  input               io_in_r_bypass_0_2_df_is_ws,
  input               io_in_r_bypass_0_2_stall,
  input      [15:0]   io_in_r_bypass_0_3_data,
  input               io_in_r_bypass_0_3_load_store,
  input               io_in_r_bypass_0_3_df_is_ws,
  input               io_in_r_bypass_0_3_stall,
  input      [15:0]   io_in_r_bypass_1_0_data,
  input               io_in_r_bypass_1_0_load_store,
  input               io_in_r_bypass_1_0_df_is_ws,
  input               io_in_r_bypass_1_0_stall,
  input      [15:0]   io_in_r_bypass_1_1_data,
  input               io_in_r_bypass_1_1_load_store,
  input               io_in_r_bypass_1_1_df_is_ws,
  input               io_in_r_bypass_1_1_stall,
  input      [15:0]   io_in_r_bypass_1_2_data,
  input               io_in_r_bypass_1_2_load_store,
  input               io_in_r_bypass_1_2_df_is_ws,
  input               io_in_r_bypass_1_2_stall,
  input      [15:0]   io_in_r_bypass_1_3_data,
  input               io_in_r_bypass_1_3_load_store,
  input               io_in_r_bypass_1_3_df_is_ws,
  input               io_in_r_bypass_1_3_stall,
  input               io_in_r_input_from_bypass_0,
  input               io_in_r_input_from_bypass_1,
  output     [15:0]   io_out_r_data_0_data,
  output              io_out_r_data_0_load_store,
  output              io_out_r_data_0_df_is_ws,
  output              io_out_r_data_0_stall,
  output     [15:0]   io_out_r_data_1_data,
  output              io_out_r_data_1_load_store,
  output              io_out_r_data_1_df_is_ws,
  output              io_out_r_data_1_stall,
  output     [15:0]   io_out_r_data_2_data,
  output              io_out_r_data_2_load_store,
  output              io_out_r_data_2_df_is_ws,
  output              io_out_r_data_2_stall,
  output     [15:0]   io_out_r_data_3_data,
  output              io_out_r_data_3_load_store,
  output              io_out_r_data_3_df_is_ws,
  output              io_out_r_data_3_stall,
  output     [15:0]   io_out_r_bypass_0_0_data,
  output              io_out_r_bypass_0_0_load_store,
  output              io_out_r_bypass_0_0_df_is_ws,
  output              io_out_r_bypass_0_0_stall,
  output     [15:0]   io_out_r_bypass_0_1_data,
  output              io_out_r_bypass_0_1_load_store,
  output              io_out_r_bypass_0_1_df_is_ws,
  output              io_out_r_bypass_0_1_stall,
  output     [15:0]   io_out_r_bypass_0_2_data,
  output              io_out_r_bypass_0_2_load_store,
  output              io_out_r_bypass_0_2_df_is_ws,
  output              io_out_r_bypass_0_2_stall,
  output     [15:0]   io_out_r_bypass_0_3_data,
  output              io_out_r_bypass_0_3_load_store,
  output              io_out_r_bypass_0_3_df_is_ws,
  output              io_out_r_bypass_0_3_stall,
  output     [15:0]   io_out_r_bypass_1_0_data,
  output              io_out_r_bypass_1_0_load_store,
  output              io_out_r_bypass_1_0_df_is_ws,
  output              io_out_r_bypass_1_0_stall,
  output     [15:0]   io_out_r_bypass_1_1_data,
  output              io_out_r_bypass_1_1_load_store,
  output              io_out_r_bypass_1_1_df_is_ws,
  output              io_out_r_bypass_1_1_stall,
  output     [15:0]   io_out_r_bypass_1_2_data,
  output              io_out_r_bypass_1_2_load_store,
  output              io_out_r_bypass_1_2_df_is_ws,
  output              io_out_r_bypass_1_2_stall,
  output     [15:0]   io_out_r_bypass_1_3_data,
  output              io_out_r_bypass_1_3_load_store,
  output              io_out_r_bypass_1_3_df_is_ws,
  output              io_out_r_bypass_1_3_stall,
  output              io_out_r_input_from_bypass_0,
  output              io_out_r_input_from_bypass_1,
  input      [15:0]   io_in_c_data_0_data,
  input               io_in_c_data_0_is_stationary,
  input      [15:0]   io_in_c_data_1_data,
  input               io_in_c_data_1_is_stationary,
  input      [15:0]   io_in_c_data_2_data,
  input               io_in_c_data_2_is_stationary,
  input      [15:0]   io_in_c_data_3_data,
  input               io_in_c_data_3_is_stationary,
  input      [15:0]   io_in_c_bypass_0_0_data,
  input               io_in_c_bypass_0_0_is_stationary,
  input      [15:0]   io_in_c_bypass_0_1_data,
  input               io_in_c_bypass_0_1_is_stationary,
  input      [15:0]   io_in_c_bypass_0_2_data,
  input               io_in_c_bypass_0_2_is_stationary,
  input      [15:0]   io_in_c_bypass_0_3_data,
  input               io_in_c_bypass_0_3_is_stationary,
  input      [15:0]   io_in_c_bypass_1_0_data,
  input               io_in_c_bypass_1_0_is_stationary,
  input      [15:0]   io_in_c_bypass_1_1_data,
  input               io_in_c_bypass_1_1_is_stationary,
  input      [15:0]   io_in_c_bypass_1_2_data,
  input               io_in_c_bypass_1_2_is_stationary,
  input      [15:0]   io_in_c_bypass_1_3_data,
  input               io_in_c_bypass_1_3_is_stationary,
  input               io_in_c_input_from_bypass_0,
  input               io_in_c_input_from_bypass_1,
  output     [15:0]   io_out_c_data_0_data,
  output              io_out_c_data_0_is_stationary,
  output     [15:0]   io_out_c_data_1_data,
  output              io_out_c_data_1_is_stationary,
  output     [15:0]   io_out_c_data_2_data,
  output              io_out_c_data_2_is_stationary,
  output     [15:0]   io_out_c_data_3_data,
  output              io_out_c_data_3_is_stationary,
  output     [15:0]   io_out_c_bypass_0_0_data,
  output              io_out_c_bypass_0_0_is_stationary,
  output     [15:0]   io_out_c_bypass_0_1_data,
  output              io_out_c_bypass_0_1_is_stationary,
  output     [15:0]   io_out_c_bypass_0_2_data,
  output              io_out_c_bypass_0_2_is_stationary,
  output     [15:0]   io_out_c_bypass_0_3_data,
  output              io_out_c_bypass_0_3_is_stationary,
  output     [15:0]   io_out_c_bypass_1_0_data,
  output              io_out_c_bypass_1_0_is_stationary,
  output     [15:0]   io_out_c_bypass_1_1_data,
  output              io_out_c_bypass_1_1_is_stationary,
  output     [15:0]   io_out_c_bypass_1_2_data,
  output              io_out_c_bypass_1_2_is_stationary,
  output     [15:0]   io_out_c_bypass_1_3_data,
  output              io_out_c_bypass_1_3_is_stationary,
  output              io_out_c_input_from_bypass_0,
  output              io_out_c_input_from_bypass_1,
  input               clk,
  input               reset
);

  wire       [15:0]   pes_0_0_io_out_r_data;
  wire                pes_0_0_io_out_r_load_store;
  wire                pes_0_0_io_out_r_df_is_ws;
  wire                pes_0_0_io_out_r_stall;
  wire       [15:0]   pes_0_0_io_out_c_data;
  wire                pes_0_0_io_out_c_is_stationary;
  wire       [15:0]   pes_0_1_io_out_r_data;
  wire                pes_0_1_io_out_r_load_store;
  wire                pes_0_1_io_out_r_df_is_ws;
  wire                pes_0_1_io_out_r_stall;
  wire       [15:0]   pes_0_1_io_out_c_data;
  wire                pes_0_1_io_out_c_is_stationary;
  wire       [15:0]   pes_0_2_io_out_r_data;
  wire                pes_0_2_io_out_r_load_store;
  wire                pes_0_2_io_out_r_df_is_ws;
  wire                pes_0_2_io_out_r_stall;
  wire       [15:0]   pes_0_2_io_out_c_data;
  wire                pes_0_2_io_out_c_is_stationary;
  wire       [15:0]   pes_0_3_io_out_r_data;
  wire                pes_0_3_io_out_r_load_store;
  wire                pes_0_3_io_out_r_df_is_ws;
  wire                pes_0_3_io_out_r_stall;
  wire       [15:0]   pes_0_3_io_out_c_data;
  wire                pes_0_3_io_out_c_is_stationary;
  wire       [15:0]   pes_1_0_io_out_r_data;
  wire                pes_1_0_io_out_r_load_store;
  wire                pes_1_0_io_out_r_df_is_ws;
  wire                pes_1_0_io_out_r_stall;
  wire       [15:0]   pes_1_0_io_out_c_data;
  wire                pes_1_0_io_out_c_is_stationary;
  wire       [15:0]   pes_1_1_io_out_r_data;
  wire                pes_1_1_io_out_r_load_store;
  wire                pes_1_1_io_out_r_df_is_ws;
  wire                pes_1_1_io_out_r_stall;
  wire       [15:0]   pes_1_1_io_out_c_data;
  wire                pes_1_1_io_out_c_is_stationary;
  wire       [15:0]   pes_1_2_io_out_r_data;
  wire                pes_1_2_io_out_r_load_store;
  wire                pes_1_2_io_out_r_df_is_ws;
  wire                pes_1_2_io_out_r_stall;
  wire       [15:0]   pes_1_2_io_out_c_data;
  wire                pes_1_2_io_out_c_is_stationary;
  wire       [15:0]   pes_1_3_io_out_r_data;
  wire                pes_1_3_io_out_r_load_store;
  wire                pes_1_3_io_out_r_df_is_ws;
  wire                pes_1_3_io_out_r_stall;
  wire       [15:0]   pes_1_3_io_out_c_data;
  wire                pes_1_3_io_out_c_is_stationary;
  wire       [15:0]   pes_2_0_io_out_r_data;
  wire                pes_2_0_io_out_r_load_store;
  wire                pes_2_0_io_out_r_df_is_ws;
  wire                pes_2_0_io_out_r_stall;
  wire       [15:0]   pes_2_0_io_out_c_data;
  wire                pes_2_0_io_out_c_is_stationary;
  wire       [15:0]   pes_2_1_io_out_r_data;
  wire                pes_2_1_io_out_r_load_store;
  wire                pes_2_1_io_out_r_df_is_ws;
  wire                pes_2_1_io_out_r_stall;
  wire       [15:0]   pes_2_1_io_out_c_data;
  wire                pes_2_1_io_out_c_is_stationary;
  wire       [15:0]   pes_2_2_io_out_r_data;
  wire                pes_2_2_io_out_r_load_store;
  wire                pes_2_2_io_out_r_df_is_ws;
  wire                pes_2_2_io_out_r_stall;
  wire       [15:0]   pes_2_2_io_out_c_data;
  wire                pes_2_2_io_out_c_is_stationary;
  wire       [15:0]   pes_2_3_io_out_r_data;
  wire                pes_2_3_io_out_r_load_store;
  wire                pes_2_3_io_out_r_df_is_ws;
  wire                pes_2_3_io_out_r_stall;
  wire       [15:0]   pes_2_3_io_out_c_data;
  wire                pes_2_3_io_out_c_is_stationary;
  wire       [15:0]   pes_3_0_io_out_r_data;
  wire                pes_3_0_io_out_r_load_store;
  wire                pes_3_0_io_out_r_df_is_ws;
  wire                pes_3_0_io_out_r_stall;
  wire       [15:0]   pes_3_0_io_out_c_data;
  wire                pes_3_0_io_out_c_is_stationary;
  wire       [15:0]   pes_3_1_io_out_r_data;
  wire                pes_3_1_io_out_r_load_store;
  wire                pes_3_1_io_out_r_df_is_ws;
  wire                pes_3_1_io_out_r_stall;
  wire       [15:0]   pes_3_1_io_out_c_data;
  wire                pes_3_1_io_out_c_is_stationary;
  wire       [15:0]   pes_3_2_io_out_r_data;
  wire                pes_3_2_io_out_r_load_store;
  wire                pes_3_2_io_out_r_df_is_ws;
  wire                pes_3_2_io_out_r_stall;
  wire       [15:0]   pes_3_2_io_out_c_data;
  wire                pes_3_2_io_out_c_is_stationary;
  wire       [15:0]   pes_3_3_io_out_r_data;
  wire                pes_3_3_io_out_r_load_store;
  wire                pes_3_3_io_out_r_df_is_ws;
  wire                pes_3_3_io_out_r_stall;
  wire       [15:0]   pes_3_3_io_out_c_data;
  wire                pes_3_3_io_out_c_is_stationary;
  wire       [15:0]   in_r_0_data;
  wire                in_r_0_load_store;
  wire                in_r_0_df_is_ws;
  wire                in_r_0_stall;
  wire       [15:0]   in_r_1_data;
  wire                in_r_1_load_store;
  wire                in_r_1_df_is_ws;
  wire                in_r_1_stall;
  wire       [15:0]   in_r_2_data;
  wire                in_r_2_load_store;
  wire                in_r_2_df_is_ws;
  wire                in_r_2_stall;
  wire       [15:0]   in_r_3_data;
  wire                in_r_3_load_store;
  wire                in_r_3_df_is_ws;
  wire                in_r_3_stall;
  wire       [15:0]   in_c_0_data;
  wire                in_c_0_is_stationary;
  wire       [15:0]   in_c_1_data;
  wire                in_c_1_is_stationary;
  wire       [15:0]   in_c_2_data;
  wire                in_c_2_is_stationary;
  wire       [15:0]   in_c_3_data;
  wire                in_c_3_is_stationary;
  wire       [15:0]   out_r_0_data;
  wire                out_r_0_load_store;
  wire                out_r_0_df_is_ws;
  wire                out_r_0_stall;
  wire       [15:0]   out_r_1_data;
  wire                out_r_1_load_store;
  wire                out_r_1_df_is_ws;
  wire                out_r_1_stall;
  wire       [15:0]   out_r_2_data;
  wire                out_r_2_load_store;
  wire                out_r_2_df_is_ws;
  wire                out_r_2_stall;
  wire       [15:0]   out_r_3_data;
  wire                out_r_3_load_store;
  wire                out_r_3_df_is_ws;
  wire                out_r_3_stall;
  wire       [15:0]   out_c_0_data;
  wire                out_c_0_is_stationary;
  wire       [15:0]   out_c_1_data;
  wire                out_c_1_is_stationary;
  wire       [15:0]   out_c_2_data;
  wire                out_c_2_is_stationary;
  wire       [15:0]   out_c_3_data;
  wire                out_c_3_is_stationary;
  reg        [15:0]   out_r_regNext_0_data;
  reg                 out_r_regNext_0_load_store;
  reg                 out_r_regNext_0_df_is_ws;
  reg                 out_r_regNext_0_stall;
  reg        [15:0]   out_r_regNext_1_data;
  reg                 out_r_regNext_1_load_store;
  reg                 out_r_regNext_1_df_is_ws;
  reg                 out_r_regNext_1_stall;
  reg        [15:0]   out_r_regNext_2_data;
  reg                 out_r_regNext_2_load_store;
  reg                 out_r_regNext_2_df_is_ws;
  reg                 out_r_regNext_2_stall;
  reg        [15:0]   out_r_regNext_3_data;
  reg                 out_r_regNext_3_load_store;
  reg                 out_r_regNext_3_df_is_ws;
  reg                 out_r_regNext_3_stall;
  reg        [15:0]   out_c_regNext_0_data;
  reg                 out_c_regNext_0_is_stationary;
  reg        [15:0]   out_c_regNext_1_data;
  reg                 out_c_regNext_1_is_stationary;
  reg        [15:0]   out_c_regNext_2_data;
  reg                 out_c_regNext_2_is_stationary;
  reg        [15:0]   out_c_regNext_3_data;
  reg                 out_c_regNext_3_is_stationary;
  reg        [15:0]   io_in_r_bypass_regNext_0_0_data;
  reg                 io_in_r_bypass_regNext_0_0_load_store;
  reg                 io_in_r_bypass_regNext_0_0_df_is_ws;
  reg                 io_in_r_bypass_regNext_0_0_stall;
  reg        [15:0]   io_in_r_bypass_regNext_0_1_data;
  reg                 io_in_r_bypass_regNext_0_1_load_store;
  reg                 io_in_r_bypass_regNext_0_1_df_is_ws;
  reg                 io_in_r_bypass_regNext_0_1_stall;
  reg        [15:0]   io_in_r_bypass_regNext_0_2_data;
  reg                 io_in_r_bypass_regNext_0_2_load_store;
  reg                 io_in_r_bypass_regNext_0_2_df_is_ws;
  reg                 io_in_r_bypass_regNext_0_2_stall;
  reg        [15:0]   io_in_r_bypass_regNext_0_3_data;
  reg                 io_in_r_bypass_regNext_0_3_load_store;
  reg                 io_in_r_bypass_regNext_0_3_df_is_ws;
  reg                 io_in_r_bypass_regNext_0_3_stall;
  reg        [15:0]   io_in_r_bypass_regNext_1_0_data;
  reg                 io_in_r_bypass_regNext_1_0_load_store;
  reg                 io_in_r_bypass_regNext_1_0_df_is_ws;
  reg                 io_in_r_bypass_regNext_1_0_stall;
  reg        [15:0]   io_in_r_bypass_regNext_1_1_data;
  reg                 io_in_r_bypass_regNext_1_1_load_store;
  reg                 io_in_r_bypass_regNext_1_1_df_is_ws;
  reg                 io_in_r_bypass_regNext_1_1_stall;
  reg        [15:0]   io_in_r_bypass_regNext_1_2_data;
  reg                 io_in_r_bypass_regNext_1_2_load_store;
  reg                 io_in_r_bypass_regNext_1_2_df_is_ws;
  reg                 io_in_r_bypass_regNext_1_2_stall;
  reg        [15:0]   io_in_r_bypass_regNext_1_3_data;
  reg                 io_in_r_bypass_regNext_1_3_load_store;
  reg                 io_in_r_bypass_regNext_1_3_df_is_ws;
  reg                 io_in_r_bypass_regNext_1_3_stall;
  reg        [15:0]   io_in_c_bypass_regNext_0_0_data;
  reg                 io_in_c_bypass_regNext_0_0_is_stationary;
  reg        [15:0]   io_in_c_bypass_regNext_0_1_data;
  reg                 io_in_c_bypass_regNext_0_1_is_stationary;
  reg        [15:0]   io_in_c_bypass_regNext_0_2_data;
  reg                 io_in_c_bypass_regNext_0_2_is_stationary;
  reg        [15:0]   io_in_c_bypass_regNext_0_3_data;
  reg                 io_in_c_bypass_regNext_0_3_is_stationary;
  reg        [15:0]   io_in_c_bypass_regNext_1_0_data;
  reg                 io_in_c_bypass_regNext_1_0_is_stationary;
  reg        [15:0]   io_in_c_bypass_regNext_1_1_data;
  reg                 io_in_c_bypass_regNext_1_1_is_stationary;
  reg        [15:0]   io_in_c_bypass_regNext_1_2_data;
  reg                 io_in_c_bypass_regNext_1_2_is_stationary;
  reg        [15:0]   io_in_c_bypass_regNext_1_3_data;
  reg                 io_in_c_bypass_regNext_1_3_is_stationary;
  reg                 io_in_r_input_from_bypass_regNext_0;
  reg                 io_in_r_input_from_bypass_regNext_1;
  reg                 io_in_c_input_from_bypass_regNext_0;
  reg                 io_in_c_input_from_bypass_regNext_1;

  PEWSOS_127 pes_0_0 (
    .io_in_r_data           (in_r_0_data[15:0]             ), //i
    .io_in_r_load_store     (in_r_0_load_store             ), //i
    .io_in_r_df_is_ws       (in_r_0_df_is_ws               ), //i
    .io_in_r_stall          (in_r_0_stall                  ), //i
    .io_out_r_data          (pes_0_0_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pes_0_0_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pes_0_0_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pes_0_0_io_out_r_stall        ), //o
    .io_in_c_data           (in_c_0_data[15:0]             ), //i
    .io_in_c_is_stationary  (in_c_0_is_stationary          ), //i
    .io_out_c_data          (pes_0_0_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pes_0_0_io_out_c_is_stationary), //o
    .clk                    (clk                           ), //i
    .reset                  (reset                         )  //i
  );
  PEWSOS_127 pes_0_1 (
    .io_in_r_data           (pes_0_0_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pes_0_0_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pes_0_0_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pes_0_0_io_out_r_stall        ), //i
    .io_out_r_data          (pes_0_1_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pes_0_1_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pes_0_1_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pes_0_1_io_out_r_stall        ), //o
    .io_in_c_data           (in_c_1_data[15:0]             ), //i
    .io_in_c_is_stationary  (in_c_1_is_stationary          ), //i
    .io_out_c_data          (pes_0_1_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pes_0_1_io_out_c_is_stationary), //o
    .clk                    (clk                           ), //i
    .reset                  (reset                         )  //i
  );
  PEWSOS_127 pes_0_2 (
    .io_in_r_data           (pes_0_1_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pes_0_1_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pes_0_1_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pes_0_1_io_out_r_stall        ), //i
    .io_out_r_data          (pes_0_2_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pes_0_2_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pes_0_2_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pes_0_2_io_out_r_stall        ), //o
    .io_in_c_data           (in_c_2_data[15:0]             ), //i
    .io_in_c_is_stationary  (in_c_2_is_stationary          ), //i
    .io_out_c_data          (pes_0_2_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pes_0_2_io_out_c_is_stationary), //o
    .clk                    (clk                           ), //i
    .reset                  (reset                         )  //i
  );
  PEWSOS_127 pes_0_3 (
    .io_in_r_data           (pes_0_2_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pes_0_2_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pes_0_2_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pes_0_2_io_out_r_stall        ), //i
    .io_out_r_data          (pes_0_3_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pes_0_3_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pes_0_3_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pes_0_3_io_out_r_stall        ), //o
    .io_in_c_data           (in_c_3_data[15:0]             ), //i
    .io_in_c_is_stationary  (in_c_3_is_stationary          ), //i
    .io_out_c_data          (pes_0_3_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pes_0_3_io_out_c_is_stationary), //o
    .clk                    (clk                           ), //i
    .reset                  (reset                         )  //i
  );
  PEWSOS_127 pes_1_0 (
    .io_in_r_data           (in_r_1_data[15:0]             ), //i
    .io_in_r_load_store     (in_r_1_load_store             ), //i
    .io_in_r_df_is_ws       (in_r_1_df_is_ws               ), //i
    .io_in_r_stall          (in_r_1_stall                  ), //i
    .io_out_r_data          (pes_1_0_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pes_1_0_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pes_1_0_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pes_1_0_io_out_r_stall        ), //o
    .io_in_c_data           (pes_0_0_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pes_0_0_io_out_c_is_stationary), //i
    .io_out_c_data          (pes_1_0_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pes_1_0_io_out_c_is_stationary), //o
    .clk                    (clk                           ), //i
    .reset                  (reset                         )  //i
  );
  PEWSOS_127 pes_1_1 (
    .io_in_r_data           (pes_1_0_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pes_1_0_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pes_1_0_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pes_1_0_io_out_r_stall        ), //i
    .io_out_r_data          (pes_1_1_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pes_1_1_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pes_1_1_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pes_1_1_io_out_r_stall        ), //o
    .io_in_c_data           (pes_0_1_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pes_0_1_io_out_c_is_stationary), //i
    .io_out_c_data          (pes_1_1_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pes_1_1_io_out_c_is_stationary), //o
    .clk                    (clk                           ), //i
    .reset                  (reset                         )  //i
  );
  PEWSOS_127 pes_1_2 (
    .io_in_r_data           (pes_1_1_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pes_1_1_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pes_1_1_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pes_1_1_io_out_r_stall        ), //i
    .io_out_r_data          (pes_1_2_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pes_1_2_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pes_1_2_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pes_1_2_io_out_r_stall        ), //o
    .io_in_c_data           (pes_0_2_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pes_0_2_io_out_c_is_stationary), //i
    .io_out_c_data          (pes_1_2_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pes_1_2_io_out_c_is_stationary), //o
    .clk                    (clk                           ), //i
    .reset                  (reset                         )  //i
  );
  PEWSOS_127 pes_1_3 (
    .io_in_r_data           (pes_1_2_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pes_1_2_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pes_1_2_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pes_1_2_io_out_r_stall        ), //i
    .io_out_r_data          (pes_1_3_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pes_1_3_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pes_1_3_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pes_1_3_io_out_r_stall        ), //o
    .io_in_c_data           (pes_0_3_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pes_0_3_io_out_c_is_stationary), //i
    .io_out_c_data          (pes_1_3_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pes_1_3_io_out_c_is_stationary), //o
    .clk                    (clk                           ), //i
    .reset                  (reset                         )  //i
  );
  PEWSOS_127 pes_2_0 (
    .io_in_r_data           (in_r_2_data[15:0]             ), //i
    .io_in_r_load_store     (in_r_2_load_store             ), //i
    .io_in_r_df_is_ws       (in_r_2_df_is_ws               ), //i
    .io_in_r_stall          (in_r_2_stall                  ), //i
    .io_out_r_data          (pes_2_0_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pes_2_0_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pes_2_0_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pes_2_0_io_out_r_stall        ), //o
    .io_in_c_data           (pes_1_0_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pes_1_0_io_out_c_is_stationary), //i
    .io_out_c_data          (pes_2_0_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pes_2_0_io_out_c_is_stationary), //o
    .clk                    (clk                           ), //i
    .reset                  (reset                         )  //i
  );
  PEWSOS_127 pes_2_1 (
    .io_in_r_data           (pes_2_0_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pes_2_0_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pes_2_0_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pes_2_0_io_out_r_stall        ), //i
    .io_out_r_data          (pes_2_1_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pes_2_1_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pes_2_1_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pes_2_1_io_out_r_stall        ), //o
    .io_in_c_data           (pes_1_1_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pes_1_1_io_out_c_is_stationary), //i
    .io_out_c_data          (pes_2_1_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pes_2_1_io_out_c_is_stationary), //o
    .clk                    (clk                           ), //i
    .reset                  (reset                         )  //i
  );
  PEWSOS_127 pes_2_2 (
    .io_in_r_data           (pes_2_1_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pes_2_1_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pes_2_1_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pes_2_1_io_out_r_stall        ), //i
    .io_out_r_data          (pes_2_2_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pes_2_2_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pes_2_2_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pes_2_2_io_out_r_stall        ), //o
    .io_in_c_data           (pes_1_2_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pes_1_2_io_out_c_is_stationary), //i
    .io_out_c_data          (pes_2_2_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pes_2_2_io_out_c_is_stationary), //o
    .clk                    (clk                           ), //i
    .reset                  (reset                         )  //i
  );
  PEWSOS_127 pes_2_3 (
    .io_in_r_data           (pes_2_2_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pes_2_2_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pes_2_2_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pes_2_2_io_out_r_stall        ), //i
    .io_out_r_data          (pes_2_3_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pes_2_3_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pes_2_3_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pes_2_3_io_out_r_stall        ), //o
    .io_in_c_data           (pes_1_3_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pes_1_3_io_out_c_is_stationary), //i
    .io_out_c_data          (pes_2_3_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pes_2_3_io_out_c_is_stationary), //o
    .clk                    (clk                           ), //i
    .reset                  (reset                         )  //i
  );
  PEWSOS_127 pes_3_0 (
    .io_in_r_data           (in_r_3_data[15:0]             ), //i
    .io_in_r_load_store     (in_r_3_load_store             ), //i
    .io_in_r_df_is_ws       (in_r_3_df_is_ws               ), //i
    .io_in_r_stall          (in_r_3_stall                  ), //i
    .io_out_r_data          (pes_3_0_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pes_3_0_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pes_3_0_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pes_3_0_io_out_r_stall        ), //o
    .io_in_c_data           (pes_2_0_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pes_2_0_io_out_c_is_stationary), //i
    .io_out_c_data          (pes_3_0_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pes_3_0_io_out_c_is_stationary), //o
    .clk                    (clk                           ), //i
    .reset                  (reset                         )  //i
  );
  PEWSOS_127 pes_3_1 (
    .io_in_r_data           (pes_3_0_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pes_3_0_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pes_3_0_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pes_3_0_io_out_r_stall        ), //i
    .io_out_r_data          (pes_3_1_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pes_3_1_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pes_3_1_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pes_3_1_io_out_r_stall        ), //o
    .io_in_c_data           (pes_2_1_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pes_2_1_io_out_c_is_stationary), //i
    .io_out_c_data          (pes_3_1_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pes_3_1_io_out_c_is_stationary), //o
    .clk                    (clk                           ), //i
    .reset                  (reset                         )  //i
  );
  PEWSOS_127 pes_3_2 (
    .io_in_r_data           (pes_3_1_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pes_3_1_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pes_3_1_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pes_3_1_io_out_r_stall        ), //i
    .io_out_r_data          (pes_3_2_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pes_3_2_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pes_3_2_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pes_3_2_io_out_r_stall        ), //o
    .io_in_c_data           (pes_2_2_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pes_2_2_io_out_c_is_stationary), //i
    .io_out_c_data          (pes_3_2_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pes_3_2_io_out_c_is_stationary), //o
    .clk                    (clk                           ), //i
    .reset                  (reset                         )  //i
  );
  PEWSOS_127 pes_3_3 (
    .io_in_r_data           (pes_3_2_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pes_3_2_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pes_3_2_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pes_3_2_io_out_r_stall        ), //i
    .io_out_r_data          (pes_3_3_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pes_3_3_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pes_3_3_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pes_3_3_io_out_r_stall        ), //o
    .io_in_c_data           (pes_2_3_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pes_2_3_io_out_c_is_stationary), //i
    .io_out_c_data          (pes_3_3_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pes_3_3_io_out_c_is_stationary), //o
    .clk                    (clk                           ), //i
    .reset                  (reset                         )  //i
  );
  assign in_r_0_data = (io_in_r_input_from_bypass_1 ? io_in_r_bypass_1_0_data : io_in_r_data_0_data); // @[Expression.scala 1420:25]
  assign in_r_0_load_store = (io_in_r_input_from_bypass_1 ? io_in_r_bypass_1_0_load_store : io_in_r_data_0_load_store); // @[Expression.scala 1420:25]
  assign in_r_0_df_is_ws = (io_in_r_input_from_bypass_1 ? io_in_r_bypass_1_0_df_is_ws : io_in_r_data_0_df_is_ws); // @[Expression.scala 1420:25]
  assign in_r_0_stall = (io_in_r_input_from_bypass_1 ? io_in_r_bypass_1_0_stall : io_in_r_data_0_stall); // @[Expression.scala 1420:25]
  assign in_r_1_data = (io_in_r_input_from_bypass_1 ? io_in_r_bypass_1_1_data : io_in_r_data_1_data); // @[Expression.scala 1420:25]
  assign in_r_1_load_store = (io_in_r_input_from_bypass_1 ? io_in_r_bypass_1_1_load_store : io_in_r_data_1_load_store); // @[Expression.scala 1420:25]
  assign in_r_1_df_is_ws = (io_in_r_input_from_bypass_1 ? io_in_r_bypass_1_1_df_is_ws : io_in_r_data_1_df_is_ws); // @[Expression.scala 1420:25]
  assign in_r_1_stall = (io_in_r_input_from_bypass_1 ? io_in_r_bypass_1_1_stall : io_in_r_data_1_stall); // @[Expression.scala 1420:25]
  assign in_r_2_data = (io_in_r_input_from_bypass_1 ? io_in_r_bypass_1_2_data : io_in_r_data_2_data); // @[Expression.scala 1420:25]
  assign in_r_2_load_store = (io_in_r_input_from_bypass_1 ? io_in_r_bypass_1_2_load_store : io_in_r_data_2_load_store); // @[Expression.scala 1420:25]
  assign in_r_2_df_is_ws = (io_in_r_input_from_bypass_1 ? io_in_r_bypass_1_2_df_is_ws : io_in_r_data_2_df_is_ws); // @[Expression.scala 1420:25]
  assign in_r_2_stall = (io_in_r_input_from_bypass_1 ? io_in_r_bypass_1_2_stall : io_in_r_data_2_stall); // @[Expression.scala 1420:25]
  assign in_r_3_data = (io_in_r_input_from_bypass_1 ? io_in_r_bypass_1_3_data : io_in_r_data_3_data); // @[Expression.scala 1420:25]
  assign in_r_3_load_store = (io_in_r_input_from_bypass_1 ? io_in_r_bypass_1_3_load_store : io_in_r_data_3_load_store); // @[Expression.scala 1420:25]
  assign in_r_3_df_is_ws = (io_in_r_input_from_bypass_1 ? io_in_r_bypass_1_3_df_is_ws : io_in_r_data_3_df_is_ws); // @[Expression.scala 1420:25]
  assign in_r_3_stall = (io_in_r_input_from_bypass_1 ? io_in_r_bypass_1_3_stall : io_in_r_data_3_stall); // @[Expression.scala 1420:25]
  assign in_c_0_data = (io_in_c_input_from_bypass_1 ? io_in_c_bypass_1_0_data : io_in_c_data_0_data); // @[Expression.scala 1420:25]
  assign in_c_0_is_stationary = (io_in_c_input_from_bypass_1 ? io_in_c_bypass_1_0_is_stationary : io_in_c_data_0_is_stationary); // @[Expression.scala 1420:25]
  assign in_c_1_data = (io_in_c_input_from_bypass_1 ? io_in_c_bypass_1_1_data : io_in_c_data_1_data); // @[Expression.scala 1420:25]
  assign in_c_1_is_stationary = (io_in_c_input_from_bypass_1 ? io_in_c_bypass_1_1_is_stationary : io_in_c_data_1_is_stationary); // @[Expression.scala 1420:25]
  assign in_c_2_data = (io_in_c_input_from_bypass_1 ? io_in_c_bypass_1_2_data : io_in_c_data_2_data); // @[Expression.scala 1420:25]
  assign in_c_2_is_stationary = (io_in_c_input_from_bypass_1 ? io_in_c_bypass_1_2_is_stationary : io_in_c_data_2_is_stationary); // @[Expression.scala 1420:25]
  assign in_c_3_data = (io_in_c_input_from_bypass_1 ? io_in_c_bypass_1_3_data : io_in_c_data_3_data); // @[Expression.scala 1420:25]
  assign in_c_3_is_stationary = (io_in_c_input_from_bypass_1 ? io_in_c_bypass_1_3_is_stationary : io_in_c_data_3_is_stationary); // @[Expression.scala 1420:25]
  assign out_r_0_data = pes_0_3_io_out_r_data; // @[SystolicConnect.scala 50:16]
  assign out_r_0_load_store = pes_0_3_io_out_r_load_store; // @[SystolicConnect.scala 50:16]
  assign out_r_0_df_is_ws = pes_0_3_io_out_r_df_is_ws; // @[SystolicConnect.scala 50:16]
  assign out_r_0_stall = pes_0_3_io_out_r_stall; // @[SystolicConnect.scala 50:16]
  assign out_r_1_data = pes_1_3_io_out_r_data; // @[SystolicConnect.scala 50:16]
  assign out_r_1_load_store = pes_1_3_io_out_r_load_store; // @[SystolicConnect.scala 50:16]
  assign out_r_1_df_is_ws = pes_1_3_io_out_r_df_is_ws; // @[SystolicConnect.scala 50:16]
  assign out_r_1_stall = pes_1_3_io_out_r_stall; // @[SystolicConnect.scala 50:16]
  assign out_r_2_data = pes_2_3_io_out_r_data; // @[SystolicConnect.scala 50:16]
  assign out_r_2_load_store = pes_2_3_io_out_r_load_store; // @[SystolicConnect.scala 50:16]
  assign out_r_2_df_is_ws = pes_2_3_io_out_r_df_is_ws; // @[SystolicConnect.scala 50:16]
  assign out_r_2_stall = pes_2_3_io_out_r_stall; // @[SystolicConnect.scala 50:16]
  assign out_r_3_data = pes_3_3_io_out_r_data; // @[SystolicConnect.scala 50:16]
  assign out_r_3_load_store = pes_3_3_io_out_r_load_store; // @[SystolicConnect.scala 50:16]
  assign out_r_3_df_is_ws = pes_3_3_io_out_r_df_is_ws; // @[SystolicConnect.scala 50:16]
  assign out_r_3_stall = pes_3_3_io_out_r_stall; // @[SystolicConnect.scala 50:16]
  assign out_c_0_data = pes_3_0_io_out_c_data; // @[SystolicConnect.scala 56:16]
  assign out_c_0_is_stationary = pes_3_0_io_out_c_is_stationary; // @[SystolicConnect.scala 56:16]
  assign out_c_1_data = pes_3_1_io_out_c_data; // @[SystolicConnect.scala 56:16]
  assign out_c_1_is_stationary = pes_3_1_io_out_c_is_stationary; // @[SystolicConnect.scala 56:16]
  assign out_c_2_data = pes_3_2_io_out_c_data; // @[SystolicConnect.scala 56:16]
  assign out_c_2_is_stationary = pes_3_2_io_out_c_is_stationary; // @[SystolicConnect.scala 56:16]
  assign out_c_3_data = pes_3_3_io_out_c_data; // @[SystolicConnect.scala 56:16]
  assign out_c_3_is_stationary = pes_3_3_io_out_c_is_stationary; // @[SystolicConnect.scala 56:16]
  assign io_out_r_data_0_data = out_r_0_data; // @[ArraySARA.scala 90:17]
  assign io_out_r_data_0_load_store = out_r_0_load_store; // @[ArraySARA.scala 90:17]
  assign io_out_r_data_0_df_is_ws = out_r_0_df_is_ws; // @[ArraySARA.scala 90:17]
  assign io_out_r_data_0_stall = out_r_0_stall; // @[ArraySARA.scala 90:17]
  assign io_out_r_data_1_data = out_r_1_data; // @[ArraySARA.scala 90:17]
  assign io_out_r_data_1_load_store = out_r_1_load_store; // @[ArraySARA.scala 90:17]
  assign io_out_r_data_1_df_is_ws = out_r_1_df_is_ws; // @[ArraySARA.scala 90:17]
  assign io_out_r_data_1_stall = out_r_1_stall; // @[ArraySARA.scala 90:17]
  assign io_out_r_data_2_data = out_r_2_data; // @[ArraySARA.scala 90:17]
  assign io_out_r_data_2_load_store = out_r_2_load_store; // @[ArraySARA.scala 90:17]
  assign io_out_r_data_2_df_is_ws = out_r_2_df_is_ws; // @[ArraySARA.scala 90:17]
  assign io_out_r_data_2_stall = out_r_2_stall; // @[ArraySARA.scala 90:17]
  assign io_out_r_data_3_data = out_r_3_data; // @[ArraySARA.scala 90:17]
  assign io_out_r_data_3_load_store = out_r_3_load_store; // @[ArraySARA.scala 90:17]
  assign io_out_r_data_3_df_is_ws = out_r_3_df_is_ws; // @[ArraySARA.scala 90:17]
  assign io_out_r_data_3_stall = out_r_3_stall; // @[ArraySARA.scala 90:17]
  assign io_out_c_data_0_data = out_c_0_data; // @[ArraySARA.scala 91:17]
  assign io_out_c_data_0_is_stationary = out_c_0_is_stationary; // @[ArraySARA.scala 91:17]
  assign io_out_c_data_1_data = out_c_1_data; // @[ArraySARA.scala 91:17]
  assign io_out_c_data_1_is_stationary = out_c_1_is_stationary; // @[ArraySARA.scala 91:17]
  assign io_out_c_data_2_data = out_c_2_data; // @[ArraySARA.scala 91:17]
  assign io_out_c_data_2_is_stationary = out_c_2_is_stationary; // @[ArraySARA.scala 91:17]
  assign io_out_c_data_3_data = out_c_3_data; // @[ArraySARA.scala 91:17]
  assign io_out_c_data_3_is_stationary = out_c_3_is_stationary; // @[ArraySARA.scala 91:17]
  assign io_out_r_bypass_1_0_data = out_r_regNext_0_data; // @[ArraySARA.scala 92:31]
  assign io_out_r_bypass_1_0_load_store = out_r_regNext_0_load_store; // @[ArraySARA.scala 92:31]
  assign io_out_r_bypass_1_0_df_is_ws = out_r_regNext_0_df_is_ws; // @[ArraySARA.scala 92:31]
  assign io_out_r_bypass_1_0_stall = out_r_regNext_0_stall; // @[ArraySARA.scala 92:31]
  assign io_out_r_bypass_1_1_data = out_r_regNext_1_data; // @[ArraySARA.scala 92:31]
  assign io_out_r_bypass_1_1_load_store = out_r_regNext_1_load_store; // @[ArraySARA.scala 92:31]
  assign io_out_r_bypass_1_1_df_is_ws = out_r_regNext_1_df_is_ws; // @[ArraySARA.scala 92:31]
  assign io_out_r_bypass_1_1_stall = out_r_regNext_1_stall; // @[ArraySARA.scala 92:31]
  assign io_out_r_bypass_1_2_data = out_r_regNext_2_data; // @[ArraySARA.scala 92:31]
  assign io_out_r_bypass_1_2_load_store = out_r_regNext_2_load_store; // @[ArraySARA.scala 92:31]
  assign io_out_r_bypass_1_2_df_is_ws = out_r_regNext_2_df_is_ws; // @[ArraySARA.scala 92:31]
  assign io_out_r_bypass_1_2_stall = out_r_regNext_2_stall; // @[ArraySARA.scala 92:31]
  assign io_out_r_bypass_1_3_data = out_r_regNext_3_data; // @[ArraySARA.scala 92:31]
  assign io_out_r_bypass_1_3_load_store = out_r_regNext_3_load_store; // @[ArraySARA.scala 92:31]
  assign io_out_r_bypass_1_3_df_is_ws = out_r_regNext_3_df_is_ws; // @[ArraySARA.scala 92:31]
  assign io_out_r_bypass_1_3_stall = out_r_regNext_3_stall; // @[ArraySARA.scala 92:31]
  assign io_out_c_bypass_1_0_data = out_c_regNext_0_data; // @[ArraySARA.scala 93:31]
  assign io_out_c_bypass_1_0_is_stationary = out_c_regNext_0_is_stationary; // @[ArraySARA.scala 93:31]
  assign io_out_c_bypass_1_1_data = out_c_regNext_1_data; // @[ArraySARA.scala 93:31]
  assign io_out_c_bypass_1_1_is_stationary = out_c_regNext_1_is_stationary; // @[ArraySARA.scala 93:31]
  assign io_out_c_bypass_1_2_data = out_c_regNext_2_data; // @[ArraySARA.scala 93:31]
  assign io_out_c_bypass_1_2_is_stationary = out_c_regNext_2_is_stationary; // @[ArraySARA.scala 93:31]
  assign io_out_c_bypass_1_3_data = out_c_regNext_3_data; // @[ArraySARA.scala 93:31]
  assign io_out_c_bypass_1_3_is_stationary = out_c_regNext_3_is_stationary; // @[ArraySARA.scala 93:31]
  assign io_out_r_bypass_0_0_data = io_in_r_bypass_regNext_0_0_data; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_0_0_load_store = io_in_r_bypass_regNext_0_0_load_store; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_0_0_df_is_ws = io_in_r_bypass_regNext_0_0_df_is_ws; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_0_0_stall = io_in_r_bypass_regNext_0_0_stall; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_0_1_data = io_in_r_bypass_regNext_0_1_data; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_0_1_load_store = io_in_r_bypass_regNext_0_1_load_store; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_0_1_df_is_ws = io_in_r_bypass_regNext_0_1_df_is_ws; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_0_1_stall = io_in_r_bypass_regNext_0_1_stall; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_0_2_data = io_in_r_bypass_regNext_0_2_data; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_0_2_load_store = io_in_r_bypass_regNext_0_2_load_store; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_0_2_df_is_ws = io_in_r_bypass_regNext_0_2_df_is_ws; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_0_2_stall = io_in_r_bypass_regNext_0_2_stall; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_0_3_data = io_in_r_bypass_regNext_0_3_data; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_0_3_load_store = io_in_r_bypass_regNext_0_3_load_store; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_0_3_df_is_ws = io_in_r_bypass_regNext_0_3_df_is_ws; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_0_3_stall = io_in_r_bypass_regNext_0_3_stall; // @[ArraySARA.scala 97:26]
  assign io_out_c_bypass_0_0_data = io_in_c_bypass_regNext_0_0_data; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_0_0_is_stationary = io_in_c_bypass_regNext_0_0_is_stationary; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_0_1_data = io_in_c_bypass_regNext_0_1_data; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_0_1_is_stationary = io_in_c_bypass_regNext_0_1_is_stationary; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_0_2_data = io_in_c_bypass_regNext_0_2_data; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_0_2_is_stationary = io_in_c_bypass_regNext_0_2_is_stationary; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_0_3_data = io_in_c_bypass_regNext_0_3_data; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_0_3_is_stationary = io_in_c_bypass_regNext_0_3_is_stationary; // @[ArraySARA.scala 101:26]
  assign io_out_r_input_from_bypass_0 = io_in_r_input_from_bypass_regNext_0; // @[ArraySARA.scala 103:30]
  assign io_out_r_input_from_bypass_1 = io_in_r_input_from_bypass_regNext_1; // @[ArraySARA.scala 103:30]
  assign io_out_c_input_from_bypass_0 = io_in_c_input_from_bypass_regNext_0; // @[ArraySARA.scala 104:30]
  assign io_out_c_input_from_bypass_1 = io_in_c_input_from_bypass_regNext_1; // @[ArraySARA.scala 104:30]
  always @(posedge clk) begin
    out_r_regNext_0_data <= out_r_0_data; // @[Reg.scala 39:30]
    out_r_regNext_0_load_store <= out_r_0_load_store; // @[Reg.scala 39:30]
    out_r_regNext_0_df_is_ws <= out_r_0_df_is_ws; // @[Reg.scala 39:30]
    out_r_regNext_0_stall <= out_r_0_stall; // @[Reg.scala 39:30]
    out_r_regNext_1_data <= out_r_1_data; // @[Reg.scala 39:30]
    out_r_regNext_1_load_store <= out_r_1_load_store; // @[Reg.scala 39:30]
    out_r_regNext_1_df_is_ws <= out_r_1_df_is_ws; // @[Reg.scala 39:30]
    out_r_regNext_1_stall <= out_r_1_stall; // @[Reg.scala 39:30]
    out_r_regNext_2_data <= out_r_2_data; // @[Reg.scala 39:30]
    out_r_regNext_2_load_store <= out_r_2_load_store; // @[Reg.scala 39:30]
    out_r_regNext_2_df_is_ws <= out_r_2_df_is_ws; // @[Reg.scala 39:30]
    out_r_regNext_2_stall <= out_r_2_stall; // @[Reg.scala 39:30]
    out_r_regNext_3_data <= out_r_3_data; // @[Reg.scala 39:30]
    out_r_regNext_3_load_store <= out_r_3_load_store; // @[Reg.scala 39:30]
    out_r_regNext_3_df_is_ws <= out_r_3_df_is_ws; // @[Reg.scala 39:30]
    out_r_regNext_3_stall <= out_r_3_stall; // @[Reg.scala 39:30]
    out_c_regNext_0_data <= out_c_0_data; // @[Reg.scala 39:30]
    out_c_regNext_0_is_stationary <= out_c_0_is_stationary; // @[Reg.scala 39:30]
    out_c_regNext_1_data <= out_c_1_data; // @[Reg.scala 39:30]
    out_c_regNext_1_is_stationary <= out_c_1_is_stationary; // @[Reg.scala 39:30]
    out_c_regNext_2_data <= out_c_2_data; // @[Reg.scala 39:30]
    out_c_regNext_2_is_stationary <= out_c_2_is_stationary; // @[Reg.scala 39:30]
    out_c_regNext_3_data <= out_c_3_data; // @[Reg.scala 39:30]
    out_c_regNext_3_is_stationary <= out_c_3_is_stationary; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_0_data <= io_in_r_bypass_0_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_0_load_store <= io_in_r_bypass_0_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_0_df_is_ws <= io_in_r_bypass_0_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_0_stall <= io_in_r_bypass_0_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_1_data <= io_in_r_bypass_0_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_1_load_store <= io_in_r_bypass_0_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_1_df_is_ws <= io_in_r_bypass_0_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_1_stall <= io_in_r_bypass_0_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_2_data <= io_in_r_bypass_0_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_2_load_store <= io_in_r_bypass_0_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_2_df_is_ws <= io_in_r_bypass_0_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_2_stall <= io_in_r_bypass_0_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_3_data <= io_in_r_bypass_0_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_3_load_store <= io_in_r_bypass_0_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_3_df_is_ws <= io_in_r_bypass_0_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_3_stall <= io_in_r_bypass_0_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_0_data <= io_in_r_bypass_1_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_0_load_store <= io_in_r_bypass_1_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_0_df_is_ws <= io_in_r_bypass_1_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_0_stall <= io_in_r_bypass_1_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_1_data <= io_in_r_bypass_1_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_1_load_store <= io_in_r_bypass_1_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_1_df_is_ws <= io_in_r_bypass_1_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_1_stall <= io_in_r_bypass_1_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_2_data <= io_in_r_bypass_1_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_2_load_store <= io_in_r_bypass_1_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_2_df_is_ws <= io_in_r_bypass_1_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_2_stall <= io_in_r_bypass_1_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_3_data <= io_in_r_bypass_1_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_3_load_store <= io_in_r_bypass_1_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_3_df_is_ws <= io_in_r_bypass_1_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_3_stall <= io_in_r_bypass_1_3_stall; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_0_data <= io_in_c_bypass_0_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_0_is_stationary <= io_in_c_bypass_0_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_1_data <= io_in_c_bypass_0_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_1_is_stationary <= io_in_c_bypass_0_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_2_data <= io_in_c_bypass_0_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_2_is_stationary <= io_in_c_bypass_0_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_3_data <= io_in_c_bypass_0_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_3_is_stationary <= io_in_c_bypass_0_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_0_data <= io_in_c_bypass_1_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_0_is_stationary <= io_in_c_bypass_1_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_1_data <= io_in_c_bypass_1_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_1_is_stationary <= io_in_c_bypass_1_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_2_data <= io_in_c_bypass_1_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_2_is_stationary <= io_in_c_bypass_1_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_3_data <= io_in_c_bypass_1_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_3_is_stationary <= io_in_c_bypass_1_3_is_stationary; // @[Reg.scala 39:30]
    io_in_r_input_from_bypass_regNext_0 <= io_in_r_input_from_bypass_0; // @[Reg.scala 39:30]
    io_in_r_input_from_bypass_regNext_1 <= io_in_r_input_from_bypass_1; // @[Reg.scala 39:30]
    io_in_c_input_from_bypass_regNext_0 <= io_in_c_input_from_bypass_0; // @[Reg.scala 39:30]
    io_in_c_input_from_bypass_regNext_1 <= io_in_c_input_from_bypass_1; // @[Reg.scala 39:30]
  end


endmodule

module CellSARA_1 (
  input      [15:0]   io_in_r_data_0_data,
  input               io_in_r_data_0_load_store,
  input               io_in_r_data_0_df_is_ws,
  input               io_in_r_data_0_stall,
  input      [15:0]   io_in_r_data_1_data,
  input               io_in_r_data_1_load_store,
  input               io_in_r_data_1_df_is_ws,
  input               io_in_r_data_1_stall,
  input      [15:0]   io_in_r_data_2_data,
  input               io_in_r_data_2_load_store,
  input               io_in_r_data_2_df_is_ws,
  input               io_in_r_data_2_stall,
  input      [15:0]   io_in_r_data_3_data,
  input               io_in_r_data_3_load_store,
  input               io_in_r_data_3_df_is_ws,
  input               io_in_r_data_3_stall,
  input      [15:0]   io_in_r_bypass_0_0_data,
  input               io_in_r_bypass_0_0_load_store,
  input               io_in_r_bypass_0_0_df_is_ws,
  input               io_in_r_bypass_0_0_stall,
  input      [15:0]   io_in_r_bypass_0_1_data,
  input               io_in_r_bypass_0_1_load_store,
  input               io_in_r_bypass_0_1_df_is_ws,
  input               io_in_r_bypass_0_1_stall,
  input      [15:0]   io_in_r_bypass_0_2_data,
  input               io_in_r_bypass_0_2_load_store,
  input               io_in_r_bypass_0_2_df_is_ws,
  input               io_in_r_bypass_0_2_stall,
  input      [15:0]   io_in_r_bypass_0_3_data,
  input               io_in_r_bypass_0_3_load_store,
  input               io_in_r_bypass_0_3_df_is_ws,
  input               io_in_r_bypass_0_3_stall,
  input      [15:0]   io_in_r_bypass_1_0_data,
  input               io_in_r_bypass_1_0_load_store,
  input               io_in_r_bypass_1_0_df_is_ws,
  input               io_in_r_bypass_1_0_stall,
  input      [15:0]   io_in_r_bypass_1_1_data,
  input               io_in_r_bypass_1_1_load_store,
  input               io_in_r_bypass_1_1_df_is_ws,
  input               io_in_r_bypass_1_1_stall,
  input      [15:0]   io_in_r_bypass_1_2_data,
  input               io_in_r_bypass_1_2_load_store,
  input               io_in_r_bypass_1_2_df_is_ws,
  input               io_in_r_bypass_1_2_stall,
  input      [15:0]   io_in_r_bypass_1_3_data,
  input               io_in_r_bypass_1_3_load_store,
  input               io_in_r_bypass_1_3_df_is_ws,
  input               io_in_r_bypass_1_3_stall,
  input               io_in_r_input_from_bypass_0,
  input               io_in_r_input_from_bypass_1,
  output     [15:0]   io_out_r_data_0_data,
  output              io_out_r_data_0_load_store,
  output              io_out_r_data_0_df_is_ws,
  output              io_out_r_data_0_stall,
  output     [15:0]   io_out_r_data_1_data,
  output              io_out_r_data_1_load_store,
  output              io_out_r_data_1_df_is_ws,
  output              io_out_r_data_1_stall,
  output     [15:0]   io_out_r_data_2_data,
  output              io_out_r_data_2_load_store,
  output              io_out_r_data_2_df_is_ws,
  output              io_out_r_data_2_stall,
  output     [15:0]   io_out_r_data_3_data,
  output              io_out_r_data_3_load_store,
  output              io_out_r_data_3_df_is_ws,
  output              io_out_r_data_3_stall,
  output     [15:0]   io_out_r_bypass_0_0_data,
  output              io_out_r_bypass_0_0_load_store,
  output              io_out_r_bypass_0_0_df_is_ws,
  output              io_out_r_bypass_0_0_stall,
  output     [15:0]   io_out_r_bypass_0_1_data,
  output              io_out_r_bypass_0_1_load_store,
  output              io_out_r_bypass_0_1_df_is_ws,
  output              io_out_r_bypass_0_1_stall,
  output     [15:0]   io_out_r_bypass_0_2_data,
  output              io_out_r_bypass_0_2_load_store,
  output              io_out_r_bypass_0_2_df_is_ws,
  output              io_out_r_bypass_0_2_stall,
  output     [15:0]   io_out_r_bypass_0_3_data,
  output              io_out_r_bypass_0_3_load_store,
  output              io_out_r_bypass_0_3_df_is_ws,
  output              io_out_r_bypass_0_3_stall,
  output     [15:0]   io_out_r_bypass_1_0_data,
  output              io_out_r_bypass_1_0_load_store,
  output              io_out_r_bypass_1_0_df_is_ws,
  output              io_out_r_bypass_1_0_stall,
  output     [15:0]   io_out_r_bypass_1_1_data,
  output              io_out_r_bypass_1_1_load_store,
  output              io_out_r_bypass_1_1_df_is_ws,
  output              io_out_r_bypass_1_1_stall,
  output     [15:0]   io_out_r_bypass_1_2_data,
  output              io_out_r_bypass_1_2_load_store,
  output              io_out_r_bypass_1_2_df_is_ws,
  output              io_out_r_bypass_1_2_stall,
  output     [15:0]   io_out_r_bypass_1_3_data,
  output              io_out_r_bypass_1_3_load_store,
  output              io_out_r_bypass_1_3_df_is_ws,
  output              io_out_r_bypass_1_3_stall,
  output              io_out_r_input_from_bypass_0,
  output              io_out_r_input_from_bypass_1,
  input      [15:0]   io_in_c_data_0_data,
  input               io_in_c_data_0_is_stationary,
  input      [15:0]   io_in_c_data_1_data,
  input               io_in_c_data_1_is_stationary,
  input      [15:0]   io_in_c_data_2_data,
  input               io_in_c_data_2_is_stationary,
  input      [15:0]   io_in_c_data_3_data,
  input               io_in_c_data_3_is_stationary,
  input      [15:0]   io_in_c_bypass_0_0_data,
  input               io_in_c_bypass_0_0_is_stationary,
  input      [15:0]   io_in_c_bypass_0_1_data,
  input               io_in_c_bypass_0_1_is_stationary,
  input      [15:0]   io_in_c_bypass_0_2_data,
  input               io_in_c_bypass_0_2_is_stationary,
  input      [15:0]   io_in_c_bypass_0_3_data,
  input               io_in_c_bypass_0_3_is_stationary,
  input      [15:0]   io_in_c_bypass_1_0_data,
  input               io_in_c_bypass_1_0_is_stationary,
  input      [15:0]   io_in_c_bypass_1_1_data,
  input               io_in_c_bypass_1_1_is_stationary,
  input      [15:0]   io_in_c_bypass_1_2_data,
  input               io_in_c_bypass_1_2_is_stationary,
  input      [15:0]   io_in_c_bypass_1_3_data,
  input               io_in_c_bypass_1_3_is_stationary,
  input               io_in_c_input_from_bypass_0,
  input               io_in_c_input_from_bypass_1,
  output     [15:0]   io_out_c_data_0_data,
  output              io_out_c_data_0_is_stationary,
  output     [15:0]   io_out_c_data_1_data,
  output              io_out_c_data_1_is_stationary,
  output     [15:0]   io_out_c_data_2_data,
  output              io_out_c_data_2_is_stationary,
  output     [15:0]   io_out_c_data_3_data,
  output              io_out_c_data_3_is_stationary,
  output     [15:0]   io_out_c_bypass_0_0_data,
  output              io_out_c_bypass_0_0_is_stationary,
  output     [15:0]   io_out_c_bypass_0_1_data,
  output              io_out_c_bypass_0_1_is_stationary,
  output     [15:0]   io_out_c_bypass_0_2_data,
  output              io_out_c_bypass_0_2_is_stationary,
  output     [15:0]   io_out_c_bypass_0_3_data,
  output              io_out_c_bypass_0_3_is_stationary,
  output     [15:0]   io_out_c_bypass_1_0_data,
  output              io_out_c_bypass_1_0_is_stationary,
  output     [15:0]   io_out_c_bypass_1_1_data,
  output              io_out_c_bypass_1_1_is_stationary,
  output     [15:0]   io_out_c_bypass_1_2_data,
  output              io_out_c_bypass_1_2_is_stationary,
  output     [15:0]   io_out_c_bypass_1_3_data,
  output              io_out_c_bypass_1_3_is_stationary,
  output              io_out_c_input_from_bypass_0,
  output              io_out_c_input_from_bypass_1,
  input               clk,
  input               reset
);

  wire       [15:0]   pes_0_0_io_out_r_data;
  wire                pes_0_0_io_out_r_load_store;
  wire                pes_0_0_io_out_r_df_is_ws;
  wire                pes_0_0_io_out_r_stall;
  wire       [15:0]   pes_0_0_io_out_c_data;
  wire                pes_0_0_io_out_c_is_stationary;
  wire       [15:0]   pes_0_1_io_out_r_data;
  wire                pes_0_1_io_out_r_load_store;
  wire                pes_0_1_io_out_r_df_is_ws;
  wire                pes_0_1_io_out_r_stall;
  wire       [15:0]   pes_0_1_io_out_c_data;
  wire                pes_0_1_io_out_c_is_stationary;
  wire       [15:0]   pes_0_2_io_out_r_data;
  wire                pes_0_2_io_out_r_load_store;
  wire                pes_0_2_io_out_r_df_is_ws;
  wire                pes_0_2_io_out_r_stall;
  wire       [15:0]   pes_0_2_io_out_c_data;
  wire                pes_0_2_io_out_c_is_stationary;
  wire       [15:0]   pes_0_3_io_out_r_data;
  wire                pes_0_3_io_out_r_load_store;
  wire                pes_0_3_io_out_r_df_is_ws;
  wire                pes_0_3_io_out_r_stall;
  wire       [15:0]   pes_0_3_io_out_c_data;
  wire                pes_0_3_io_out_c_is_stationary;
  wire       [15:0]   pes_1_0_io_out_r_data;
  wire                pes_1_0_io_out_r_load_store;
  wire                pes_1_0_io_out_r_df_is_ws;
  wire                pes_1_0_io_out_r_stall;
  wire       [15:0]   pes_1_0_io_out_c_data;
  wire                pes_1_0_io_out_c_is_stationary;
  wire       [15:0]   pes_1_1_io_out_r_data;
  wire                pes_1_1_io_out_r_load_store;
  wire                pes_1_1_io_out_r_df_is_ws;
  wire                pes_1_1_io_out_r_stall;
  wire       [15:0]   pes_1_1_io_out_c_data;
  wire                pes_1_1_io_out_c_is_stationary;
  wire       [15:0]   pes_1_2_io_out_r_data;
  wire                pes_1_2_io_out_r_load_store;
  wire                pes_1_2_io_out_r_df_is_ws;
  wire                pes_1_2_io_out_r_stall;
  wire       [15:0]   pes_1_2_io_out_c_data;
  wire                pes_1_2_io_out_c_is_stationary;
  wire       [15:0]   pes_1_3_io_out_r_data;
  wire                pes_1_3_io_out_r_load_store;
  wire                pes_1_3_io_out_r_df_is_ws;
  wire                pes_1_3_io_out_r_stall;
  wire       [15:0]   pes_1_3_io_out_c_data;
  wire                pes_1_3_io_out_c_is_stationary;
  wire       [15:0]   pes_2_0_io_out_r_data;
  wire                pes_2_0_io_out_r_load_store;
  wire                pes_2_0_io_out_r_df_is_ws;
  wire                pes_2_0_io_out_r_stall;
  wire       [15:0]   pes_2_0_io_out_c_data;
  wire                pes_2_0_io_out_c_is_stationary;
  wire       [15:0]   pes_2_1_io_out_r_data;
  wire                pes_2_1_io_out_r_load_store;
  wire                pes_2_1_io_out_r_df_is_ws;
  wire                pes_2_1_io_out_r_stall;
  wire       [15:0]   pes_2_1_io_out_c_data;
  wire                pes_2_1_io_out_c_is_stationary;
  wire       [15:0]   pes_2_2_io_out_r_data;
  wire                pes_2_2_io_out_r_load_store;
  wire                pes_2_2_io_out_r_df_is_ws;
  wire                pes_2_2_io_out_r_stall;
  wire       [15:0]   pes_2_2_io_out_c_data;
  wire                pes_2_2_io_out_c_is_stationary;
  wire       [15:0]   pes_2_3_io_out_r_data;
  wire                pes_2_3_io_out_r_load_store;
  wire                pes_2_3_io_out_r_df_is_ws;
  wire                pes_2_3_io_out_r_stall;
  wire       [15:0]   pes_2_3_io_out_c_data;
  wire                pes_2_3_io_out_c_is_stationary;
  wire       [15:0]   pes_3_0_io_out_r_data;
  wire                pes_3_0_io_out_r_load_store;
  wire                pes_3_0_io_out_r_df_is_ws;
  wire                pes_3_0_io_out_r_stall;
  wire       [15:0]   pes_3_0_io_out_c_data;
  wire                pes_3_0_io_out_c_is_stationary;
  wire       [15:0]   pes_3_1_io_out_r_data;
  wire                pes_3_1_io_out_r_load_store;
  wire                pes_3_1_io_out_r_df_is_ws;
  wire                pes_3_1_io_out_r_stall;
  wire       [15:0]   pes_3_1_io_out_c_data;
  wire                pes_3_1_io_out_c_is_stationary;
  wire       [15:0]   pes_3_2_io_out_r_data;
  wire                pes_3_2_io_out_r_load_store;
  wire                pes_3_2_io_out_r_df_is_ws;
  wire                pes_3_2_io_out_r_stall;
  wire       [15:0]   pes_3_2_io_out_c_data;
  wire                pes_3_2_io_out_c_is_stationary;
  wire       [15:0]   pes_3_3_io_out_r_data;
  wire                pes_3_3_io_out_r_load_store;
  wire                pes_3_3_io_out_r_df_is_ws;
  wire                pes_3_3_io_out_r_stall;
  wire       [15:0]   pes_3_3_io_out_c_data;
  wire                pes_3_3_io_out_c_is_stationary;
  wire       [15:0]   in_r_0_data;
  wire                in_r_0_load_store;
  wire                in_r_0_df_is_ws;
  wire                in_r_0_stall;
  wire       [15:0]   in_r_1_data;
  wire                in_r_1_load_store;
  wire                in_r_1_df_is_ws;
  wire                in_r_1_stall;
  wire       [15:0]   in_r_2_data;
  wire                in_r_2_load_store;
  wire                in_r_2_df_is_ws;
  wire                in_r_2_stall;
  wire       [15:0]   in_r_3_data;
  wire                in_r_3_load_store;
  wire                in_r_3_df_is_ws;
  wire                in_r_3_stall;
  wire       [15:0]   in_c_0_data;
  wire                in_c_0_is_stationary;
  wire       [15:0]   in_c_1_data;
  wire                in_c_1_is_stationary;
  wire       [15:0]   in_c_2_data;
  wire                in_c_2_is_stationary;
  wire       [15:0]   in_c_3_data;
  wire                in_c_3_is_stationary;
  wire       [15:0]   out_r_0_data;
  wire                out_r_0_load_store;
  wire                out_r_0_df_is_ws;
  wire                out_r_0_stall;
  wire       [15:0]   out_r_1_data;
  wire                out_r_1_load_store;
  wire                out_r_1_df_is_ws;
  wire                out_r_1_stall;
  wire       [15:0]   out_r_2_data;
  wire                out_r_2_load_store;
  wire                out_r_2_df_is_ws;
  wire                out_r_2_stall;
  wire       [15:0]   out_r_3_data;
  wire                out_r_3_load_store;
  wire                out_r_3_df_is_ws;
  wire                out_r_3_stall;
  wire       [15:0]   out_c_0_data;
  wire                out_c_0_is_stationary;
  wire       [15:0]   out_c_1_data;
  wire                out_c_1_is_stationary;
  wire       [15:0]   out_c_2_data;
  wire                out_c_2_is_stationary;
  wire       [15:0]   out_c_3_data;
  wire                out_c_3_is_stationary;
  reg        [15:0]   out_r_regNext_0_data;
  reg                 out_r_regNext_0_load_store;
  reg                 out_r_regNext_0_df_is_ws;
  reg                 out_r_regNext_0_stall;
  reg        [15:0]   out_r_regNext_1_data;
  reg                 out_r_regNext_1_load_store;
  reg                 out_r_regNext_1_df_is_ws;
  reg                 out_r_regNext_1_stall;
  reg        [15:0]   out_r_regNext_2_data;
  reg                 out_r_regNext_2_load_store;
  reg                 out_r_regNext_2_df_is_ws;
  reg                 out_r_regNext_2_stall;
  reg        [15:0]   out_r_regNext_3_data;
  reg                 out_r_regNext_3_load_store;
  reg                 out_r_regNext_3_df_is_ws;
  reg                 out_r_regNext_3_stall;
  reg        [15:0]   out_c_regNext_0_data;
  reg                 out_c_regNext_0_is_stationary;
  reg        [15:0]   out_c_regNext_1_data;
  reg                 out_c_regNext_1_is_stationary;
  reg        [15:0]   out_c_regNext_2_data;
  reg                 out_c_regNext_2_is_stationary;
  reg        [15:0]   out_c_regNext_3_data;
  reg                 out_c_regNext_3_is_stationary;
  reg        [15:0]   io_in_r_bypass_regNext_0_0_data;
  reg                 io_in_r_bypass_regNext_0_0_load_store;
  reg                 io_in_r_bypass_regNext_0_0_df_is_ws;
  reg                 io_in_r_bypass_regNext_0_0_stall;
  reg        [15:0]   io_in_r_bypass_regNext_0_1_data;
  reg                 io_in_r_bypass_regNext_0_1_load_store;
  reg                 io_in_r_bypass_regNext_0_1_df_is_ws;
  reg                 io_in_r_bypass_regNext_0_1_stall;
  reg        [15:0]   io_in_r_bypass_regNext_0_2_data;
  reg                 io_in_r_bypass_regNext_0_2_load_store;
  reg                 io_in_r_bypass_regNext_0_2_df_is_ws;
  reg                 io_in_r_bypass_regNext_0_2_stall;
  reg        [15:0]   io_in_r_bypass_regNext_0_3_data;
  reg                 io_in_r_bypass_regNext_0_3_load_store;
  reg                 io_in_r_bypass_regNext_0_3_df_is_ws;
  reg                 io_in_r_bypass_regNext_0_3_stall;
  reg        [15:0]   io_in_r_bypass_regNext_1_0_data;
  reg                 io_in_r_bypass_regNext_1_0_load_store;
  reg                 io_in_r_bypass_regNext_1_0_df_is_ws;
  reg                 io_in_r_bypass_regNext_1_0_stall;
  reg        [15:0]   io_in_r_bypass_regNext_1_1_data;
  reg                 io_in_r_bypass_regNext_1_1_load_store;
  reg                 io_in_r_bypass_regNext_1_1_df_is_ws;
  reg                 io_in_r_bypass_regNext_1_1_stall;
  reg        [15:0]   io_in_r_bypass_regNext_1_2_data;
  reg                 io_in_r_bypass_regNext_1_2_load_store;
  reg                 io_in_r_bypass_regNext_1_2_df_is_ws;
  reg                 io_in_r_bypass_regNext_1_2_stall;
  reg        [15:0]   io_in_r_bypass_regNext_1_3_data;
  reg                 io_in_r_bypass_regNext_1_3_load_store;
  reg                 io_in_r_bypass_regNext_1_3_df_is_ws;
  reg                 io_in_r_bypass_regNext_1_3_stall;
  reg        [15:0]   io_in_c_bypass_regNext_0_0_data;
  reg                 io_in_c_bypass_regNext_0_0_is_stationary;
  reg        [15:0]   io_in_c_bypass_regNext_0_1_data;
  reg                 io_in_c_bypass_regNext_0_1_is_stationary;
  reg        [15:0]   io_in_c_bypass_regNext_0_2_data;
  reg                 io_in_c_bypass_regNext_0_2_is_stationary;
  reg        [15:0]   io_in_c_bypass_regNext_0_3_data;
  reg                 io_in_c_bypass_regNext_0_3_is_stationary;
  reg        [15:0]   io_in_c_bypass_regNext_1_0_data;
  reg                 io_in_c_bypass_regNext_1_0_is_stationary;
  reg        [15:0]   io_in_c_bypass_regNext_1_1_data;
  reg                 io_in_c_bypass_regNext_1_1_is_stationary;
  reg        [15:0]   io_in_c_bypass_regNext_1_2_data;
  reg                 io_in_c_bypass_regNext_1_2_is_stationary;
  reg        [15:0]   io_in_c_bypass_regNext_1_3_data;
  reg                 io_in_c_bypass_regNext_1_3_is_stationary;
  reg                 io_in_r_input_from_bypass_regNext_0;
  reg                 io_in_r_input_from_bypass_regNext_1;
  reg                 io_in_c_input_from_bypass_regNext_0;
  reg                 io_in_c_input_from_bypass_regNext_1;

  PEWSOS_127 pes_0_0 (
    .io_in_r_data           (in_r_0_data[15:0]             ), //i
    .io_in_r_load_store     (in_r_0_load_store             ), //i
    .io_in_r_df_is_ws       (in_r_0_df_is_ws               ), //i
    .io_in_r_stall          (in_r_0_stall                  ), //i
    .io_out_r_data          (pes_0_0_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pes_0_0_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pes_0_0_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pes_0_0_io_out_r_stall        ), //o
    .io_in_c_data           (in_c_0_data[15:0]             ), //i
    .io_in_c_is_stationary  (in_c_0_is_stationary          ), //i
    .io_out_c_data          (pes_0_0_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pes_0_0_io_out_c_is_stationary), //o
    .clk                    (clk                           ), //i
    .reset                  (reset                         )  //i
  );
  PEWSOS_127 pes_0_1 (
    .io_in_r_data           (pes_0_0_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pes_0_0_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pes_0_0_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pes_0_0_io_out_r_stall        ), //i
    .io_out_r_data          (pes_0_1_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pes_0_1_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pes_0_1_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pes_0_1_io_out_r_stall        ), //o
    .io_in_c_data           (in_c_1_data[15:0]             ), //i
    .io_in_c_is_stationary  (in_c_1_is_stationary          ), //i
    .io_out_c_data          (pes_0_1_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pes_0_1_io_out_c_is_stationary), //o
    .clk                    (clk                           ), //i
    .reset                  (reset                         )  //i
  );
  PEWSOS_127 pes_0_2 (
    .io_in_r_data           (pes_0_1_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pes_0_1_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pes_0_1_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pes_0_1_io_out_r_stall        ), //i
    .io_out_r_data          (pes_0_2_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pes_0_2_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pes_0_2_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pes_0_2_io_out_r_stall        ), //o
    .io_in_c_data           (in_c_2_data[15:0]             ), //i
    .io_in_c_is_stationary  (in_c_2_is_stationary          ), //i
    .io_out_c_data          (pes_0_2_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pes_0_2_io_out_c_is_stationary), //o
    .clk                    (clk                           ), //i
    .reset                  (reset                         )  //i
  );
  PEWSOS_127 pes_0_3 (
    .io_in_r_data           (pes_0_2_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pes_0_2_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pes_0_2_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pes_0_2_io_out_r_stall        ), //i
    .io_out_r_data          (pes_0_3_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pes_0_3_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pes_0_3_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pes_0_3_io_out_r_stall        ), //o
    .io_in_c_data           (in_c_3_data[15:0]             ), //i
    .io_in_c_is_stationary  (in_c_3_is_stationary          ), //i
    .io_out_c_data          (pes_0_3_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pes_0_3_io_out_c_is_stationary), //o
    .clk                    (clk                           ), //i
    .reset                  (reset                         )  //i
  );
  PEWSOS_127 pes_1_0 (
    .io_in_r_data           (in_r_1_data[15:0]             ), //i
    .io_in_r_load_store     (in_r_1_load_store             ), //i
    .io_in_r_df_is_ws       (in_r_1_df_is_ws               ), //i
    .io_in_r_stall          (in_r_1_stall                  ), //i
    .io_out_r_data          (pes_1_0_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pes_1_0_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pes_1_0_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pes_1_0_io_out_r_stall        ), //o
    .io_in_c_data           (pes_0_0_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pes_0_0_io_out_c_is_stationary), //i
    .io_out_c_data          (pes_1_0_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pes_1_0_io_out_c_is_stationary), //o
    .clk                    (clk                           ), //i
    .reset                  (reset                         )  //i
  );
  PEWSOS_127 pes_1_1 (
    .io_in_r_data           (pes_1_0_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pes_1_0_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pes_1_0_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pes_1_0_io_out_r_stall        ), //i
    .io_out_r_data          (pes_1_1_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pes_1_1_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pes_1_1_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pes_1_1_io_out_r_stall        ), //o
    .io_in_c_data           (pes_0_1_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pes_0_1_io_out_c_is_stationary), //i
    .io_out_c_data          (pes_1_1_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pes_1_1_io_out_c_is_stationary), //o
    .clk                    (clk                           ), //i
    .reset                  (reset                         )  //i
  );
  PEWSOS_127 pes_1_2 (
    .io_in_r_data           (pes_1_1_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pes_1_1_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pes_1_1_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pes_1_1_io_out_r_stall        ), //i
    .io_out_r_data          (pes_1_2_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pes_1_2_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pes_1_2_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pes_1_2_io_out_r_stall        ), //o
    .io_in_c_data           (pes_0_2_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pes_0_2_io_out_c_is_stationary), //i
    .io_out_c_data          (pes_1_2_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pes_1_2_io_out_c_is_stationary), //o
    .clk                    (clk                           ), //i
    .reset                  (reset                         )  //i
  );
  PEWSOS_127 pes_1_3 (
    .io_in_r_data           (pes_1_2_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pes_1_2_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pes_1_2_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pes_1_2_io_out_r_stall        ), //i
    .io_out_r_data          (pes_1_3_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pes_1_3_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pes_1_3_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pes_1_3_io_out_r_stall        ), //o
    .io_in_c_data           (pes_0_3_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pes_0_3_io_out_c_is_stationary), //i
    .io_out_c_data          (pes_1_3_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pes_1_3_io_out_c_is_stationary), //o
    .clk                    (clk                           ), //i
    .reset                  (reset                         )  //i
  );
  PEWSOS_127 pes_2_0 (
    .io_in_r_data           (in_r_2_data[15:0]             ), //i
    .io_in_r_load_store     (in_r_2_load_store             ), //i
    .io_in_r_df_is_ws       (in_r_2_df_is_ws               ), //i
    .io_in_r_stall          (in_r_2_stall                  ), //i
    .io_out_r_data          (pes_2_0_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pes_2_0_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pes_2_0_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pes_2_0_io_out_r_stall        ), //o
    .io_in_c_data           (pes_1_0_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pes_1_0_io_out_c_is_stationary), //i
    .io_out_c_data          (pes_2_0_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pes_2_0_io_out_c_is_stationary), //o
    .clk                    (clk                           ), //i
    .reset                  (reset                         )  //i
  );
  PEWSOS_127 pes_2_1 (
    .io_in_r_data           (pes_2_0_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pes_2_0_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pes_2_0_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pes_2_0_io_out_r_stall        ), //i
    .io_out_r_data          (pes_2_1_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pes_2_1_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pes_2_1_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pes_2_1_io_out_r_stall        ), //o
    .io_in_c_data           (pes_1_1_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pes_1_1_io_out_c_is_stationary), //i
    .io_out_c_data          (pes_2_1_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pes_2_1_io_out_c_is_stationary), //o
    .clk                    (clk                           ), //i
    .reset                  (reset                         )  //i
  );
  PEWSOS_127 pes_2_2 (
    .io_in_r_data           (pes_2_1_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pes_2_1_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pes_2_1_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pes_2_1_io_out_r_stall        ), //i
    .io_out_r_data          (pes_2_2_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pes_2_2_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pes_2_2_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pes_2_2_io_out_r_stall        ), //o
    .io_in_c_data           (pes_1_2_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pes_1_2_io_out_c_is_stationary), //i
    .io_out_c_data          (pes_2_2_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pes_2_2_io_out_c_is_stationary), //o
    .clk                    (clk                           ), //i
    .reset                  (reset                         )  //i
  );
  PEWSOS_127 pes_2_3 (
    .io_in_r_data           (pes_2_2_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pes_2_2_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pes_2_2_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pes_2_2_io_out_r_stall        ), //i
    .io_out_r_data          (pes_2_3_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pes_2_3_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pes_2_3_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pes_2_3_io_out_r_stall        ), //o
    .io_in_c_data           (pes_1_3_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pes_1_3_io_out_c_is_stationary), //i
    .io_out_c_data          (pes_2_3_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pes_2_3_io_out_c_is_stationary), //o
    .clk                    (clk                           ), //i
    .reset                  (reset                         )  //i
  );
  PEWSOS_127 pes_3_0 (
    .io_in_r_data           (in_r_3_data[15:0]             ), //i
    .io_in_r_load_store     (in_r_3_load_store             ), //i
    .io_in_r_df_is_ws       (in_r_3_df_is_ws               ), //i
    .io_in_r_stall          (in_r_3_stall                  ), //i
    .io_out_r_data          (pes_3_0_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pes_3_0_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pes_3_0_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pes_3_0_io_out_r_stall        ), //o
    .io_in_c_data           (pes_2_0_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pes_2_0_io_out_c_is_stationary), //i
    .io_out_c_data          (pes_3_0_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pes_3_0_io_out_c_is_stationary), //o
    .clk                    (clk                           ), //i
    .reset                  (reset                         )  //i
  );
  PEWSOS_127 pes_3_1 (
    .io_in_r_data           (pes_3_0_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pes_3_0_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pes_3_0_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pes_3_0_io_out_r_stall        ), //i
    .io_out_r_data          (pes_3_1_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pes_3_1_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pes_3_1_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pes_3_1_io_out_r_stall        ), //o
    .io_in_c_data           (pes_2_1_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pes_2_1_io_out_c_is_stationary), //i
    .io_out_c_data          (pes_3_1_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pes_3_1_io_out_c_is_stationary), //o
    .clk                    (clk                           ), //i
    .reset                  (reset                         )  //i
  );
  PEWSOS_127 pes_3_2 (
    .io_in_r_data           (pes_3_1_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pes_3_1_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pes_3_1_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pes_3_1_io_out_r_stall        ), //i
    .io_out_r_data          (pes_3_2_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pes_3_2_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pes_3_2_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pes_3_2_io_out_r_stall        ), //o
    .io_in_c_data           (pes_2_2_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pes_2_2_io_out_c_is_stationary), //i
    .io_out_c_data          (pes_3_2_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pes_3_2_io_out_c_is_stationary), //o
    .clk                    (clk                           ), //i
    .reset                  (reset                         )  //i
  );
  PEWSOS_127 pes_3_3 (
    .io_in_r_data           (pes_3_2_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pes_3_2_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pes_3_2_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pes_3_2_io_out_r_stall        ), //i
    .io_out_r_data          (pes_3_3_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pes_3_3_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pes_3_3_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pes_3_3_io_out_r_stall        ), //o
    .io_in_c_data           (pes_2_3_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pes_2_3_io_out_c_is_stationary), //i
    .io_out_c_data          (pes_3_3_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pes_3_3_io_out_c_is_stationary), //o
    .clk                    (clk                           ), //i
    .reset                  (reset                         )  //i
  );
  assign in_r_0_data = (io_in_r_input_from_bypass_1 ? io_in_r_bypass_1_0_data : io_in_r_data_0_data); // @[Expression.scala 1420:25]
  assign in_r_0_load_store = (io_in_r_input_from_bypass_1 ? io_in_r_bypass_1_0_load_store : io_in_r_data_0_load_store); // @[Expression.scala 1420:25]
  assign in_r_0_df_is_ws = (io_in_r_input_from_bypass_1 ? io_in_r_bypass_1_0_df_is_ws : io_in_r_data_0_df_is_ws); // @[Expression.scala 1420:25]
  assign in_r_0_stall = (io_in_r_input_from_bypass_1 ? io_in_r_bypass_1_0_stall : io_in_r_data_0_stall); // @[Expression.scala 1420:25]
  assign in_r_1_data = (io_in_r_input_from_bypass_1 ? io_in_r_bypass_1_1_data : io_in_r_data_1_data); // @[Expression.scala 1420:25]
  assign in_r_1_load_store = (io_in_r_input_from_bypass_1 ? io_in_r_bypass_1_1_load_store : io_in_r_data_1_load_store); // @[Expression.scala 1420:25]
  assign in_r_1_df_is_ws = (io_in_r_input_from_bypass_1 ? io_in_r_bypass_1_1_df_is_ws : io_in_r_data_1_df_is_ws); // @[Expression.scala 1420:25]
  assign in_r_1_stall = (io_in_r_input_from_bypass_1 ? io_in_r_bypass_1_1_stall : io_in_r_data_1_stall); // @[Expression.scala 1420:25]
  assign in_r_2_data = (io_in_r_input_from_bypass_1 ? io_in_r_bypass_1_2_data : io_in_r_data_2_data); // @[Expression.scala 1420:25]
  assign in_r_2_load_store = (io_in_r_input_from_bypass_1 ? io_in_r_bypass_1_2_load_store : io_in_r_data_2_load_store); // @[Expression.scala 1420:25]
  assign in_r_2_df_is_ws = (io_in_r_input_from_bypass_1 ? io_in_r_bypass_1_2_df_is_ws : io_in_r_data_2_df_is_ws); // @[Expression.scala 1420:25]
  assign in_r_2_stall = (io_in_r_input_from_bypass_1 ? io_in_r_bypass_1_2_stall : io_in_r_data_2_stall); // @[Expression.scala 1420:25]
  assign in_r_3_data = (io_in_r_input_from_bypass_1 ? io_in_r_bypass_1_3_data : io_in_r_data_3_data); // @[Expression.scala 1420:25]
  assign in_r_3_load_store = (io_in_r_input_from_bypass_1 ? io_in_r_bypass_1_3_load_store : io_in_r_data_3_load_store); // @[Expression.scala 1420:25]
  assign in_r_3_df_is_ws = (io_in_r_input_from_bypass_1 ? io_in_r_bypass_1_3_df_is_ws : io_in_r_data_3_df_is_ws); // @[Expression.scala 1420:25]
  assign in_r_3_stall = (io_in_r_input_from_bypass_1 ? io_in_r_bypass_1_3_stall : io_in_r_data_3_stall); // @[Expression.scala 1420:25]
  assign in_c_0_data = (io_in_c_input_from_bypass_0 ? io_in_c_bypass_0_0_data : io_in_c_data_0_data); // @[Expression.scala 1420:25]
  assign in_c_0_is_stationary = (io_in_c_input_from_bypass_0 ? io_in_c_bypass_0_0_is_stationary : io_in_c_data_0_is_stationary); // @[Expression.scala 1420:25]
  assign in_c_1_data = (io_in_c_input_from_bypass_0 ? io_in_c_bypass_0_1_data : io_in_c_data_1_data); // @[Expression.scala 1420:25]
  assign in_c_1_is_stationary = (io_in_c_input_from_bypass_0 ? io_in_c_bypass_0_1_is_stationary : io_in_c_data_1_is_stationary); // @[Expression.scala 1420:25]
  assign in_c_2_data = (io_in_c_input_from_bypass_0 ? io_in_c_bypass_0_2_data : io_in_c_data_2_data); // @[Expression.scala 1420:25]
  assign in_c_2_is_stationary = (io_in_c_input_from_bypass_0 ? io_in_c_bypass_0_2_is_stationary : io_in_c_data_2_is_stationary); // @[Expression.scala 1420:25]
  assign in_c_3_data = (io_in_c_input_from_bypass_0 ? io_in_c_bypass_0_3_data : io_in_c_data_3_data); // @[Expression.scala 1420:25]
  assign in_c_3_is_stationary = (io_in_c_input_from_bypass_0 ? io_in_c_bypass_0_3_is_stationary : io_in_c_data_3_is_stationary); // @[Expression.scala 1420:25]
  assign out_r_0_data = pes_0_3_io_out_r_data; // @[SystolicConnect.scala 50:16]
  assign out_r_0_load_store = pes_0_3_io_out_r_load_store; // @[SystolicConnect.scala 50:16]
  assign out_r_0_df_is_ws = pes_0_3_io_out_r_df_is_ws; // @[SystolicConnect.scala 50:16]
  assign out_r_0_stall = pes_0_3_io_out_r_stall; // @[SystolicConnect.scala 50:16]
  assign out_r_1_data = pes_1_3_io_out_r_data; // @[SystolicConnect.scala 50:16]
  assign out_r_1_load_store = pes_1_3_io_out_r_load_store; // @[SystolicConnect.scala 50:16]
  assign out_r_1_df_is_ws = pes_1_3_io_out_r_df_is_ws; // @[SystolicConnect.scala 50:16]
  assign out_r_1_stall = pes_1_3_io_out_r_stall; // @[SystolicConnect.scala 50:16]
  assign out_r_2_data = pes_2_3_io_out_r_data; // @[SystolicConnect.scala 50:16]
  assign out_r_2_load_store = pes_2_3_io_out_r_load_store; // @[SystolicConnect.scala 50:16]
  assign out_r_2_df_is_ws = pes_2_3_io_out_r_df_is_ws; // @[SystolicConnect.scala 50:16]
  assign out_r_2_stall = pes_2_3_io_out_r_stall; // @[SystolicConnect.scala 50:16]
  assign out_r_3_data = pes_3_3_io_out_r_data; // @[SystolicConnect.scala 50:16]
  assign out_r_3_load_store = pes_3_3_io_out_r_load_store; // @[SystolicConnect.scala 50:16]
  assign out_r_3_df_is_ws = pes_3_3_io_out_r_df_is_ws; // @[SystolicConnect.scala 50:16]
  assign out_r_3_stall = pes_3_3_io_out_r_stall; // @[SystolicConnect.scala 50:16]
  assign out_c_0_data = pes_3_0_io_out_c_data; // @[SystolicConnect.scala 56:16]
  assign out_c_0_is_stationary = pes_3_0_io_out_c_is_stationary; // @[SystolicConnect.scala 56:16]
  assign out_c_1_data = pes_3_1_io_out_c_data; // @[SystolicConnect.scala 56:16]
  assign out_c_1_is_stationary = pes_3_1_io_out_c_is_stationary; // @[SystolicConnect.scala 56:16]
  assign out_c_2_data = pes_3_2_io_out_c_data; // @[SystolicConnect.scala 56:16]
  assign out_c_2_is_stationary = pes_3_2_io_out_c_is_stationary; // @[SystolicConnect.scala 56:16]
  assign out_c_3_data = pes_3_3_io_out_c_data; // @[SystolicConnect.scala 56:16]
  assign out_c_3_is_stationary = pes_3_3_io_out_c_is_stationary; // @[SystolicConnect.scala 56:16]
  assign io_out_r_data_0_data = out_r_0_data; // @[ArraySARA.scala 90:17]
  assign io_out_r_data_0_load_store = out_r_0_load_store; // @[ArraySARA.scala 90:17]
  assign io_out_r_data_0_df_is_ws = out_r_0_df_is_ws; // @[ArraySARA.scala 90:17]
  assign io_out_r_data_0_stall = out_r_0_stall; // @[ArraySARA.scala 90:17]
  assign io_out_r_data_1_data = out_r_1_data; // @[ArraySARA.scala 90:17]
  assign io_out_r_data_1_load_store = out_r_1_load_store; // @[ArraySARA.scala 90:17]
  assign io_out_r_data_1_df_is_ws = out_r_1_df_is_ws; // @[ArraySARA.scala 90:17]
  assign io_out_r_data_1_stall = out_r_1_stall; // @[ArraySARA.scala 90:17]
  assign io_out_r_data_2_data = out_r_2_data; // @[ArraySARA.scala 90:17]
  assign io_out_r_data_2_load_store = out_r_2_load_store; // @[ArraySARA.scala 90:17]
  assign io_out_r_data_2_df_is_ws = out_r_2_df_is_ws; // @[ArraySARA.scala 90:17]
  assign io_out_r_data_2_stall = out_r_2_stall; // @[ArraySARA.scala 90:17]
  assign io_out_r_data_3_data = out_r_3_data; // @[ArraySARA.scala 90:17]
  assign io_out_r_data_3_load_store = out_r_3_load_store; // @[ArraySARA.scala 90:17]
  assign io_out_r_data_3_df_is_ws = out_r_3_df_is_ws; // @[ArraySARA.scala 90:17]
  assign io_out_r_data_3_stall = out_r_3_stall; // @[ArraySARA.scala 90:17]
  assign io_out_c_data_0_data = out_c_0_data; // @[ArraySARA.scala 91:17]
  assign io_out_c_data_0_is_stationary = out_c_0_is_stationary; // @[ArraySARA.scala 91:17]
  assign io_out_c_data_1_data = out_c_1_data; // @[ArraySARA.scala 91:17]
  assign io_out_c_data_1_is_stationary = out_c_1_is_stationary; // @[ArraySARA.scala 91:17]
  assign io_out_c_data_2_data = out_c_2_data; // @[ArraySARA.scala 91:17]
  assign io_out_c_data_2_is_stationary = out_c_2_is_stationary; // @[ArraySARA.scala 91:17]
  assign io_out_c_data_3_data = out_c_3_data; // @[ArraySARA.scala 91:17]
  assign io_out_c_data_3_is_stationary = out_c_3_is_stationary; // @[ArraySARA.scala 91:17]
  assign io_out_r_bypass_1_0_data = out_r_regNext_0_data; // @[ArraySARA.scala 92:31]
  assign io_out_r_bypass_1_0_load_store = out_r_regNext_0_load_store; // @[ArraySARA.scala 92:31]
  assign io_out_r_bypass_1_0_df_is_ws = out_r_regNext_0_df_is_ws; // @[ArraySARA.scala 92:31]
  assign io_out_r_bypass_1_0_stall = out_r_regNext_0_stall; // @[ArraySARA.scala 92:31]
  assign io_out_r_bypass_1_1_data = out_r_regNext_1_data; // @[ArraySARA.scala 92:31]
  assign io_out_r_bypass_1_1_load_store = out_r_regNext_1_load_store; // @[ArraySARA.scala 92:31]
  assign io_out_r_bypass_1_1_df_is_ws = out_r_regNext_1_df_is_ws; // @[ArraySARA.scala 92:31]
  assign io_out_r_bypass_1_1_stall = out_r_regNext_1_stall; // @[ArraySARA.scala 92:31]
  assign io_out_r_bypass_1_2_data = out_r_regNext_2_data; // @[ArraySARA.scala 92:31]
  assign io_out_r_bypass_1_2_load_store = out_r_regNext_2_load_store; // @[ArraySARA.scala 92:31]
  assign io_out_r_bypass_1_2_df_is_ws = out_r_regNext_2_df_is_ws; // @[ArraySARA.scala 92:31]
  assign io_out_r_bypass_1_2_stall = out_r_regNext_2_stall; // @[ArraySARA.scala 92:31]
  assign io_out_r_bypass_1_3_data = out_r_regNext_3_data; // @[ArraySARA.scala 92:31]
  assign io_out_r_bypass_1_3_load_store = out_r_regNext_3_load_store; // @[ArraySARA.scala 92:31]
  assign io_out_r_bypass_1_3_df_is_ws = out_r_regNext_3_df_is_ws; // @[ArraySARA.scala 92:31]
  assign io_out_r_bypass_1_3_stall = out_r_regNext_3_stall; // @[ArraySARA.scala 92:31]
  assign io_out_c_bypass_0_0_data = out_c_regNext_0_data; // @[ArraySARA.scala 93:31]
  assign io_out_c_bypass_0_0_is_stationary = out_c_regNext_0_is_stationary; // @[ArraySARA.scala 93:31]
  assign io_out_c_bypass_0_1_data = out_c_regNext_1_data; // @[ArraySARA.scala 93:31]
  assign io_out_c_bypass_0_1_is_stationary = out_c_regNext_1_is_stationary; // @[ArraySARA.scala 93:31]
  assign io_out_c_bypass_0_2_data = out_c_regNext_2_data; // @[ArraySARA.scala 93:31]
  assign io_out_c_bypass_0_2_is_stationary = out_c_regNext_2_is_stationary; // @[ArraySARA.scala 93:31]
  assign io_out_c_bypass_0_3_data = out_c_regNext_3_data; // @[ArraySARA.scala 93:31]
  assign io_out_c_bypass_0_3_is_stationary = out_c_regNext_3_is_stationary; // @[ArraySARA.scala 93:31]
  assign io_out_r_bypass_0_0_data = io_in_r_bypass_regNext_0_0_data; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_0_0_load_store = io_in_r_bypass_regNext_0_0_load_store; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_0_0_df_is_ws = io_in_r_bypass_regNext_0_0_df_is_ws; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_0_0_stall = io_in_r_bypass_regNext_0_0_stall; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_0_1_data = io_in_r_bypass_regNext_0_1_data; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_0_1_load_store = io_in_r_bypass_regNext_0_1_load_store; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_0_1_df_is_ws = io_in_r_bypass_regNext_0_1_df_is_ws; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_0_1_stall = io_in_r_bypass_regNext_0_1_stall; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_0_2_data = io_in_r_bypass_regNext_0_2_data; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_0_2_load_store = io_in_r_bypass_regNext_0_2_load_store; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_0_2_df_is_ws = io_in_r_bypass_regNext_0_2_df_is_ws; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_0_2_stall = io_in_r_bypass_regNext_0_2_stall; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_0_3_data = io_in_r_bypass_regNext_0_3_data; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_0_3_load_store = io_in_r_bypass_regNext_0_3_load_store; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_0_3_df_is_ws = io_in_r_bypass_regNext_0_3_df_is_ws; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_0_3_stall = io_in_r_bypass_regNext_0_3_stall; // @[ArraySARA.scala 97:26]
  assign io_out_c_bypass_1_0_data = io_in_c_bypass_regNext_1_0_data; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_1_0_is_stationary = io_in_c_bypass_regNext_1_0_is_stationary; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_1_1_data = io_in_c_bypass_regNext_1_1_data; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_1_1_is_stationary = io_in_c_bypass_regNext_1_1_is_stationary; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_1_2_data = io_in_c_bypass_regNext_1_2_data; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_1_2_is_stationary = io_in_c_bypass_regNext_1_2_is_stationary; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_1_3_data = io_in_c_bypass_regNext_1_3_data; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_1_3_is_stationary = io_in_c_bypass_regNext_1_3_is_stationary; // @[ArraySARA.scala 101:26]
  assign io_out_r_input_from_bypass_0 = io_in_r_input_from_bypass_regNext_0; // @[ArraySARA.scala 103:30]
  assign io_out_r_input_from_bypass_1 = io_in_r_input_from_bypass_regNext_1; // @[ArraySARA.scala 103:30]
  assign io_out_c_input_from_bypass_0 = io_in_c_input_from_bypass_regNext_0; // @[ArraySARA.scala 104:30]
  assign io_out_c_input_from_bypass_1 = io_in_c_input_from_bypass_regNext_1; // @[ArraySARA.scala 104:30]
  always @(posedge clk) begin
    out_r_regNext_0_data <= out_r_0_data; // @[Reg.scala 39:30]
    out_r_regNext_0_load_store <= out_r_0_load_store; // @[Reg.scala 39:30]
    out_r_regNext_0_df_is_ws <= out_r_0_df_is_ws; // @[Reg.scala 39:30]
    out_r_regNext_0_stall <= out_r_0_stall; // @[Reg.scala 39:30]
    out_r_regNext_1_data <= out_r_1_data; // @[Reg.scala 39:30]
    out_r_regNext_1_load_store <= out_r_1_load_store; // @[Reg.scala 39:30]
    out_r_regNext_1_df_is_ws <= out_r_1_df_is_ws; // @[Reg.scala 39:30]
    out_r_regNext_1_stall <= out_r_1_stall; // @[Reg.scala 39:30]
    out_r_regNext_2_data <= out_r_2_data; // @[Reg.scala 39:30]
    out_r_regNext_2_load_store <= out_r_2_load_store; // @[Reg.scala 39:30]
    out_r_regNext_2_df_is_ws <= out_r_2_df_is_ws; // @[Reg.scala 39:30]
    out_r_regNext_2_stall <= out_r_2_stall; // @[Reg.scala 39:30]
    out_r_regNext_3_data <= out_r_3_data; // @[Reg.scala 39:30]
    out_r_regNext_3_load_store <= out_r_3_load_store; // @[Reg.scala 39:30]
    out_r_regNext_3_df_is_ws <= out_r_3_df_is_ws; // @[Reg.scala 39:30]
    out_r_regNext_3_stall <= out_r_3_stall; // @[Reg.scala 39:30]
    out_c_regNext_0_data <= out_c_0_data; // @[Reg.scala 39:30]
    out_c_regNext_0_is_stationary <= out_c_0_is_stationary; // @[Reg.scala 39:30]
    out_c_regNext_1_data <= out_c_1_data; // @[Reg.scala 39:30]
    out_c_regNext_1_is_stationary <= out_c_1_is_stationary; // @[Reg.scala 39:30]
    out_c_regNext_2_data <= out_c_2_data; // @[Reg.scala 39:30]
    out_c_regNext_2_is_stationary <= out_c_2_is_stationary; // @[Reg.scala 39:30]
    out_c_regNext_3_data <= out_c_3_data; // @[Reg.scala 39:30]
    out_c_regNext_3_is_stationary <= out_c_3_is_stationary; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_0_data <= io_in_r_bypass_0_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_0_load_store <= io_in_r_bypass_0_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_0_df_is_ws <= io_in_r_bypass_0_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_0_stall <= io_in_r_bypass_0_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_1_data <= io_in_r_bypass_0_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_1_load_store <= io_in_r_bypass_0_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_1_df_is_ws <= io_in_r_bypass_0_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_1_stall <= io_in_r_bypass_0_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_2_data <= io_in_r_bypass_0_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_2_load_store <= io_in_r_bypass_0_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_2_df_is_ws <= io_in_r_bypass_0_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_2_stall <= io_in_r_bypass_0_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_3_data <= io_in_r_bypass_0_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_3_load_store <= io_in_r_bypass_0_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_3_df_is_ws <= io_in_r_bypass_0_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_3_stall <= io_in_r_bypass_0_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_0_data <= io_in_r_bypass_1_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_0_load_store <= io_in_r_bypass_1_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_0_df_is_ws <= io_in_r_bypass_1_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_0_stall <= io_in_r_bypass_1_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_1_data <= io_in_r_bypass_1_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_1_load_store <= io_in_r_bypass_1_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_1_df_is_ws <= io_in_r_bypass_1_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_1_stall <= io_in_r_bypass_1_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_2_data <= io_in_r_bypass_1_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_2_load_store <= io_in_r_bypass_1_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_2_df_is_ws <= io_in_r_bypass_1_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_2_stall <= io_in_r_bypass_1_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_3_data <= io_in_r_bypass_1_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_3_load_store <= io_in_r_bypass_1_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_3_df_is_ws <= io_in_r_bypass_1_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_3_stall <= io_in_r_bypass_1_3_stall; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_0_data <= io_in_c_bypass_0_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_0_is_stationary <= io_in_c_bypass_0_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_1_data <= io_in_c_bypass_0_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_1_is_stationary <= io_in_c_bypass_0_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_2_data <= io_in_c_bypass_0_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_2_is_stationary <= io_in_c_bypass_0_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_3_data <= io_in_c_bypass_0_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_3_is_stationary <= io_in_c_bypass_0_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_0_data <= io_in_c_bypass_1_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_0_is_stationary <= io_in_c_bypass_1_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_1_data <= io_in_c_bypass_1_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_1_is_stationary <= io_in_c_bypass_1_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_2_data <= io_in_c_bypass_1_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_2_is_stationary <= io_in_c_bypass_1_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_3_data <= io_in_c_bypass_1_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_3_is_stationary <= io_in_c_bypass_1_3_is_stationary; // @[Reg.scala 39:30]
    io_in_r_input_from_bypass_regNext_0 <= io_in_r_input_from_bypass_0; // @[Reg.scala 39:30]
    io_in_r_input_from_bypass_regNext_1 <= io_in_r_input_from_bypass_1; // @[Reg.scala 39:30]
    io_in_c_input_from_bypass_regNext_0 <= io_in_c_input_from_bypass_0; // @[Reg.scala 39:30]
    io_in_c_input_from_bypass_regNext_1 <= io_in_c_input_from_bypass_1; // @[Reg.scala 39:30]
  end


endmodule

module CellSARA_2 (
  input      [15:0]   io_in_r_data_0_data,
  input               io_in_r_data_0_load_store,
  input               io_in_r_data_0_df_is_ws,
  input               io_in_r_data_0_stall,
  input      [15:0]   io_in_r_data_1_data,
  input               io_in_r_data_1_load_store,
  input               io_in_r_data_1_df_is_ws,
  input               io_in_r_data_1_stall,
  input      [15:0]   io_in_r_data_2_data,
  input               io_in_r_data_2_load_store,
  input               io_in_r_data_2_df_is_ws,
  input               io_in_r_data_2_stall,
  input      [15:0]   io_in_r_data_3_data,
  input               io_in_r_data_3_load_store,
  input               io_in_r_data_3_df_is_ws,
  input               io_in_r_data_3_stall,
  input      [15:0]   io_in_r_bypass_0_0_data,
  input               io_in_r_bypass_0_0_load_store,
  input               io_in_r_bypass_0_0_df_is_ws,
  input               io_in_r_bypass_0_0_stall,
  input      [15:0]   io_in_r_bypass_0_1_data,
  input               io_in_r_bypass_0_1_load_store,
  input               io_in_r_bypass_0_1_df_is_ws,
  input               io_in_r_bypass_0_1_stall,
  input      [15:0]   io_in_r_bypass_0_2_data,
  input               io_in_r_bypass_0_2_load_store,
  input               io_in_r_bypass_0_2_df_is_ws,
  input               io_in_r_bypass_0_2_stall,
  input      [15:0]   io_in_r_bypass_0_3_data,
  input               io_in_r_bypass_0_3_load_store,
  input               io_in_r_bypass_0_3_df_is_ws,
  input               io_in_r_bypass_0_3_stall,
  input      [15:0]   io_in_r_bypass_1_0_data,
  input               io_in_r_bypass_1_0_load_store,
  input               io_in_r_bypass_1_0_df_is_ws,
  input               io_in_r_bypass_1_0_stall,
  input      [15:0]   io_in_r_bypass_1_1_data,
  input               io_in_r_bypass_1_1_load_store,
  input               io_in_r_bypass_1_1_df_is_ws,
  input               io_in_r_bypass_1_1_stall,
  input      [15:0]   io_in_r_bypass_1_2_data,
  input               io_in_r_bypass_1_2_load_store,
  input               io_in_r_bypass_1_2_df_is_ws,
  input               io_in_r_bypass_1_2_stall,
  input      [15:0]   io_in_r_bypass_1_3_data,
  input               io_in_r_bypass_1_3_load_store,
  input               io_in_r_bypass_1_3_df_is_ws,
  input               io_in_r_bypass_1_3_stall,
  input               io_in_r_input_from_bypass_0,
  input               io_in_r_input_from_bypass_1,
  output     [15:0]   io_out_r_data_0_data,
  output              io_out_r_data_0_load_store,
  output              io_out_r_data_0_df_is_ws,
  output              io_out_r_data_0_stall,
  output     [15:0]   io_out_r_data_1_data,
  output              io_out_r_data_1_load_store,
  output              io_out_r_data_1_df_is_ws,
  output              io_out_r_data_1_stall,
  output     [15:0]   io_out_r_data_2_data,
  output              io_out_r_data_2_load_store,
  output              io_out_r_data_2_df_is_ws,
  output              io_out_r_data_2_stall,
  output     [15:0]   io_out_r_data_3_data,
  output              io_out_r_data_3_load_store,
  output              io_out_r_data_3_df_is_ws,
  output              io_out_r_data_3_stall,
  output     [15:0]   io_out_r_bypass_0_0_data,
  output              io_out_r_bypass_0_0_load_store,
  output              io_out_r_bypass_0_0_df_is_ws,
  output              io_out_r_bypass_0_0_stall,
  output     [15:0]   io_out_r_bypass_0_1_data,
  output              io_out_r_bypass_0_1_load_store,
  output              io_out_r_bypass_0_1_df_is_ws,
  output              io_out_r_bypass_0_1_stall,
  output     [15:0]   io_out_r_bypass_0_2_data,
  output              io_out_r_bypass_0_2_load_store,
  output              io_out_r_bypass_0_2_df_is_ws,
  output              io_out_r_bypass_0_2_stall,
  output     [15:0]   io_out_r_bypass_0_3_data,
  output              io_out_r_bypass_0_3_load_store,
  output              io_out_r_bypass_0_3_df_is_ws,
  output              io_out_r_bypass_0_3_stall,
  output     [15:0]   io_out_r_bypass_1_0_data,
  output              io_out_r_bypass_1_0_load_store,
  output              io_out_r_bypass_1_0_df_is_ws,
  output              io_out_r_bypass_1_0_stall,
  output     [15:0]   io_out_r_bypass_1_1_data,
  output              io_out_r_bypass_1_1_load_store,
  output              io_out_r_bypass_1_1_df_is_ws,
  output              io_out_r_bypass_1_1_stall,
  output     [15:0]   io_out_r_bypass_1_2_data,
  output              io_out_r_bypass_1_2_load_store,
  output              io_out_r_bypass_1_2_df_is_ws,
  output              io_out_r_bypass_1_2_stall,
  output     [15:0]   io_out_r_bypass_1_3_data,
  output              io_out_r_bypass_1_3_load_store,
  output              io_out_r_bypass_1_3_df_is_ws,
  output              io_out_r_bypass_1_3_stall,
  output              io_out_r_input_from_bypass_0,
  output              io_out_r_input_from_bypass_1,
  input      [15:0]   io_in_c_data_0_data,
  input               io_in_c_data_0_is_stationary,
  input      [15:0]   io_in_c_data_1_data,
  input               io_in_c_data_1_is_stationary,
  input      [15:0]   io_in_c_data_2_data,
  input               io_in_c_data_2_is_stationary,
  input      [15:0]   io_in_c_data_3_data,
  input               io_in_c_data_3_is_stationary,
  input      [15:0]   io_in_c_bypass_0_0_data,
  input               io_in_c_bypass_0_0_is_stationary,
  input      [15:0]   io_in_c_bypass_0_1_data,
  input               io_in_c_bypass_0_1_is_stationary,
  input      [15:0]   io_in_c_bypass_0_2_data,
  input               io_in_c_bypass_0_2_is_stationary,
  input      [15:0]   io_in_c_bypass_0_3_data,
  input               io_in_c_bypass_0_3_is_stationary,
  input      [15:0]   io_in_c_bypass_1_0_data,
  input               io_in_c_bypass_1_0_is_stationary,
  input      [15:0]   io_in_c_bypass_1_1_data,
  input               io_in_c_bypass_1_1_is_stationary,
  input      [15:0]   io_in_c_bypass_1_2_data,
  input               io_in_c_bypass_1_2_is_stationary,
  input      [15:0]   io_in_c_bypass_1_3_data,
  input               io_in_c_bypass_1_3_is_stationary,
  input               io_in_c_input_from_bypass_0,
  input               io_in_c_input_from_bypass_1,
  output     [15:0]   io_out_c_data_0_data,
  output              io_out_c_data_0_is_stationary,
  output     [15:0]   io_out_c_data_1_data,
  output              io_out_c_data_1_is_stationary,
  output     [15:0]   io_out_c_data_2_data,
  output              io_out_c_data_2_is_stationary,
  output     [15:0]   io_out_c_data_3_data,
  output              io_out_c_data_3_is_stationary,
  output     [15:0]   io_out_c_bypass_0_0_data,
  output              io_out_c_bypass_0_0_is_stationary,
  output     [15:0]   io_out_c_bypass_0_1_data,
  output              io_out_c_bypass_0_1_is_stationary,
  output     [15:0]   io_out_c_bypass_0_2_data,
  output              io_out_c_bypass_0_2_is_stationary,
  output     [15:0]   io_out_c_bypass_0_3_data,
  output              io_out_c_bypass_0_3_is_stationary,
  output     [15:0]   io_out_c_bypass_1_0_data,
  output              io_out_c_bypass_1_0_is_stationary,
  output     [15:0]   io_out_c_bypass_1_1_data,
  output              io_out_c_bypass_1_1_is_stationary,
  output     [15:0]   io_out_c_bypass_1_2_data,
  output              io_out_c_bypass_1_2_is_stationary,
  output     [15:0]   io_out_c_bypass_1_3_data,
  output              io_out_c_bypass_1_3_is_stationary,
  output              io_out_c_input_from_bypass_0,
  output              io_out_c_input_from_bypass_1,
  input               clk,
  input               reset
);

  wire       [15:0]   pes_0_0_io_out_r_data;
  wire                pes_0_0_io_out_r_load_store;
  wire                pes_0_0_io_out_r_df_is_ws;
  wire                pes_0_0_io_out_r_stall;
  wire       [15:0]   pes_0_0_io_out_c_data;
  wire                pes_0_0_io_out_c_is_stationary;
  wire       [15:0]   pes_0_1_io_out_r_data;
  wire                pes_0_1_io_out_r_load_store;
  wire                pes_0_1_io_out_r_df_is_ws;
  wire                pes_0_1_io_out_r_stall;
  wire       [15:0]   pes_0_1_io_out_c_data;
  wire                pes_0_1_io_out_c_is_stationary;
  wire       [15:0]   pes_0_2_io_out_r_data;
  wire                pes_0_2_io_out_r_load_store;
  wire                pes_0_2_io_out_r_df_is_ws;
  wire                pes_0_2_io_out_r_stall;
  wire       [15:0]   pes_0_2_io_out_c_data;
  wire                pes_0_2_io_out_c_is_stationary;
  wire       [15:0]   pes_0_3_io_out_r_data;
  wire                pes_0_3_io_out_r_load_store;
  wire                pes_0_3_io_out_r_df_is_ws;
  wire                pes_0_3_io_out_r_stall;
  wire       [15:0]   pes_0_3_io_out_c_data;
  wire                pes_0_3_io_out_c_is_stationary;
  wire       [15:0]   pes_1_0_io_out_r_data;
  wire                pes_1_0_io_out_r_load_store;
  wire                pes_1_0_io_out_r_df_is_ws;
  wire                pes_1_0_io_out_r_stall;
  wire       [15:0]   pes_1_0_io_out_c_data;
  wire                pes_1_0_io_out_c_is_stationary;
  wire       [15:0]   pes_1_1_io_out_r_data;
  wire                pes_1_1_io_out_r_load_store;
  wire                pes_1_1_io_out_r_df_is_ws;
  wire                pes_1_1_io_out_r_stall;
  wire       [15:0]   pes_1_1_io_out_c_data;
  wire                pes_1_1_io_out_c_is_stationary;
  wire       [15:0]   pes_1_2_io_out_r_data;
  wire                pes_1_2_io_out_r_load_store;
  wire                pes_1_2_io_out_r_df_is_ws;
  wire                pes_1_2_io_out_r_stall;
  wire       [15:0]   pes_1_2_io_out_c_data;
  wire                pes_1_2_io_out_c_is_stationary;
  wire       [15:0]   pes_1_3_io_out_r_data;
  wire                pes_1_3_io_out_r_load_store;
  wire                pes_1_3_io_out_r_df_is_ws;
  wire                pes_1_3_io_out_r_stall;
  wire       [15:0]   pes_1_3_io_out_c_data;
  wire                pes_1_3_io_out_c_is_stationary;
  wire       [15:0]   pes_2_0_io_out_r_data;
  wire                pes_2_0_io_out_r_load_store;
  wire                pes_2_0_io_out_r_df_is_ws;
  wire                pes_2_0_io_out_r_stall;
  wire       [15:0]   pes_2_0_io_out_c_data;
  wire                pes_2_0_io_out_c_is_stationary;
  wire       [15:0]   pes_2_1_io_out_r_data;
  wire                pes_2_1_io_out_r_load_store;
  wire                pes_2_1_io_out_r_df_is_ws;
  wire                pes_2_1_io_out_r_stall;
  wire       [15:0]   pes_2_1_io_out_c_data;
  wire                pes_2_1_io_out_c_is_stationary;
  wire       [15:0]   pes_2_2_io_out_r_data;
  wire                pes_2_2_io_out_r_load_store;
  wire                pes_2_2_io_out_r_df_is_ws;
  wire                pes_2_2_io_out_r_stall;
  wire       [15:0]   pes_2_2_io_out_c_data;
  wire                pes_2_2_io_out_c_is_stationary;
  wire       [15:0]   pes_2_3_io_out_r_data;
  wire                pes_2_3_io_out_r_load_store;
  wire                pes_2_3_io_out_r_df_is_ws;
  wire                pes_2_3_io_out_r_stall;
  wire       [15:0]   pes_2_3_io_out_c_data;
  wire                pes_2_3_io_out_c_is_stationary;
  wire       [15:0]   pes_3_0_io_out_r_data;
  wire                pes_3_0_io_out_r_load_store;
  wire                pes_3_0_io_out_r_df_is_ws;
  wire                pes_3_0_io_out_r_stall;
  wire       [15:0]   pes_3_0_io_out_c_data;
  wire                pes_3_0_io_out_c_is_stationary;
  wire       [15:0]   pes_3_1_io_out_r_data;
  wire                pes_3_1_io_out_r_load_store;
  wire                pes_3_1_io_out_r_df_is_ws;
  wire                pes_3_1_io_out_r_stall;
  wire       [15:0]   pes_3_1_io_out_c_data;
  wire                pes_3_1_io_out_c_is_stationary;
  wire       [15:0]   pes_3_2_io_out_r_data;
  wire                pes_3_2_io_out_r_load_store;
  wire                pes_3_2_io_out_r_df_is_ws;
  wire                pes_3_2_io_out_r_stall;
  wire       [15:0]   pes_3_2_io_out_c_data;
  wire                pes_3_2_io_out_c_is_stationary;
  wire       [15:0]   pes_3_3_io_out_r_data;
  wire                pes_3_3_io_out_r_load_store;
  wire                pes_3_3_io_out_r_df_is_ws;
  wire                pes_3_3_io_out_r_stall;
  wire       [15:0]   pes_3_3_io_out_c_data;
  wire                pes_3_3_io_out_c_is_stationary;
  wire       [15:0]   in_r_0_data;
  wire                in_r_0_load_store;
  wire                in_r_0_df_is_ws;
  wire                in_r_0_stall;
  wire       [15:0]   in_r_1_data;
  wire                in_r_1_load_store;
  wire                in_r_1_df_is_ws;
  wire                in_r_1_stall;
  wire       [15:0]   in_r_2_data;
  wire                in_r_2_load_store;
  wire                in_r_2_df_is_ws;
  wire                in_r_2_stall;
  wire       [15:0]   in_r_3_data;
  wire                in_r_3_load_store;
  wire                in_r_3_df_is_ws;
  wire                in_r_3_stall;
  wire       [15:0]   in_c_0_data;
  wire                in_c_0_is_stationary;
  wire       [15:0]   in_c_1_data;
  wire                in_c_1_is_stationary;
  wire       [15:0]   in_c_2_data;
  wire                in_c_2_is_stationary;
  wire       [15:0]   in_c_3_data;
  wire                in_c_3_is_stationary;
  wire       [15:0]   out_r_0_data;
  wire                out_r_0_load_store;
  wire                out_r_0_df_is_ws;
  wire                out_r_0_stall;
  wire       [15:0]   out_r_1_data;
  wire                out_r_1_load_store;
  wire                out_r_1_df_is_ws;
  wire                out_r_1_stall;
  wire       [15:0]   out_r_2_data;
  wire                out_r_2_load_store;
  wire                out_r_2_df_is_ws;
  wire                out_r_2_stall;
  wire       [15:0]   out_r_3_data;
  wire                out_r_3_load_store;
  wire                out_r_3_df_is_ws;
  wire                out_r_3_stall;
  wire       [15:0]   out_c_0_data;
  wire                out_c_0_is_stationary;
  wire       [15:0]   out_c_1_data;
  wire                out_c_1_is_stationary;
  wire       [15:0]   out_c_2_data;
  wire                out_c_2_is_stationary;
  wire       [15:0]   out_c_3_data;
  wire                out_c_3_is_stationary;
  reg        [15:0]   out_r_regNext_0_data;
  reg                 out_r_regNext_0_load_store;
  reg                 out_r_regNext_0_df_is_ws;
  reg                 out_r_regNext_0_stall;
  reg        [15:0]   out_r_regNext_1_data;
  reg                 out_r_regNext_1_load_store;
  reg                 out_r_regNext_1_df_is_ws;
  reg                 out_r_regNext_1_stall;
  reg        [15:0]   out_r_regNext_2_data;
  reg                 out_r_regNext_2_load_store;
  reg                 out_r_regNext_2_df_is_ws;
  reg                 out_r_regNext_2_stall;
  reg        [15:0]   out_r_regNext_3_data;
  reg                 out_r_regNext_3_load_store;
  reg                 out_r_regNext_3_df_is_ws;
  reg                 out_r_regNext_3_stall;
  reg        [15:0]   out_c_regNext_0_data;
  reg                 out_c_regNext_0_is_stationary;
  reg        [15:0]   out_c_regNext_1_data;
  reg                 out_c_regNext_1_is_stationary;
  reg        [15:0]   out_c_regNext_2_data;
  reg                 out_c_regNext_2_is_stationary;
  reg        [15:0]   out_c_regNext_3_data;
  reg                 out_c_regNext_3_is_stationary;
  reg        [15:0]   io_in_r_bypass_regNext_0_0_data;
  reg                 io_in_r_bypass_regNext_0_0_load_store;
  reg                 io_in_r_bypass_regNext_0_0_df_is_ws;
  reg                 io_in_r_bypass_regNext_0_0_stall;
  reg        [15:0]   io_in_r_bypass_regNext_0_1_data;
  reg                 io_in_r_bypass_regNext_0_1_load_store;
  reg                 io_in_r_bypass_regNext_0_1_df_is_ws;
  reg                 io_in_r_bypass_regNext_0_1_stall;
  reg        [15:0]   io_in_r_bypass_regNext_0_2_data;
  reg                 io_in_r_bypass_regNext_0_2_load_store;
  reg                 io_in_r_bypass_regNext_0_2_df_is_ws;
  reg                 io_in_r_bypass_regNext_0_2_stall;
  reg        [15:0]   io_in_r_bypass_regNext_0_3_data;
  reg                 io_in_r_bypass_regNext_0_3_load_store;
  reg                 io_in_r_bypass_regNext_0_3_df_is_ws;
  reg                 io_in_r_bypass_regNext_0_3_stall;
  reg        [15:0]   io_in_r_bypass_regNext_1_0_data;
  reg                 io_in_r_bypass_regNext_1_0_load_store;
  reg                 io_in_r_bypass_regNext_1_0_df_is_ws;
  reg                 io_in_r_bypass_regNext_1_0_stall;
  reg        [15:0]   io_in_r_bypass_regNext_1_1_data;
  reg                 io_in_r_bypass_regNext_1_1_load_store;
  reg                 io_in_r_bypass_regNext_1_1_df_is_ws;
  reg                 io_in_r_bypass_regNext_1_1_stall;
  reg        [15:0]   io_in_r_bypass_regNext_1_2_data;
  reg                 io_in_r_bypass_regNext_1_2_load_store;
  reg                 io_in_r_bypass_regNext_1_2_df_is_ws;
  reg                 io_in_r_bypass_regNext_1_2_stall;
  reg        [15:0]   io_in_r_bypass_regNext_1_3_data;
  reg                 io_in_r_bypass_regNext_1_3_load_store;
  reg                 io_in_r_bypass_regNext_1_3_df_is_ws;
  reg                 io_in_r_bypass_regNext_1_3_stall;
  reg        [15:0]   io_in_c_bypass_regNext_0_0_data;
  reg                 io_in_c_bypass_regNext_0_0_is_stationary;
  reg        [15:0]   io_in_c_bypass_regNext_0_1_data;
  reg                 io_in_c_bypass_regNext_0_1_is_stationary;
  reg        [15:0]   io_in_c_bypass_regNext_0_2_data;
  reg                 io_in_c_bypass_regNext_0_2_is_stationary;
  reg        [15:0]   io_in_c_bypass_regNext_0_3_data;
  reg                 io_in_c_bypass_regNext_0_3_is_stationary;
  reg        [15:0]   io_in_c_bypass_regNext_1_0_data;
  reg                 io_in_c_bypass_regNext_1_0_is_stationary;
  reg        [15:0]   io_in_c_bypass_regNext_1_1_data;
  reg                 io_in_c_bypass_regNext_1_1_is_stationary;
  reg        [15:0]   io_in_c_bypass_regNext_1_2_data;
  reg                 io_in_c_bypass_regNext_1_2_is_stationary;
  reg        [15:0]   io_in_c_bypass_regNext_1_3_data;
  reg                 io_in_c_bypass_regNext_1_3_is_stationary;
  reg                 io_in_r_input_from_bypass_regNext_0;
  reg                 io_in_r_input_from_bypass_regNext_1;
  reg                 io_in_c_input_from_bypass_regNext_0;
  reg                 io_in_c_input_from_bypass_regNext_1;

  PEWSOS_127 pes_0_0 (
    .io_in_r_data           (in_r_0_data[15:0]             ), //i
    .io_in_r_load_store     (in_r_0_load_store             ), //i
    .io_in_r_df_is_ws       (in_r_0_df_is_ws               ), //i
    .io_in_r_stall          (in_r_0_stall                  ), //i
    .io_out_r_data          (pes_0_0_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pes_0_0_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pes_0_0_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pes_0_0_io_out_r_stall        ), //o
    .io_in_c_data           (in_c_0_data[15:0]             ), //i
    .io_in_c_is_stationary  (in_c_0_is_stationary          ), //i
    .io_out_c_data          (pes_0_0_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pes_0_0_io_out_c_is_stationary), //o
    .clk                    (clk                           ), //i
    .reset                  (reset                         )  //i
  );
  PEWSOS_127 pes_0_1 (
    .io_in_r_data           (pes_0_0_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pes_0_0_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pes_0_0_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pes_0_0_io_out_r_stall        ), //i
    .io_out_r_data          (pes_0_1_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pes_0_1_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pes_0_1_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pes_0_1_io_out_r_stall        ), //o
    .io_in_c_data           (in_c_1_data[15:0]             ), //i
    .io_in_c_is_stationary  (in_c_1_is_stationary          ), //i
    .io_out_c_data          (pes_0_1_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pes_0_1_io_out_c_is_stationary), //o
    .clk                    (clk                           ), //i
    .reset                  (reset                         )  //i
  );
  PEWSOS_127 pes_0_2 (
    .io_in_r_data           (pes_0_1_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pes_0_1_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pes_0_1_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pes_0_1_io_out_r_stall        ), //i
    .io_out_r_data          (pes_0_2_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pes_0_2_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pes_0_2_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pes_0_2_io_out_r_stall        ), //o
    .io_in_c_data           (in_c_2_data[15:0]             ), //i
    .io_in_c_is_stationary  (in_c_2_is_stationary          ), //i
    .io_out_c_data          (pes_0_2_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pes_0_2_io_out_c_is_stationary), //o
    .clk                    (clk                           ), //i
    .reset                  (reset                         )  //i
  );
  PEWSOS_127 pes_0_3 (
    .io_in_r_data           (pes_0_2_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pes_0_2_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pes_0_2_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pes_0_2_io_out_r_stall        ), //i
    .io_out_r_data          (pes_0_3_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pes_0_3_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pes_0_3_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pes_0_3_io_out_r_stall        ), //o
    .io_in_c_data           (in_c_3_data[15:0]             ), //i
    .io_in_c_is_stationary  (in_c_3_is_stationary          ), //i
    .io_out_c_data          (pes_0_3_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pes_0_3_io_out_c_is_stationary), //o
    .clk                    (clk                           ), //i
    .reset                  (reset                         )  //i
  );
  PEWSOS_127 pes_1_0 (
    .io_in_r_data           (in_r_1_data[15:0]             ), //i
    .io_in_r_load_store     (in_r_1_load_store             ), //i
    .io_in_r_df_is_ws       (in_r_1_df_is_ws               ), //i
    .io_in_r_stall          (in_r_1_stall                  ), //i
    .io_out_r_data          (pes_1_0_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pes_1_0_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pes_1_0_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pes_1_0_io_out_r_stall        ), //o
    .io_in_c_data           (pes_0_0_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pes_0_0_io_out_c_is_stationary), //i
    .io_out_c_data          (pes_1_0_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pes_1_0_io_out_c_is_stationary), //o
    .clk                    (clk                           ), //i
    .reset                  (reset                         )  //i
  );
  PEWSOS_127 pes_1_1 (
    .io_in_r_data           (pes_1_0_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pes_1_0_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pes_1_0_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pes_1_0_io_out_r_stall        ), //i
    .io_out_r_data          (pes_1_1_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pes_1_1_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pes_1_1_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pes_1_1_io_out_r_stall        ), //o
    .io_in_c_data           (pes_0_1_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pes_0_1_io_out_c_is_stationary), //i
    .io_out_c_data          (pes_1_1_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pes_1_1_io_out_c_is_stationary), //o
    .clk                    (clk                           ), //i
    .reset                  (reset                         )  //i
  );
  PEWSOS_127 pes_1_2 (
    .io_in_r_data           (pes_1_1_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pes_1_1_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pes_1_1_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pes_1_1_io_out_r_stall        ), //i
    .io_out_r_data          (pes_1_2_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pes_1_2_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pes_1_2_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pes_1_2_io_out_r_stall        ), //o
    .io_in_c_data           (pes_0_2_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pes_0_2_io_out_c_is_stationary), //i
    .io_out_c_data          (pes_1_2_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pes_1_2_io_out_c_is_stationary), //o
    .clk                    (clk                           ), //i
    .reset                  (reset                         )  //i
  );
  PEWSOS_127 pes_1_3 (
    .io_in_r_data           (pes_1_2_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pes_1_2_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pes_1_2_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pes_1_2_io_out_r_stall        ), //i
    .io_out_r_data          (pes_1_3_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pes_1_3_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pes_1_3_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pes_1_3_io_out_r_stall        ), //o
    .io_in_c_data           (pes_0_3_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pes_0_3_io_out_c_is_stationary), //i
    .io_out_c_data          (pes_1_3_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pes_1_3_io_out_c_is_stationary), //o
    .clk                    (clk                           ), //i
    .reset                  (reset                         )  //i
  );
  PEWSOS_127 pes_2_0 (
    .io_in_r_data           (in_r_2_data[15:0]             ), //i
    .io_in_r_load_store     (in_r_2_load_store             ), //i
    .io_in_r_df_is_ws       (in_r_2_df_is_ws               ), //i
    .io_in_r_stall          (in_r_2_stall                  ), //i
    .io_out_r_data          (pes_2_0_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pes_2_0_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pes_2_0_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pes_2_0_io_out_r_stall        ), //o
    .io_in_c_data           (pes_1_0_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pes_1_0_io_out_c_is_stationary), //i
    .io_out_c_data          (pes_2_0_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pes_2_0_io_out_c_is_stationary), //o
    .clk                    (clk                           ), //i
    .reset                  (reset                         )  //i
  );
  PEWSOS_127 pes_2_1 (
    .io_in_r_data           (pes_2_0_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pes_2_0_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pes_2_0_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pes_2_0_io_out_r_stall        ), //i
    .io_out_r_data          (pes_2_1_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pes_2_1_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pes_2_1_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pes_2_1_io_out_r_stall        ), //o
    .io_in_c_data           (pes_1_1_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pes_1_1_io_out_c_is_stationary), //i
    .io_out_c_data          (pes_2_1_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pes_2_1_io_out_c_is_stationary), //o
    .clk                    (clk                           ), //i
    .reset                  (reset                         )  //i
  );
  PEWSOS_127 pes_2_2 (
    .io_in_r_data           (pes_2_1_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pes_2_1_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pes_2_1_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pes_2_1_io_out_r_stall        ), //i
    .io_out_r_data          (pes_2_2_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pes_2_2_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pes_2_2_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pes_2_2_io_out_r_stall        ), //o
    .io_in_c_data           (pes_1_2_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pes_1_2_io_out_c_is_stationary), //i
    .io_out_c_data          (pes_2_2_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pes_2_2_io_out_c_is_stationary), //o
    .clk                    (clk                           ), //i
    .reset                  (reset                         )  //i
  );
  PEWSOS_127 pes_2_3 (
    .io_in_r_data           (pes_2_2_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pes_2_2_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pes_2_2_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pes_2_2_io_out_r_stall        ), //i
    .io_out_r_data          (pes_2_3_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pes_2_3_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pes_2_3_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pes_2_3_io_out_r_stall        ), //o
    .io_in_c_data           (pes_1_3_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pes_1_3_io_out_c_is_stationary), //i
    .io_out_c_data          (pes_2_3_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pes_2_3_io_out_c_is_stationary), //o
    .clk                    (clk                           ), //i
    .reset                  (reset                         )  //i
  );
  PEWSOS_127 pes_3_0 (
    .io_in_r_data           (in_r_3_data[15:0]             ), //i
    .io_in_r_load_store     (in_r_3_load_store             ), //i
    .io_in_r_df_is_ws       (in_r_3_df_is_ws               ), //i
    .io_in_r_stall          (in_r_3_stall                  ), //i
    .io_out_r_data          (pes_3_0_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pes_3_0_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pes_3_0_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pes_3_0_io_out_r_stall        ), //o
    .io_in_c_data           (pes_2_0_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pes_2_0_io_out_c_is_stationary), //i
    .io_out_c_data          (pes_3_0_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pes_3_0_io_out_c_is_stationary), //o
    .clk                    (clk                           ), //i
    .reset                  (reset                         )  //i
  );
  PEWSOS_127 pes_3_1 (
    .io_in_r_data           (pes_3_0_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pes_3_0_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pes_3_0_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pes_3_0_io_out_r_stall        ), //i
    .io_out_r_data          (pes_3_1_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pes_3_1_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pes_3_1_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pes_3_1_io_out_r_stall        ), //o
    .io_in_c_data           (pes_2_1_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pes_2_1_io_out_c_is_stationary), //i
    .io_out_c_data          (pes_3_1_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pes_3_1_io_out_c_is_stationary), //o
    .clk                    (clk                           ), //i
    .reset                  (reset                         )  //i
  );
  PEWSOS_127 pes_3_2 (
    .io_in_r_data           (pes_3_1_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pes_3_1_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pes_3_1_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pes_3_1_io_out_r_stall        ), //i
    .io_out_r_data          (pes_3_2_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pes_3_2_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pes_3_2_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pes_3_2_io_out_r_stall        ), //o
    .io_in_c_data           (pes_2_2_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pes_2_2_io_out_c_is_stationary), //i
    .io_out_c_data          (pes_3_2_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pes_3_2_io_out_c_is_stationary), //o
    .clk                    (clk                           ), //i
    .reset                  (reset                         )  //i
  );
  PEWSOS_127 pes_3_3 (
    .io_in_r_data           (pes_3_2_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pes_3_2_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pes_3_2_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pes_3_2_io_out_r_stall        ), //i
    .io_out_r_data          (pes_3_3_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pes_3_3_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pes_3_3_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pes_3_3_io_out_r_stall        ), //o
    .io_in_c_data           (pes_2_3_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pes_2_3_io_out_c_is_stationary), //i
    .io_out_c_data          (pes_3_3_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pes_3_3_io_out_c_is_stationary), //o
    .clk                    (clk                           ), //i
    .reset                  (reset                         )  //i
  );
  assign in_r_0_data = (io_in_r_input_from_bypass_0 ? io_in_r_bypass_0_0_data : io_in_r_data_0_data); // @[Expression.scala 1420:25]
  assign in_r_0_load_store = (io_in_r_input_from_bypass_0 ? io_in_r_bypass_0_0_load_store : io_in_r_data_0_load_store); // @[Expression.scala 1420:25]
  assign in_r_0_df_is_ws = (io_in_r_input_from_bypass_0 ? io_in_r_bypass_0_0_df_is_ws : io_in_r_data_0_df_is_ws); // @[Expression.scala 1420:25]
  assign in_r_0_stall = (io_in_r_input_from_bypass_0 ? io_in_r_bypass_0_0_stall : io_in_r_data_0_stall); // @[Expression.scala 1420:25]
  assign in_r_1_data = (io_in_r_input_from_bypass_0 ? io_in_r_bypass_0_1_data : io_in_r_data_1_data); // @[Expression.scala 1420:25]
  assign in_r_1_load_store = (io_in_r_input_from_bypass_0 ? io_in_r_bypass_0_1_load_store : io_in_r_data_1_load_store); // @[Expression.scala 1420:25]
  assign in_r_1_df_is_ws = (io_in_r_input_from_bypass_0 ? io_in_r_bypass_0_1_df_is_ws : io_in_r_data_1_df_is_ws); // @[Expression.scala 1420:25]
  assign in_r_1_stall = (io_in_r_input_from_bypass_0 ? io_in_r_bypass_0_1_stall : io_in_r_data_1_stall); // @[Expression.scala 1420:25]
  assign in_r_2_data = (io_in_r_input_from_bypass_0 ? io_in_r_bypass_0_2_data : io_in_r_data_2_data); // @[Expression.scala 1420:25]
  assign in_r_2_load_store = (io_in_r_input_from_bypass_0 ? io_in_r_bypass_0_2_load_store : io_in_r_data_2_load_store); // @[Expression.scala 1420:25]
  assign in_r_2_df_is_ws = (io_in_r_input_from_bypass_0 ? io_in_r_bypass_0_2_df_is_ws : io_in_r_data_2_df_is_ws); // @[Expression.scala 1420:25]
  assign in_r_2_stall = (io_in_r_input_from_bypass_0 ? io_in_r_bypass_0_2_stall : io_in_r_data_2_stall); // @[Expression.scala 1420:25]
  assign in_r_3_data = (io_in_r_input_from_bypass_0 ? io_in_r_bypass_0_3_data : io_in_r_data_3_data); // @[Expression.scala 1420:25]
  assign in_r_3_load_store = (io_in_r_input_from_bypass_0 ? io_in_r_bypass_0_3_load_store : io_in_r_data_3_load_store); // @[Expression.scala 1420:25]
  assign in_r_3_df_is_ws = (io_in_r_input_from_bypass_0 ? io_in_r_bypass_0_3_df_is_ws : io_in_r_data_3_df_is_ws); // @[Expression.scala 1420:25]
  assign in_r_3_stall = (io_in_r_input_from_bypass_0 ? io_in_r_bypass_0_3_stall : io_in_r_data_3_stall); // @[Expression.scala 1420:25]
  assign in_c_0_data = (io_in_c_input_from_bypass_1 ? io_in_c_bypass_1_0_data : io_in_c_data_0_data); // @[Expression.scala 1420:25]
  assign in_c_0_is_stationary = (io_in_c_input_from_bypass_1 ? io_in_c_bypass_1_0_is_stationary : io_in_c_data_0_is_stationary); // @[Expression.scala 1420:25]
  assign in_c_1_data = (io_in_c_input_from_bypass_1 ? io_in_c_bypass_1_1_data : io_in_c_data_1_data); // @[Expression.scala 1420:25]
  assign in_c_1_is_stationary = (io_in_c_input_from_bypass_1 ? io_in_c_bypass_1_1_is_stationary : io_in_c_data_1_is_stationary); // @[Expression.scala 1420:25]
  assign in_c_2_data = (io_in_c_input_from_bypass_1 ? io_in_c_bypass_1_2_data : io_in_c_data_2_data); // @[Expression.scala 1420:25]
  assign in_c_2_is_stationary = (io_in_c_input_from_bypass_1 ? io_in_c_bypass_1_2_is_stationary : io_in_c_data_2_is_stationary); // @[Expression.scala 1420:25]
  assign in_c_3_data = (io_in_c_input_from_bypass_1 ? io_in_c_bypass_1_3_data : io_in_c_data_3_data); // @[Expression.scala 1420:25]
  assign in_c_3_is_stationary = (io_in_c_input_from_bypass_1 ? io_in_c_bypass_1_3_is_stationary : io_in_c_data_3_is_stationary); // @[Expression.scala 1420:25]
  assign out_r_0_data = pes_0_3_io_out_r_data; // @[SystolicConnect.scala 50:16]
  assign out_r_0_load_store = pes_0_3_io_out_r_load_store; // @[SystolicConnect.scala 50:16]
  assign out_r_0_df_is_ws = pes_0_3_io_out_r_df_is_ws; // @[SystolicConnect.scala 50:16]
  assign out_r_0_stall = pes_0_3_io_out_r_stall; // @[SystolicConnect.scala 50:16]
  assign out_r_1_data = pes_1_3_io_out_r_data; // @[SystolicConnect.scala 50:16]
  assign out_r_1_load_store = pes_1_3_io_out_r_load_store; // @[SystolicConnect.scala 50:16]
  assign out_r_1_df_is_ws = pes_1_3_io_out_r_df_is_ws; // @[SystolicConnect.scala 50:16]
  assign out_r_1_stall = pes_1_3_io_out_r_stall; // @[SystolicConnect.scala 50:16]
  assign out_r_2_data = pes_2_3_io_out_r_data; // @[SystolicConnect.scala 50:16]
  assign out_r_2_load_store = pes_2_3_io_out_r_load_store; // @[SystolicConnect.scala 50:16]
  assign out_r_2_df_is_ws = pes_2_3_io_out_r_df_is_ws; // @[SystolicConnect.scala 50:16]
  assign out_r_2_stall = pes_2_3_io_out_r_stall; // @[SystolicConnect.scala 50:16]
  assign out_r_3_data = pes_3_3_io_out_r_data; // @[SystolicConnect.scala 50:16]
  assign out_r_3_load_store = pes_3_3_io_out_r_load_store; // @[SystolicConnect.scala 50:16]
  assign out_r_3_df_is_ws = pes_3_3_io_out_r_df_is_ws; // @[SystolicConnect.scala 50:16]
  assign out_r_3_stall = pes_3_3_io_out_r_stall; // @[SystolicConnect.scala 50:16]
  assign out_c_0_data = pes_3_0_io_out_c_data; // @[SystolicConnect.scala 56:16]
  assign out_c_0_is_stationary = pes_3_0_io_out_c_is_stationary; // @[SystolicConnect.scala 56:16]
  assign out_c_1_data = pes_3_1_io_out_c_data; // @[SystolicConnect.scala 56:16]
  assign out_c_1_is_stationary = pes_3_1_io_out_c_is_stationary; // @[SystolicConnect.scala 56:16]
  assign out_c_2_data = pes_3_2_io_out_c_data; // @[SystolicConnect.scala 56:16]
  assign out_c_2_is_stationary = pes_3_2_io_out_c_is_stationary; // @[SystolicConnect.scala 56:16]
  assign out_c_3_data = pes_3_3_io_out_c_data; // @[SystolicConnect.scala 56:16]
  assign out_c_3_is_stationary = pes_3_3_io_out_c_is_stationary; // @[SystolicConnect.scala 56:16]
  assign io_out_r_data_0_data = out_r_0_data; // @[ArraySARA.scala 90:17]
  assign io_out_r_data_0_load_store = out_r_0_load_store; // @[ArraySARA.scala 90:17]
  assign io_out_r_data_0_df_is_ws = out_r_0_df_is_ws; // @[ArraySARA.scala 90:17]
  assign io_out_r_data_0_stall = out_r_0_stall; // @[ArraySARA.scala 90:17]
  assign io_out_r_data_1_data = out_r_1_data; // @[ArraySARA.scala 90:17]
  assign io_out_r_data_1_load_store = out_r_1_load_store; // @[ArraySARA.scala 90:17]
  assign io_out_r_data_1_df_is_ws = out_r_1_df_is_ws; // @[ArraySARA.scala 90:17]
  assign io_out_r_data_1_stall = out_r_1_stall; // @[ArraySARA.scala 90:17]
  assign io_out_r_data_2_data = out_r_2_data; // @[ArraySARA.scala 90:17]
  assign io_out_r_data_2_load_store = out_r_2_load_store; // @[ArraySARA.scala 90:17]
  assign io_out_r_data_2_df_is_ws = out_r_2_df_is_ws; // @[ArraySARA.scala 90:17]
  assign io_out_r_data_2_stall = out_r_2_stall; // @[ArraySARA.scala 90:17]
  assign io_out_r_data_3_data = out_r_3_data; // @[ArraySARA.scala 90:17]
  assign io_out_r_data_3_load_store = out_r_3_load_store; // @[ArraySARA.scala 90:17]
  assign io_out_r_data_3_df_is_ws = out_r_3_df_is_ws; // @[ArraySARA.scala 90:17]
  assign io_out_r_data_3_stall = out_r_3_stall; // @[ArraySARA.scala 90:17]
  assign io_out_c_data_0_data = out_c_0_data; // @[ArraySARA.scala 91:17]
  assign io_out_c_data_0_is_stationary = out_c_0_is_stationary; // @[ArraySARA.scala 91:17]
  assign io_out_c_data_1_data = out_c_1_data; // @[ArraySARA.scala 91:17]
  assign io_out_c_data_1_is_stationary = out_c_1_is_stationary; // @[ArraySARA.scala 91:17]
  assign io_out_c_data_2_data = out_c_2_data; // @[ArraySARA.scala 91:17]
  assign io_out_c_data_2_is_stationary = out_c_2_is_stationary; // @[ArraySARA.scala 91:17]
  assign io_out_c_data_3_data = out_c_3_data; // @[ArraySARA.scala 91:17]
  assign io_out_c_data_3_is_stationary = out_c_3_is_stationary; // @[ArraySARA.scala 91:17]
  assign io_out_r_bypass_0_0_data = out_r_regNext_0_data; // @[ArraySARA.scala 92:31]
  assign io_out_r_bypass_0_0_load_store = out_r_regNext_0_load_store; // @[ArraySARA.scala 92:31]
  assign io_out_r_bypass_0_0_df_is_ws = out_r_regNext_0_df_is_ws; // @[ArraySARA.scala 92:31]
  assign io_out_r_bypass_0_0_stall = out_r_regNext_0_stall; // @[ArraySARA.scala 92:31]
  assign io_out_r_bypass_0_1_data = out_r_regNext_1_data; // @[ArraySARA.scala 92:31]
  assign io_out_r_bypass_0_1_load_store = out_r_regNext_1_load_store; // @[ArraySARA.scala 92:31]
  assign io_out_r_bypass_0_1_df_is_ws = out_r_regNext_1_df_is_ws; // @[ArraySARA.scala 92:31]
  assign io_out_r_bypass_0_1_stall = out_r_regNext_1_stall; // @[ArraySARA.scala 92:31]
  assign io_out_r_bypass_0_2_data = out_r_regNext_2_data; // @[ArraySARA.scala 92:31]
  assign io_out_r_bypass_0_2_load_store = out_r_regNext_2_load_store; // @[ArraySARA.scala 92:31]
  assign io_out_r_bypass_0_2_df_is_ws = out_r_regNext_2_df_is_ws; // @[ArraySARA.scala 92:31]
  assign io_out_r_bypass_0_2_stall = out_r_regNext_2_stall; // @[ArraySARA.scala 92:31]
  assign io_out_r_bypass_0_3_data = out_r_regNext_3_data; // @[ArraySARA.scala 92:31]
  assign io_out_r_bypass_0_3_load_store = out_r_regNext_3_load_store; // @[ArraySARA.scala 92:31]
  assign io_out_r_bypass_0_3_df_is_ws = out_r_regNext_3_df_is_ws; // @[ArraySARA.scala 92:31]
  assign io_out_r_bypass_0_3_stall = out_r_regNext_3_stall; // @[ArraySARA.scala 92:31]
  assign io_out_c_bypass_1_0_data = out_c_regNext_0_data; // @[ArraySARA.scala 93:31]
  assign io_out_c_bypass_1_0_is_stationary = out_c_regNext_0_is_stationary; // @[ArraySARA.scala 93:31]
  assign io_out_c_bypass_1_1_data = out_c_regNext_1_data; // @[ArraySARA.scala 93:31]
  assign io_out_c_bypass_1_1_is_stationary = out_c_regNext_1_is_stationary; // @[ArraySARA.scala 93:31]
  assign io_out_c_bypass_1_2_data = out_c_regNext_2_data; // @[ArraySARA.scala 93:31]
  assign io_out_c_bypass_1_2_is_stationary = out_c_regNext_2_is_stationary; // @[ArraySARA.scala 93:31]
  assign io_out_c_bypass_1_3_data = out_c_regNext_3_data; // @[ArraySARA.scala 93:31]
  assign io_out_c_bypass_1_3_is_stationary = out_c_regNext_3_is_stationary; // @[ArraySARA.scala 93:31]
  assign io_out_r_bypass_1_0_data = io_in_r_bypass_regNext_1_0_data; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_1_0_load_store = io_in_r_bypass_regNext_1_0_load_store; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_1_0_df_is_ws = io_in_r_bypass_regNext_1_0_df_is_ws; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_1_0_stall = io_in_r_bypass_regNext_1_0_stall; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_1_1_data = io_in_r_bypass_regNext_1_1_data; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_1_1_load_store = io_in_r_bypass_regNext_1_1_load_store; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_1_1_df_is_ws = io_in_r_bypass_regNext_1_1_df_is_ws; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_1_1_stall = io_in_r_bypass_regNext_1_1_stall; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_1_2_data = io_in_r_bypass_regNext_1_2_data; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_1_2_load_store = io_in_r_bypass_regNext_1_2_load_store; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_1_2_df_is_ws = io_in_r_bypass_regNext_1_2_df_is_ws; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_1_2_stall = io_in_r_bypass_regNext_1_2_stall; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_1_3_data = io_in_r_bypass_regNext_1_3_data; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_1_3_load_store = io_in_r_bypass_regNext_1_3_load_store; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_1_3_df_is_ws = io_in_r_bypass_regNext_1_3_df_is_ws; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_1_3_stall = io_in_r_bypass_regNext_1_3_stall; // @[ArraySARA.scala 97:26]
  assign io_out_c_bypass_0_0_data = io_in_c_bypass_regNext_0_0_data; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_0_0_is_stationary = io_in_c_bypass_regNext_0_0_is_stationary; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_0_1_data = io_in_c_bypass_regNext_0_1_data; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_0_1_is_stationary = io_in_c_bypass_regNext_0_1_is_stationary; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_0_2_data = io_in_c_bypass_regNext_0_2_data; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_0_2_is_stationary = io_in_c_bypass_regNext_0_2_is_stationary; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_0_3_data = io_in_c_bypass_regNext_0_3_data; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_0_3_is_stationary = io_in_c_bypass_regNext_0_3_is_stationary; // @[ArraySARA.scala 101:26]
  assign io_out_r_input_from_bypass_0 = io_in_r_input_from_bypass_regNext_0; // @[ArraySARA.scala 103:30]
  assign io_out_r_input_from_bypass_1 = io_in_r_input_from_bypass_regNext_1; // @[ArraySARA.scala 103:30]
  assign io_out_c_input_from_bypass_0 = io_in_c_input_from_bypass_regNext_0; // @[ArraySARA.scala 104:30]
  assign io_out_c_input_from_bypass_1 = io_in_c_input_from_bypass_regNext_1; // @[ArraySARA.scala 104:30]
  always @(posedge clk) begin
    out_r_regNext_0_data <= out_r_0_data; // @[Reg.scala 39:30]
    out_r_regNext_0_load_store <= out_r_0_load_store; // @[Reg.scala 39:30]
    out_r_regNext_0_df_is_ws <= out_r_0_df_is_ws; // @[Reg.scala 39:30]
    out_r_regNext_0_stall <= out_r_0_stall; // @[Reg.scala 39:30]
    out_r_regNext_1_data <= out_r_1_data; // @[Reg.scala 39:30]
    out_r_regNext_1_load_store <= out_r_1_load_store; // @[Reg.scala 39:30]
    out_r_regNext_1_df_is_ws <= out_r_1_df_is_ws; // @[Reg.scala 39:30]
    out_r_regNext_1_stall <= out_r_1_stall; // @[Reg.scala 39:30]
    out_r_regNext_2_data <= out_r_2_data; // @[Reg.scala 39:30]
    out_r_regNext_2_load_store <= out_r_2_load_store; // @[Reg.scala 39:30]
    out_r_regNext_2_df_is_ws <= out_r_2_df_is_ws; // @[Reg.scala 39:30]
    out_r_regNext_2_stall <= out_r_2_stall; // @[Reg.scala 39:30]
    out_r_regNext_3_data <= out_r_3_data; // @[Reg.scala 39:30]
    out_r_regNext_3_load_store <= out_r_3_load_store; // @[Reg.scala 39:30]
    out_r_regNext_3_df_is_ws <= out_r_3_df_is_ws; // @[Reg.scala 39:30]
    out_r_regNext_3_stall <= out_r_3_stall; // @[Reg.scala 39:30]
    out_c_regNext_0_data <= out_c_0_data; // @[Reg.scala 39:30]
    out_c_regNext_0_is_stationary <= out_c_0_is_stationary; // @[Reg.scala 39:30]
    out_c_regNext_1_data <= out_c_1_data; // @[Reg.scala 39:30]
    out_c_regNext_1_is_stationary <= out_c_1_is_stationary; // @[Reg.scala 39:30]
    out_c_regNext_2_data <= out_c_2_data; // @[Reg.scala 39:30]
    out_c_regNext_2_is_stationary <= out_c_2_is_stationary; // @[Reg.scala 39:30]
    out_c_regNext_3_data <= out_c_3_data; // @[Reg.scala 39:30]
    out_c_regNext_3_is_stationary <= out_c_3_is_stationary; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_0_data <= io_in_r_bypass_0_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_0_load_store <= io_in_r_bypass_0_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_0_df_is_ws <= io_in_r_bypass_0_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_0_stall <= io_in_r_bypass_0_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_1_data <= io_in_r_bypass_0_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_1_load_store <= io_in_r_bypass_0_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_1_df_is_ws <= io_in_r_bypass_0_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_1_stall <= io_in_r_bypass_0_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_2_data <= io_in_r_bypass_0_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_2_load_store <= io_in_r_bypass_0_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_2_df_is_ws <= io_in_r_bypass_0_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_2_stall <= io_in_r_bypass_0_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_3_data <= io_in_r_bypass_0_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_3_load_store <= io_in_r_bypass_0_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_3_df_is_ws <= io_in_r_bypass_0_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_3_stall <= io_in_r_bypass_0_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_0_data <= io_in_r_bypass_1_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_0_load_store <= io_in_r_bypass_1_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_0_df_is_ws <= io_in_r_bypass_1_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_0_stall <= io_in_r_bypass_1_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_1_data <= io_in_r_bypass_1_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_1_load_store <= io_in_r_bypass_1_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_1_df_is_ws <= io_in_r_bypass_1_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_1_stall <= io_in_r_bypass_1_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_2_data <= io_in_r_bypass_1_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_2_load_store <= io_in_r_bypass_1_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_2_df_is_ws <= io_in_r_bypass_1_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_2_stall <= io_in_r_bypass_1_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_3_data <= io_in_r_bypass_1_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_3_load_store <= io_in_r_bypass_1_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_3_df_is_ws <= io_in_r_bypass_1_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_3_stall <= io_in_r_bypass_1_3_stall; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_0_data <= io_in_c_bypass_0_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_0_is_stationary <= io_in_c_bypass_0_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_1_data <= io_in_c_bypass_0_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_1_is_stationary <= io_in_c_bypass_0_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_2_data <= io_in_c_bypass_0_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_2_is_stationary <= io_in_c_bypass_0_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_3_data <= io_in_c_bypass_0_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_3_is_stationary <= io_in_c_bypass_0_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_0_data <= io_in_c_bypass_1_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_0_is_stationary <= io_in_c_bypass_1_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_1_data <= io_in_c_bypass_1_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_1_is_stationary <= io_in_c_bypass_1_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_2_data <= io_in_c_bypass_1_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_2_is_stationary <= io_in_c_bypass_1_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_3_data <= io_in_c_bypass_1_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_3_is_stationary <= io_in_c_bypass_1_3_is_stationary; // @[Reg.scala 39:30]
    io_in_r_input_from_bypass_regNext_0 <= io_in_r_input_from_bypass_0; // @[Reg.scala 39:30]
    io_in_r_input_from_bypass_regNext_1 <= io_in_r_input_from_bypass_1; // @[Reg.scala 39:30]
    io_in_c_input_from_bypass_regNext_0 <= io_in_c_input_from_bypass_0; // @[Reg.scala 39:30]
    io_in_c_input_from_bypass_regNext_1 <= io_in_c_input_from_bypass_1; // @[Reg.scala 39:30]
  end


endmodule

//CellSARA_7 replaced by CellSARA_7

//CellSARA_7 replaced by CellSARA_7

//CellSARA_7 replaced by CellSARA_7

//CellSARA_7 replaced by CellSARA_7

module CellSARA_7 (
  input      [15:0]   io_in_r_data_0_data,
  input               io_in_r_data_0_load_store,
  input               io_in_r_data_0_df_is_ws,
  input               io_in_r_data_0_stall,
  input      [15:0]   io_in_r_data_1_data,
  input               io_in_r_data_1_load_store,
  input               io_in_r_data_1_df_is_ws,
  input               io_in_r_data_1_stall,
  input      [15:0]   io_in_r_data_2_data,
  input               io_in_r_data_2_load_store,
  input               io_in_r_data_2_df_is_ws,
  input               io_in_r_data_2_stall,
  input      [15:0]   io_in_r_data_3_data,
  input               io_in_r_data_3_load_store,
  input               io_in_r_data_3_df_is_ws,
  input               io_in_r_data_3_stall,
  input      [15:0]   io_in_r_bypass_0_0_data,
  input               io_in_r_bypass_0_0_load_store,
  input               io_in_r_bypass_0_0_df_is_ws,
  input               io_in_r_bypass_0_0_stall,
  input      [15:0]   io_in_r_bypass_0_1_data,
  input               io_in_r_bypass_0_1_load_store,
  input               io_in_r_bypass_0_1_df_is_ws,
  input               io_in_r_bypass_0_1_stall,
  input      [15:0]   io_in_r_bypass_0_2_data,
  input               io_in_r_bypass_0_2_load_store,
  input               io_in_r_bypass_0_2_df_is_ws,
  input               io_in_r_bypass_0_2_stall,
  input      [15:0]   io_in_r_bypass_0_3_data,
  input               io_in_r_bypass_0_3_load_store,
  input               io_in_r_bypass_0_3_df_is_ws,
  input               io_in_r_bypass_0_3_stall,
  input      [15:0]   io_in_r_bypass_1_0_data,
  input               io_in_r_bypass_1_0_load_store,
  input               io_in_r_bypass_1_0_df_is_ws,
  input               io_in_r_bypass_1_0_stall,
  input      [15:0]   io_in_r_bypass_1_1_data,
  input               io_in_r_bypass_1_1_load_store,
  input               io_in_r_bypass_1_1_df_is_ws,
  input               io_in_r_bypass_1_1_stall,
  input      [15:0]   io_in_r_bypass_1_2_data,
  input               io_in_r_bypass_1_2_load_store,
  input               io_in_r_bypass_1_2_df_is_ws,
  input               io_in_r_bypass_1_2_stall,
  input      [15:0]   io_in_r_bypass_1_3_data,
  input               io_in_r_bypass_1_3_load_store,
  input               io_in_r_bypass_1_3_df_is_ws,
  input               io_in_r_bypass_1_3_stall,
  input               io_in_r_input_from_bypass_0,
  input               io_in_r_input_from_bypass_1,
  output     [15:0]   io_out_r_data_0_data,
  output              io_out_r_data_0_load_store,
  output              io_out_r_data_0_df_is_ws,
  output              io_out_r_data_0_stall,
  output     [15:0]   io_out_r_data_1_data,
  output              io_out_r_data_1_load_store,
  output              io_out_r_data_1_df_is_ws,
  output              io_out_r_data_1_stall,
  output     [15:0]   io_out_r_data_2_data,
  output              io_out_r_data_2_load_store,
  output              io_out_r_data_2_df_is_ws,
  output              io_out_r_data_2_stall,
  output     [15:0]   io_out_r_data_3_data,
  output              io_out_r_data_3_load_store,
  output              io_out_r_data_3_df_is_ws,
  output              io_out_r_data_3_stall,
  output     [15:0]   io_out_r_bypass_0_0_data,
  output              io_out_r_bypass_0_0_load_store,
  output              io_out_r_bypass_0_0_df_is_ws,
  output              io_out_r_bypass_0_0_stall,
  output     [15:0]   io_out_r_bypass_0_1_data,
  output              io_out_r_bypass_0_1_load_store,
  output              io_out_r_bypass_0_1_df_is_ws,
  output              io_out_r_bypass_0_1_stall,
  output     [15:0]   io_out_r_bypass_0_2_data,
  output              io_out_r_bypass_0_2_load_store,
  output              io_out_r_bypass_0_2_df_is_ws,
  output              io_out_r_bypass_0_2_stall,
  output     [15:0]   io_out_r_bypass_0_3_data,
  output              io_out_r_bypass_0_3_load_store,
  output              io_out_r_bypass_0_3_df_is_ws,
  output              io_out_r_bypass_0_3_stall,
  output     [15:0]   io_out_r_bypass_1_0_data,
  output              io_out_r_bypass_1_0_load_store,
  output              io_out_r_bypass_1_0_df_is_ws,
  output              io_out_r_bypass_1_0_stall,
  output     [15:0]   io_out_r_bypass_1_1_data,
  output              io_out_r_bypass_1_1_load_store,
  output              io_out_r_bypass_1_1_df_is_ws,
  output              io_out_r_bypass_1_1_stall,
  output     [15:0]   io_out_r_bypass_1_2_data,
  output              io_out_r_bypass_1_2_load_store,
  output              io_out_r_bypass_1_2_df_is_ws,
  output              io_out_r_bypass_1_2_stall,
  output     [15:0]   io_out_r_bypass_1_3_data,
  output              io_out_r_bypass_1_3_load_store,
  output              io_out_r_bypass_1_3_df_is_ws,
  output              io_out_r_bypass_1_3_stall,
  output              io_out_r_input_from_bypass_0,
  output              io_out_r_input_from_bypass_1,
  input      [15:0]   io_in_c_data_0_data,
  input               io_in_c_data_0_is_stationary,
  input      [15:0]   io_in_c_data_1_data,
  input               io_in_c_data_1_is_stationary,
  input      [15:0]   io_in_c_data_2_data,
  input               io_in_c_data_2_is_stationary,
  input      [15:0]   io_in_c_data_3_data,
  input               io_in_c_data_3_is_stationary,
  input      [15:0]   io_in_c_bypass_0_0_data,
  input               io_in_c_bypass_0_0_is_stationary,
  input      [15:0]   io_in_c_bypass_0_1_data,
  input               io_in_c_bypass_0_1_is_stationary,
  input      [15:0]   io_in_c_bypass_0_2_data,
  input               io_in_c_bypass_0_2_is_stationary,
  input      [15:0]   io_in_c_bypass_0_3_data,
  input               io_in_c_bypass_0_3_is_stationary,
  input      [15:0]   io_in_c_bypass_1_0_data,
  input               io_in_c_bypass_1_0_is_stationary,
  input      [15:0]   io_in_c_bypass_1_1_data,
  input               io_in_c_bypass_1_1_is_stationary,
  input      [15:0]   io_in_c_bypass_1_2_data,
  input               io_in_c_bypass_1_2_is_stationary,
  input      [15:0]   io_in_c_bypass_1_3_data,
  input               io_in_c_bypass_1_3_is_stationary,
  input               io_in_c_input_from_bypass_0,
  input               io_in_c_input_from_bypass_1,
  output     [15:0]   io_out_c_data_0_data,
  output              io_out_c_data_0_is_stationary,
  output     [15:0]   io_out_c_data_1_data,
  output              io_out_c_data_1_is_stationary,
  output     [15:0]   io_out_c_data_2_data,
  output              io_out_c_data_2_is_stationary,
  output     [15:0]   io_out_c_data_3_data,
  output              io_out_c_data_3_is_stationary,
  output     [15:0]   io_out_c_bypass_0_0_data,
  output              io_out_c_bypass_0_0_is_stationary,
  output     [15:0]   io_out_c_bypass_0_1_data,
  output              io_out_c_bypass_0_1_is_stationary,
  output     [15:0]   io_out_c_bypass_0_2_data,
  output              io_out_c_bypass_0_2_is_stationary,
  output     [15:0]   io_out_c_bypass_0_3_data,
  output              io_out_c_bypass_0_3_is_stationary,
  output     [15:0]   io_out_c_bypass_1_0_data,
  output              io_out_c_bypass_1_0_is_stationary,
  output     [15:0]   io_out_c_bypass_1_1_data,
  output              io_out_c_bypass_1_1_is_stationary,
  output     [15:0]   io_out_c_bypass_1_2_data,
  output              io_out_c_bypass_1_2_is_stationary,
  output     [15:0]   io_out_c_bypass_1_3_data,
  output              io_out_c_bypass_1_3_is_stationary,
  output              io_out_c_input_from_bypass_0,
  output              io_out_c_input_from_bypass_1,
  input               clk,
  input               reset
);

  wire       [15:0]   pes_0_0_io_out_r_data;
  wire                pes_0_0_io_out_r_load_store;
  wire                pes_0_0_io_out_r_df_is_ws;
  wire                pes_0_0_io_out_r_stall;
  wire       [15:0]   pes_0_0_io_out_c_data;
  wire                pes_0_0_io_out_c_is_stationary;
  wire       [15:0]   pes_0_1_io_out_r_data;
  wire                pes_0_1_io_out_r_load_store;
  wire                pes_0_1_io_out_r_df_is_ws;
  wire                pes_0_1_io_out_r_stall;
  wire       [15:0]   pes_0_1_io_out_c_data;
  wire                pes_0_1_io_out_c_is_stationary;
  wire       [15:0]   pes_0_2_io_out_r_data;
  wire                pes_0_2_io_out_r_load_store;
  wire                pes_0_2_io_out_r_df_is_ws;
  wire                pes_0_2_io_out_r_stall;
  wire       [15:0]   pes_0_2_io_out_c_data;
  wire                pes_0_2_io_out_c_is_stationary;
  wire       [15:0]   pes_0_3_io_out_r_data;
  wire                pes_0_3_io_out_r_load_store;
  wire                pes_0_3_io_out_r_df_is_ws;
  wire                pes_0_3_io_out_r_stall;
  wire       [15:0]   pes_0_3_io_out_c_data;
  wire                pes_0_3_io_out_c_is_stationary;
  wire       [15:0]   pes_1_0_io_out_r_data;
  wire                pes_1_0_io_out_r_load_store;
  wire                pes_1_0_io_out_r_df_is_ws;
  wire                pes_1_0_io_out_r_stall;
  wire       [15:0]   pes_1_0_io_out_c_data;
  wire                pes_1_0_io_out_c_is_stationary;
  wire       [15:0]   pes_1_1_io_out_r_data;
  wire                pes_1_1_io_out_r_load_store;
  wire                pes_1_1_io_out_r_df_is_ws;
  wire                pes_1_1_io_out_r_stall;
  wire       [15:0]   pes_1_1_io_out_c_data;
  wire                pes_1_1_io_out_c_is_stationary;
  wire       [15:0]   pes_1_2_io_out_r_data;
  wire                pes_1_2_io_out_r_load_store;
  wire                pes_1_2_io_out_r_df_is_ws;
  wire                pes_1_2_io_out_r_stall;
  wire       [15:0]   pes_1_2_io_out_c_data;
  wire                pes_1_2_io_out_c_is_stationary;
  wire       [15:0]   pes_1_3_io_out_r_data;
  wire                pes_1_3_io_out_r_load_store;
  wire                pes_1_3_io_out_r_df_is_ws;
  wire                pes_1_3_io_out_r_stall;
  wire       [15:0]   pes_1_3_io_out_c_data;
  wire                pes_1_3_io_out_c_is_stationary;
  wire       [15:0]   pes_2_0_io_out_r_data;
  wire                pes_2_0_io_out_r_load_store;
  wire                pes_2_0_io_out_r_df_is_ws;
  wire                pes_2_0_io_out_r_stall;
  wire       [15:0]   pes_2_0_io_out_c_data;
  wire                pes_2_0_io_out_c_is_stationary;
  wire       [15:0]   pes_2_1_io_out_r_data;
  wire                pes_2_1_io_out_r_load_store;
  wire                pes_2_1_io_out_r_df_is_ws;
  wire                pes_2_1_io_out_r_stall;
  wire       [15:0]   pes_2_1_io_out_c_data;
  wire                pes_2_1_io_out_c_is_stationary;
  wire       [15:0]   pes_2_2_io_out_r_data;
  wire                pes_2_2_io_out_r_load_store;
  wire                pes_2_2_io_out_r_df_is_ws;
  wire                pes_2_2_io_out_r_stall;
  wire       [15:0]   pes_2_2_io_out_c_data;
  wire                pes_2_2_io_out_c_is_stationary;
  wire       [15:0]   pes_2_3_io_out_r_data;
  wire                pes_2_3_io_out_r_load_store;
  wire                pes_2_3_io_out_r_df_is_ws;
  wire                pes_2_3_io_out_r_stall;
  wire       [15:0]   pes_2_3_io_out_c_data;
  wire                pes_2_3_io_out_c_is_stationary;
  wire       [15:0]   pes_3_0_io_out_r_data;
  wire                pes_3_0_io_out_r_load_store;
  wire                pes_3_0_io_out_r_df_is_ws;
  wire                pes_3_0_io_out_r_stall;
  wire       [15:0]   pes_3_0_io_out_c_data;
  wire                pes_3_0_io_out_c_is_stationary;
  wire       [15:0]   pes_3_1_io_out_r_data;
  wire                pes_3_1_io_out_r_load_store;
  wire                pes_3_1_io_out_r_df_is_ws;
  wire                pes_3_1_io_out_r_stall;
  wire       [15:0]   pes_3_1_io_out_c_data;
  wire                pes_3_1_io_out_c_is_stationary;
  wire       [15:0]   pes_3_2_io_out_r_data;
  wire                pes_3_2_io_out_r_load_store;
  wire                pes_3_2_io_out_r_df_is_ws;
  wire                pes_3_2_io_out_r_stall;
  wire       [15:0]   pes_3_2_io_out_c_data;
  wire                pes_3_2_io_out_c_is_stationary;
  wire       [15:0]   pes_3_3_io_out_r_data;
  wire                pes_3_3_io_out_r_load_store;
  wire                pes_3_3_io_out_r_df_is_ws;
  wire                pes_3_3_io_out_r_stall;
  wire       [15:0]   pes_3_3_io_out_c_data;
  wire                pes_3_3_io_out_c_is_stationary;
  wire       [15:0]   in_r_0_data;
  wire                in_r_0_load_store;
  wire                in_r_0_df_is_ws;
  wire                in_r_0_stall;
  wire       [15:0]   in_r_1_data;
  wire                in_r_1_load_store;
  wire                in_r_1_df_is_ws;
  wire                in_r_1_stall;
  wire       [15:0]   in_r_2_data;
  wire                in_r_2_load_store;
  wire                in_r_2_df_is_ws;
  wire                in_r_2_stall;
  wire       [15:0]   in_r_3_data;
  wire                in_r_3_load_store;
  wire                in_r_3_df_is_ws;
  wire                in_r_3_stall;
  wire       [15:0]   in_c_0_data;
  wire                in_c_0_is_stationary;
  wire       [15:0]   in_c_1_data;
  wire                in_c_1_is_stationary;
  wire       [15:0]   in_c_2_data;
  wire                in_c_2_is_stationary;
  wire       [15:0]   in_c_3_data;
  wire                in_c_3_is_stationary;
  wire       [15:0]   out_r_0_data;
  wire                out_r_0_load_store;
  wire                out_r_0_df_is_ws;
  wire                out_r_0_stall;
  wire       [15:0]   out_r_1_data;
  wire                out_r_1_load_store;
  wire                out_r_1_df_is_ws;
  wire                out_r_1_stall;
  wire       [15:0]   out_r_2_data;
  wire                out_r_2_load_store;
  wire                out_r_2_df_is_ws;
  wire                out_r_2_stall;
  wire       [15:0]   out_r_3_data;
  wire                out_r_3_load_store;
  wire                out_r_3_df_is_ws;
  wire                out_r_3_stall;
  wire       [15:0]   out_c_0_data;
  wire                out_c_0_is_stationary;
  wire       [15:0]   out_c_1_data;
  wire                out_c_1_is_stationary;
  wire       [15:0]   out_c_2_data;
  wire                out_c_2_is_stationary;
  wire       [15:0]   out_c_3_data;
  wire                out_c_3_is_stationary;
  reg        [15:0]   out_r_regNext_0_data;
  reg                 out_r_regNext_0_load_store;
  reg                 out_r_regNext_0_df_is_ws;
  reg                 out_r_regNext_0_stall;
  reg        [15:0]   out_r_regNext_1_data;
  reg                 out_r_regNext_1_load_store;
  reg                 out_r_regNext_1_df_is_ws;
  reg                 out_r_regNext_1_stall;
  reg        [15:0]   out_r_regNext_2_data;
  reg                 out_r_regNext_2_load_store;
  reg                 out_r_regNext_2_df_is_ws;
  reg                 out_r_regNext_2_stall;
  reg        [15:0]   out_r_regNext_3_data;
  reg                 out_r_regNext_3_load_store;
  reg                 out_r_regNext_3_df_is_ws;
  reg                 out_r_regNext_3_stall;
  reg        [15:0]   out_c_regNext_0_data;
  reg                 out_c_regNext_0_is_stationary;
  reg        [15:0]   out_c_regNext_1_data;
  reg                 out_c_regNext_1_is_stationary;
  reg        [15:0]   out_c_regNext_2_data;
  reg                 out_c_regNext_2_is_stationary;
  reg        [15:0]   out_c_regNext_3_data;
  reg                 out_c_regNext_3_is_stationary;
  reg        [15:0]   io_in_r_bypass_regNext_0_0_data;
  reg                 io_in_r_bypass_regNext_0_0_load_store;
  reg                 io_in_r_bypass_regNext_0_0_df_is_ws;
  reg                 io_in_r_bypass_regNext_0_0_stall;
  reg        [15:0]   io_in_r_bypass_regNext_0_1_data;
  reg                 io_in_r_bypass_regNext_0_1_load_store;
  reg                 io_in_r_bypass_regNext_0_1_df_is_ws;
  reg                 io_in_r_bypass_regNext_0_1_stall;
  reg        [15:0]   io_in_r_bypass_regNext_0_2_data;
  reg                 io_in_r_bypass_regNext_0_2_load_store;
  reg                 io_in_r_bypass_regNext_0_2_df_is_ws;
  reg                 io_in_r_bypass_regNext_0_2_stall;
  reg        [15:0]   io_in_r_bypass_regNext_0_3_data;
  reg                 io_in_r_bypass_regNext_0_3_load_store;
  reg                 io_in_r_bypass_regNext_0_3_df_is_ws;
  reg                 io_in_r_bypass_regNext_0_3_stall;
  reg        [15:0]   io_in_r_bypass_regNext_1_0_data;
  reg                 io_in_r_bypass_regNext_1_0_load_store;
  reg                 io_in_r_bypass_regNext_1_0_df_is_ws;
  reg                 io_in_r_bypass_regNext_1_0_stall;
  reg        [15:0]   io_in_r_bypass_regNext_1_1_data;
  reg                 io_in_r_bypass_regNext_1_1_load_store;
  reg                 io_in_r_bypass_regNext_1_1_df_is_ws;
  reg                 io_in_r_bypass_regNext_1_1_stall;
  reg        [15:0]   io_in_r_bypass_regNext_1_2_data;
  reg                 io_in_r_bypass_regNext_1_2_load_store;
  reg                 io_in_r_bypass_regNext_1_2_df_is_ws;
  reg                 io_in_r_bypass_regNext_1_2_stall;
  reg        [15:0]   io_in_r_bypass_regNext_1_3_data;
  reg                 io_in_r_bypass_regNext_1_3_load_store;
  reg                 io_in_r_bypass_regNext_1_3_df_is_ws;
  reg                 io_in_r_bypass_regNext_1_3_stall;
  reg        [15:0]   io_in_c_bypass_regNext_0_0_data;
  reg                 io_in_c_bypass_regNext_0_0_is_stationary;
  reg        [15:0]   io_in_c_bypass_regNext_0_1_data;
  reg                 io_in_c_bypass_regNext_0_1_is_stationary;
  reg        [15:0]   io_in_c_bypass_regNext_0_2_data;
  reg                 io_in_c_bypass_regNext_0_2_is_stationary;
  reg        [15:0]   io_in_c_bypass_regNext_0_3_data;
  reg                 io_in_c_bypass_regNext_0_3_is_stationary;
  reg        [15:0]   io_in_c_bypass_regNext_1_0_data;
  reg                 io_in_c_bypass_regNext_1_0_is_stationary;
  reg        [15:0]   io_in_c_bypass_regNext_1_1_data;
  reg                 io_in_c_bypass_regNext_1_1_is_stationary;
  reg        [15:0]   io_in_c_bypass_regNext_1_2_data;
  reg                 io_in_c_bypass_regNext_1_2_is_stationary;
  reg        [15:0]   io_in_c_bypass_regNext_1_3_data;
  reg                 io_in_c_bypass_regNext_1_3_is_stationary;
  reg                 io_in_r_input_from_bypass_regNext_0;
  reg                 io_in_r_input_from_bypass_regNext_1;
  reg                 io_in_c_input_from_bypass_regNext_0;
  reg                 io_in_c_input_from_bypass_regNext_1;

  PEWSOS_127 pes_0_0 (
    .io_in_r_data           (in_r_0_data[15:0]             ), //i
    .io_in_r_load_store     (in_r_0_load_store             ), //i
    .io_in_r_df_is_ws       (in_r_0_df_is_ws               ), //i
    .io_in_r_stall          (in_r_0_stall                  ), //i
    .io_out_r_data          (pes_0_0_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pes_0_0_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pes_0_0_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pes_0_0_io_out_r_stall        ), //o
    .io_in_c_data           (in_c_0_data[15:0]             ), //i
    .io_in_c_is_stationary  (in_c_0_is_stationary          ), //i
    .io_out_c_data          (pes_0_0_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pes_0_0_io_out_c_is_stationary), //o
    .clk                    (clk                           ), //i
    .reset                  (reset                         )  //i
  );
  PEWSOS_127 pes_0_1 (
    .io_in_r_data           (pes_0_0_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pes_0_0_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pes_0_0_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pes_0_0_io_out_r_stall        ), //i
    .io_out_r_data          (pes_0_1_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pes_0_1_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pes_0_1_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pes_0_1_io_out_r_stall        ), //o
    .io_in_c_data           (in_c_1_data[15:0]             ), //i
    .io_in_c_is_stationary  (in_c_1_is_stationary          ), //i
    .io_out_c_data          (pes_0_1_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pes_0_1_io_out_c_is_stationary), //o
    .clk                    (clk                           ), //i
    .reset                  (reset                         )  //i
  );
  PEWSOS_127 pes_0_2 (
    .io_in_r_data           (pes_0_1_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pes_0_1_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pes_0_1_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pes_0_1_io_out_r_stall        ), //i
    .io_out_r_data          (pes_0_2_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pes_0_2_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pes_0_2_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pes_0_2_io_out_r_stall        ), //o
    .io_in_c_data           (in_c_2_data[15:0]             ), //i
    .io_in_c_is_stationary  (in_c_2_is_stationary          ), //i
    .io_out_c_data          (pes_0_2_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pes_0_2_io_out_c_is_stationary), //o
    .clk                    (clk                           ), //i
    .reset                  (reset                         )  //i
  );
  PEWSOS_127 pes_0_3 (
    .io_in_r_data           (pes_0_2_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pes_0_2_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pes_0_2_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pes_0_2_io_out_r_stall        ), //i
    .io_out_r_data          (pes_0_3_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pes_0_3_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pes_0_3_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pes_0_3_io_out_r_stall        ), //o
    .io_in_c_data           (in_c_3_data[15:0]             ), //i
    .io_in_c_is_stationary  (in_c_3_is_stationary          ), //i
    .io_out_c_data          (pes_0_3_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pes_0_3_io_out_c_is_stationary), //o
    .clk                    (clk                           ), //i
    .reset                  (reset                         )  //i
  );
  PEWSOS_127 pes_1_0 (
    .io_in_r_data           (in_r_1_data[15:0]             ), //i
    .io_in_r_load_store     (in_r_1_load_store             ), //i
    .io_in_r_df_is_ws       (in_r_1_df_is_ws               ), //i
    .io_in_r_stall          (in_r_1_stall                  ), //i
    .io_out_r_data          (pes_1_0_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pes_1_0_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pes_1_0_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pes_1_0_io_out_r_stall        ), //o
    .io_in_c_data           (pes_0_0_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pes_0_0_io_out_c_is_stationary), //i
    .io_out_c_data          (pes_1_0_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pes_1_0_io_out_c_is_stationary), //o
    .clk                    (clk                           ), //i
    .reset                  (reset                         )  //i
  );
  PEWSOS_127 pes_1_1 (
    .io_in_r_data           (pes_1_0_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pes_1_0_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pes_1_0_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pes_1_0_io_out_r_stall        ), //i
    .io_out_r_data          (pes_1_1_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pes_1_1_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pes_1_1_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pes_1_1_io_out_r_stall        ), //o
    .io_in_c_data           (pes_0_1_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pes_0_1_io_out_c_is_stationary), //i
    .io_out_c_data          (pes_1_1_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pes_1_1_io_out_c_is_stationary), //o
    .clk                    (clk                           ), //i
    .reset                  (reset                         )  //i
  );
  PEWSOS_127 pes_1_2 (
    .io_in_r_data           (pes_1_1_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pes_1_1_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pes_1_1_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pes_1_1_io_out_r_stall        ), //i
    .io_out_r_data          (pes_1_2_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pes_1_2_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pes_1_2_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pes_1_2_io_out_r_stall        ), //o
    .io_in_c_data           (pes_0_2_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pes_0_2_io_out_c_is_stationary), //i
    .io_out_c_data          (pes_1_2_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pes_1_2_io_out_c_is_stationary), //o
    .clk                    (clk                           ), //i
    .reset                  (reset                         )  //i
  );
  PEWSOS_127 pes_1_3 (
    .io_in_r_data           (pes_1_2_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pes_1_2_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pes_1_2_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pes_1_2_io_out_r_stall        ), //i
    .io_out_r_data          (pes_1_3_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pes_1_3_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pes_1_3_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pes_1_3_io_out_r_stall        ), //o
    .io_in_c_data           (pes_0_3_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pes_0_3_io_out_c_is_stationary), //i
    .io_out_c_data          (pes_1_3_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pes_1_3_io_out_c_is_stationary), //o
    .clk                    (clk                           ), //i
    .reset                  (reset                         )  //i
  );
  PEWSOS_127 pes_2_0 (
    .io_in_r_data           (in_r_2_data[15:0]             ), //i
    .io_in_r_load_store     (in_r_2_load_store             ), //i
    .io_in_r_df_is_ws       (in_r_2_df_is_ws               ), //i
    .io_in_r_stall          (in_r_2_stall                  ), //i
    .io_out_r_data          (pes_2_0_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pes_2_0_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pes_2_0_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pes_2_0_io_out_r_stall        ), //o
    .io_in_c_data           (pes_1_0_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pes_1_0_io_out_c_is_stationary), //i
    .io_out_c_data          (pes_2_0_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pes_2_0_io_out_c_is_stationary), //o
    .clk                    (clk                           ), //i
    .reset                  (reset                         )  //i
  );
  PEWSOS_127 pes_2_1 (
    .io_in_r_data           (pes_2_0_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pes_2_0_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pes_2_0_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pes_2_0_io_out_r_stall        ), //i
    .io_out_r_data          (pes_2_1_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pes_2_1_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pes_2_1_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pes_2_1_io_out_r_stall        ), //o
    .io_in_c_data           (pes_1_1_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pes_1_1_io_out_c_is_stationary), //i
    .io_out_c_data          (pes_2_1_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pes_2_1_io_out_c_is_stationary), //o
    .clk                    (clk                           ), //i
    .reset                  (reset                         )  //i
  );
  PEWSOS_127 pes_2_2 (
    .io_in_r_data           (pes_2_1_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pes_2_1_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pes_2_1_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pes_2_1_io_out_r_stall        ), //i
    .io_out_r_data          (pes_2_2_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pes_2_2_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pes_2_2_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pes_2_2_io_out_r_stall        ), //o
    .io_in_c_data           (pes_1_2_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pes_1_2_io_out_c_is_stationary), //i
    .io_out_c_data          (pes_2_2_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pes_2_2_io_out_c_is_stationary), //o
    .clk                    (clk                           ), //i
    .reset                  (reset                         )  //i
  );
  PEWSOS_127 pes_2_3 (
    .io_in_r_data           (pes_2_2_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pes_2_2_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pes_2_2_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pes_2_2_io_out_r_stall        ), //i
    .io_out_r_data          (pes_2_3_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pes_2_3_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pes_2_3_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pes_2_3_io_out_r_stall        ), //o
    .io_in_c_data           (pes_1_3_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pes_1_3_io_out_c_is_stationary), //i
    .io_out_c_data          (pes_2_3_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pes_2_3_io_out_c_is_stationary), //o
    .clk                    (clk                           ), //i
    .reset                  (reset                         )  //i
  );
  PEWSOS_127 pes_3_0 (
    .io_in_r_data           (in_r_3_data[15:0]             ), //i
    .io_in_r_load_store     (in_r_3_load_store             ), //i
    .io_in_r_df_is_ws       (in_r_3_df_is_ws               ), //i
    .io_in_r_stall          (in_r_3_stall                  ), //i
    .io_out_r_data          (pes_3_0_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pes_3_0_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pes_3_0_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pes_3_0_io_out_r_stall        ), //o
    .io_in_c_data           (pes_2_0_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pes_2_0_io_out_c_is_stationary), //i
    .io_out_c_data          (pes_3_0_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pes_3_0_io_out_c_is_stationary), //o
    .clk                    (clk                           ), //i
    .reset                  (reset                         )  //i
  );
  PEWSOS_127 pes_3_1 (
    .io_in_r_data           (pes_3_0_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pes_3_0_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pes_3_0_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pes_3_0_io_out_r_stall        ), //i
    .io_out_r_data          (pes_3_1_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pes_3_1_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pes_3_1_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pes_3_1_io_out_r_stall        ), //o
    .io_in_c_data           (pes_2_1_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pes_2_1_io_out_c_is_stationary), //i
    .io_out_c_data          (pes_3_1_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pes_3_1_io_out_c_is_stationary), //o
    .clk                    (clk                           ), //i
    .reset                  (reset                         )  //i
  );
  PEWSOS_127 pes_3_2 (
    .io_in_r_data           (pes_3_1_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pes_3_1_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pes_3_1_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pes_3_1_io_out_r_stall        ), //i
    .io_out_r_data          (pes_3_2_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pes_3_2_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pes_3_2_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pes_3_2_io_out_r_stall        ), //o
    .io_in_c_data           (pes_2_2_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pes_2_2_io_out_c_is_stationary), //i
    .io_out_c_data          (pes_3_2_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pes_3_2_io_out_c_is_stationary), //o
    .clk                    (clk                           ), //i
    .reset                  (reset                         )  //i
  );
  PEWSOS_127 pes_3_3 (
    .io_in_r_data           (pes_3_2_io_out_r_data[15:0]   ), //i
    .io_in_r_load_store     (pes_3_2_io_out_r_load_store   ), //i
    .io_in_r_df_is_ws       (pes_3_2_io_out_r_df_is_ws     ), //i
    .io_in_r_stall          (pes_3_2_io_out_r_stall        ), //i
    .io_out_r_data          (pes_3_3_io_out_r_data[15:0]   ), //o
    .io_out_r_load_store    (pes_3_3_io_out_r_load_store   ), //o
    .io_out_r_df_is_ws      (pes_3_3_io_out_r_df_is_ws     ), //o
    .io_out_r_stall         (pes_3_3_io_out_r_stall        ), //o
    .io_in_c_data           (pes_2_3_io_out_c_data[15:0]   ), //i
    .io_in_c_is_stationary  (pes_2_3_io_out_c_is_stationary), //i
    .io_out_c_data          (pes_3_3_io_out_c_data[15:0]   ), //o
    .io_out_c_is_stationary (pes_3_3_io_out_c_is_stationary), //o
    .clk                    (clk                           ), //i
    .reset                  (reset                         )  //i
  );
  assign in_r_0_data = (io_in_r_input_from_bypass_0 ? io_in_r_bypass_0_0_data : io_in_r_data_0_data); // @[Expression.scala 1420:25]
  assign in_r_0_load_store = (io_in_r_input_from_bypass_0 ? io_in_r_bypass_0_0_load_store : io_in_r_data_0_load_store); // @[Expression.scala 1420:25]
  assign in_r_0_df_is_ws = (io_in_r_input_from_bypass_0 ? io_in_r_bypass_0_0_df_is_ws : io_in_r_data_0_df_is_ws); // @[Expression.scala 1420:25]
  assign in_r_0_stall = (io_in_r_input_from_bypass_0 ? io_in_r_bypass_0_0_stall : io_in_r_data_0_stall); // @[Expression.scala 1420:25]
  assign in_r_1_data = (io_in_r_input_from_bypass_0 ? io_in_r_bypass_0_1_data : io_in_r_data_1_data); // @[Expression.scala 1420:25]
  assign in_r_1_load_store = (io_in_r_input_from_bypass_0 ? io_in_r_bypass_0_1_load_store : io_in_r_data_1_load_store); // @[Expression.scala 1420:25]
  assign in_r_1_df_is_ws = (io_in_r_input_from_bypass_0 ? io_in_r_bypass_0_1_df_is_ws : io_in_r_data_1_df_is_ws); // @[Expression.scala 1420:25]
  assign in_r_1_stall = (io_in_r_input_from_bypass_0 ? io_in_r_bypass_0_1_stall : io_in_r_data_1_stall); // @[Expression.scala 1420:25]
  assign in_r_2_data = (io_in_r_input_from_bypass_0 ? io_in_r_bypass_0_2_data : io_in_r_data_2_data); // @[Expression.scala 1420:25]
  assign in_r_2_load_store = (io_in_r_input_from_bypass_0 ? io_in_r_bypass_0_2_load_store : io_in_r_data_2_load_store); // @[Expression.scala 1420:25]
  assign in_r_2_df_is_ws = (io_in_r_input_from_bypass_0 ? io_in_r_bypass_0_2_df_is_ws : io_in_r_data_2_df_is_ws); // @[Expression.scala 1420:25]
  assign in_r_2_stall = (io_in_r_input_from_bypass_0 ? io_in_r_bypass_0_2_stall : io_in_r_data_2_stall); // @[Expression.scala 1420:25]
  assign in_r_3_data = (io_in_r_input_from_bypass_0 ? io_in_r_bypass_0_3_data : io_in_r_data_3_data); // @[Expression.scala 1420:25]
  assign in_r_3_load_store = (io_in_r_input_from_bypass_0 ? io_in_r_bypass_0_3_load_store : io_in_r_data_3_load_store); // @[Expression.scala 1420:25]
  assign in_r_3_df_is_ws = (io_in_r_input_from_bypass_0 ? io_in_r_bypass_0_3_df_is_ws : io_in_r_data_3_df_is_ws); // @[Expression.scala 1420:25]
  assign in_r_3_stall = (io_in_r_input_from_bypass_0 ? io_in_r_bypass_0_3_stall : io_in_r_data_3_stall); // @[Expression.scala 1420:25]
  assign in_c_0_data = (io_in_c_input_from_bypass_0 ? io_in_c_bypass_0_0_data : io_in_c_data_0_data); // @[Expression.scala 1420:25]
  assign in_c_0_is_stationary = (io_in_c_input_from_bypass_0 ? io_in_c_bypass_0_0_is_stationary : io_in_c_data_0_is_stationary); // @[Expression.scala 1420:25]
  assign in_c_1_data = (io_in_c_input_from_bypass_0 ? io_in_c_bypass_0_1_data : io_in_c_data_1_data); // @[Expression.scala 1420:25]
  assign in_c_1_is_stationary = (io_in_c_input_from_bypass_0 ? io_in_c_bypass_0_1_is_stationary : io_in_c_data_1_is_stationary); // @[Expression.scala 1420:25]
  assign in_c_2_data = (io_in_c_input_from_bypass_0 ? io_in_c_bypass_0_2_data : io_in_c_data_2_data); // @[Expression.scala 1420:25]
  assign in_c_2_is_stationary = (io_in_c_input_from_bypass_0 ? io_in_c_bypass_0_2_is_stationary : io_in_c_data_2_is_stationary); // @[Expression.scala 1420:25]
  assign in_c_3_data = (io_in_c_input_from_bypass_0 ? io_in_c_bypass_0_3_data : io_in_c_data_3_data); // @[Expression.scala 1420:25]
  assign in_c_3_is_stationary = (io_in_c_input_from_bypass_0 ? io_in_c_bypass_0_3_is_stationary : io_in_c_data_3_is_stationary); // @[Expression.scala 1420:25]
  assign out_r_0_data = pes_0_3_io_out_r_data; // @[SystolicConnect.scala 50:16]
  assign out_r_0_load_store = pes_0_3_io_out_r_load_store; // @[SystolicConnect.scala 50:16]
  assign out_r_0_df_is_ws = pes_0_3_io_out_r_df_is_ws; // @[SystolicConnect.scala 50:16]
  assign out_r_0_stall = pes_0_3_io_out_r_stall; // @[SystolicConnect.scala 50:16]
  assign out_r_1_data = pes_1_3_io_out_r_data; // @[SystolicConnect.scala 50:16]
  assign out_r_1_load_store = pes_1_3_io_out_r_load_store; // @[SystolicConnect.scala 50:16]
  assign out_r_1_df_is_ws = pes_1_3_io_out_r_df_is_ws; // @[SystolicConnect.scala 50:16]
  assign out_r_1_stall = pes_1_3_io_out_r_stall; // @[SystolicConnect.scala 50:16]
  assign out_r_2_data = pes_2_3_io_out_r_data; // @[SystolicConnect.scala 50:16]
  assign out_r_2_load_store = pes_2_3_io_out_r_load_store; // @[SystolicConnect.scala 50:16]
  assign out_r_2_df_is_ws = pes_2_3_io_out_r_df_is_ws; // @[SystolicConnect.scala 50:16]
  assign out_r_2_stall = pes_2_3_io_out_r_stall; // @[SystolicConnect.scala 50:16]
  assign out_r_3_data = pes_3_3_io_out_r_data; // @[SystolicConnect.scala 50:16]
  assign out_r_3_load_store = pes_3_3_io_out_r_load_store; // @[SystolicConnect.scala 50:16]
  assign out_r_3_df_is_ws = pes_3_3_io_out_r_df_is_ws; // @[SystolicConnect.scala 50:16]
  assign out_r_3_stall = pes_3_3_io_out_r_stall; // @[SystolicConnect.scala 50:16]
  assign out_c_0_data = pes_3_0_io_out_c_data; // @[SystolicConnect.scala 56:16]
  assign out_c_0_is_stationary = pes_3_0_io_out_c_is_stationary; // @[SystolicConnect.scala 56:16]
  assign out_c_1_data = pes_3_1_io_out_c_data; // @[SystolicConnect.scala 56:16]
  assign out_c_1_is_stationary = pes_3_1_io_out_c_is_stationary; // @[SystolicConnect.scala 56:16]
  assign out_c_2_data = pes_3_2_io_out_c_data; // @[SystolicConnect.scala 56:16]
  assign out_c_2_is_stationary = pes_3_2_io_out_c_is_stationary; // @[SystolicConnect.scala 56:16]
  assign out_c_3_data = pes_3_3_io_out_c_data; // @[SystolicConnect.scala 56:16]
  assign out_c_3_is_stationary = pes_3_3_io_out_c_is_stationary; // @[SystolicConnect.scala 56:16]
  assign io_out_r_data_0_data = out_r_0_data; // @[ArraySARA.scala 90:17]
  assign io_out_r_data_0_load_store = out_r_0_load_store; // @[ArraySARA.scala 90:17]
  assign io_out_r_data_0_df_is_ws = out_r_0_df_is_ws; // @[ArraySARA.scala 90:17]
  assign io_out_r_data_0_stall = out_r_0_stall; // @[ArraySARA.scala 90:17]
  assign io_out_r_data_1_data = out_r_1_data; // @[ArraySARA.scala 90:17]
  assign io_out_r_data_1_load_store = out_r_1_load_store; // @[ArraySARA.scala 90:17]
  assign io_out_r_data_1_df_is_ws = out_r_1_df_is_ws; // @[ArraySARA.scala 90:17]
  assign io_out_r_data_1_stall = out_r_1_stall; // @[ArraySARA.scala 90:17]
  assign io_out_r_data_2_data = out_r_2_data; // @[ArraySARA.scala 90:17]
  assign io_out_r_data_2_load_store = out_r_2_load_store; // @[ArraySARA.scala 90:17]
  assign io_out_r_data_2_df_is_ws = out_r_2_df_is_ws; // @[ArraySARA.scala 90:17]
  assign io_out_r_data_2_stall = out_r_2_stall; // @[ArraySARA.scala 90:17]
  assign io_out_r_data_3_data = out_r_3_data; // @[ArraySARA.scala 90:17]
  assign io_out_r_data_3_load_store = out_r_3_load_store; // @[ArraySARA.scala 90:17]
  assign io_out_r_data_3_df_is_ws = out_r_3_df_is_ws; // @[ArraySARA.scala 90:17]
  assign io_out_r_data_3_stall = out_r_3_stall; // @[ArraySARA.scala 90:17]
  assign io_out_c_data_0_data = out_c_0_data; // @[ArraySARA.scala 91:17]
  assign io_out_c_data_0_is_stationary = out_c_0_is_stationary; // @[ArraySARA.scala 91:17]
  assign io_out_c_data_1_data = out_c_1_data; // @[ArraySARA.scala 91:17]
  assign io_out_c_data_1_is_stationary = out_c_1_is_stationary; // @[ArraySARA.scala 91:17]
  assign io_out_c_data_2_data = out_c_2_data; // @[ArraySARA.scala 91:17]
  assign io_out_c_data_2_is_stationary = out_c_2_is_stationary; // @[ArraySARA.scala 91:17]
  assign io_out_c_data_3_data = out_c_3_data; // @[ArraySARA.scala 91:17]
  assign io_out_c_data_3_is_stationary = out_c_3_is_stationary; // @[ArraySARA.scala 91:17]
  assign io_out_r_bypass_0_0_data = out_r_regNext_0_data; // @[ArraySARA.scala 92:31]
  assign io_out_r_bypass_0_0_load_store = out_r_regNext_0_load_store; // @[ArraySARA.scala 92:31]
  assign io_out_r_bypass_0_0_df_is_ws = out_r_regNext_0_df_is_ws; // @[ArraySARA.scala 92:31]
  assign io_out_r_bypass_0_0_stall = out_r_regNext_0_stall; // @[ArraySARA.scala 92:31]
  assign io_out_r_bypass_0_1_data = out_r_regNext_1_data; // @[ArraySARA.scala 92:31]
  assign io_out_r_bypass_0_1_load_store = out_r_regNext_1_load_store; // @[ArraySARA.scala 92:31]
  assign io_out_r_bypass_0_1_df_is_ws = out_r_regNext_1_df_is_ws; // @[ArraySARA.scala 92:31]
  assign io_out_r_bypass_0_1_stall = out_r_regNext_1_stall; // @[ArraySARA.scala 92:31]
  assign io_out_r_bypass_0_2_data = out_r_regNext_2_data; // @[ArraySARA.scala 92:31]
  assign io_out_r_bypass_0_2_load_store = out_r_regNext_2_load_store; // @[ArraySARA.scala 92:31]
  assign io_out_r_bypass_0_2_df_is_ws = out_r_regNext_2_df_is_ws; // @[ArraySARA.scala 92:31]
  assign io_out_r_bypass_0_2_stall = out_r_regNext_2_stall; // @[ArraySARA.scala 92:31]
  assign io_out_r_bypass_0_3_data = out_r_regNext_3_data; // @[ArraySARA.scala 92:31]
  assign io_out_r_bypass_0_3_load_store = out_r_regNext_3_load_store; // @[ArraySARA.scala 92:31]
  assign io_out_r_bypass_0_3_df_is_ws = out_r_regNext_3_df_is_ws; // @[ArraySARA.scala 92:31]
  assign io_out_r_bypass_0_3_stall = out_r_regNext_3_stall; // @[ArraySARA.scala 92:31]
  assign io_out_c_bypass_0_0_data = out_c_regNext_0_data; // @[ArraySARA.scala 93:31]
  assign io_out_c_bypass_0_0_is_stationary = out_c_regNext_0_is_stationary; // @[ArraySARA.scala 93:31]
  assign io_out_c_bypass_0_1_data = out_c_regNext_1_data; // @[ArraySARA.scala 93:31]
  assign io_out_c_bypass_0_1_is_stationary = out_c_regNext_1_is_stationary; // @[ArraySARA.scala 93:31]
  assign io_out_c_bypass_0_2_data = out_c_regNext_2_data; // @[ArraySARA.scala 93:31]
  assign io_out_c_bypass_0_2_is_stationary = out_c_regNext_2_is_stationary; // @[ArraySARA.scala 93:31]
  assign io_out_c_bypass_0_3_data = out_c_regNext_3_data; // @[ArraySARA.scala 93:31]
  assign io_out_c_bypass_0_3_is_stationary = out_c_regNext_3_is_stationary; // @[ArraySARA.scala 93:31]
  assign io_out_r_bypass_1_0_data = io_in_r_bypass_regNext_1_0_data; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_1_0_load_store = io_in_r_bypass_regNext_1_0_load_store; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_1_0_df_is_ws = io_in_r_bypass_regNext_1_0_df_is_ws; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_1_0_stall = io_in_r_bypass_regNext_1_0_stall; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_1_1_data = io_in_r_bypass_regNext_1_1_data; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_1_1_load_store = io_in_r_bypass_regNext_1_1_load_store; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_1_1_df_is_ws = io_in_r_bypass_regNext_1_1_df_is_ws; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_1_1_stall = io_in_r_bypass_regNext_1_1_stall; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_1_2_data = io_in_r_bypass_regNext_1_2_data; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_1_2_load_store = io_in_r_bypass_regNext_1_2_load_store; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_1_2_df_is_ws = io_in_r_bypass_regNext_1_2_df_is_ws; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_1_2_stall = io_in_r_bypass_regNext_1_2_stall; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_1_3_data = io_in_r_bypass_regNext_1_3_data; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_1_3_load_store = io_in_r_bypass_regNext_1_3_load_store; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_1_3_df_is_ws = io_in_r_bypass_regNext_1_3_df_is_ws; // @[ArraySARA.scala 97:26]
  assign io_out_r_bypass_1_3_stall = io_in_r_bypass_regNext_1_3_stall; // @[ArraySARA.scala 97:26]
  assign io_out_c_bypass_1_0_data = io_in_c_bypass_regNext_1_0_data; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_1_0_is_stationary = io_in_c_bypass_regNext_1_0_is_stationary; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_1_1_data = io_in_c_bypass_regNext_1_1_data; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_1_1_is_stationary = io_in_c_bypass_regNext_1_1_is_stationary; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_1_2_data = io_in_c_bypass_regNext_1_2_data; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_1_2_is_stationary = io_in_c_bypass_regNext_1_2_is_stationary; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_1_3_data = io_in_c_bypass_regNext_1_3_data; // @[ArraySARA.scala 101:26]
  assign io_out_c_bypass_1_3_is_stationary = io_in_c_bypass_regNext_1_3_is_stationary; // @[ArraySARA.scala 101:26]
  assign io_out_r_input_from_bypass_0 = io_in_r_input_from_bypass_regNext_0; // @[ArraySARA.scala 103:30]
  assign io_out_r_input_from_bypass_1 = io_in_r_input_from_bypass_regNext_1; // @[ArraySARA.scala 103:30]
  assign io_out_c_input_from_bypass_0 = io_in_c_input_from_bypass_regNext_0; // @[ArraySARA.scala 104:30]
  assign io_out_c_input_from_bypass_1 = io_in_c_input_from_bypass_regNext_1; // @[ArraySARA.scala 104:30]
  always @(posedge clk) begin
    out_r_regNext_0_data <= out_r_0_data; // @[Reg.scala 39:30]
    out_r_regNext_0_load_store <= out_r_0_load_store; // @[Reg.scala 39:30]
    out_r_regNext_0_df_is_ws <= out_r_0_df_is_ws; // @[Reg.scala 39:30]
    out_r_regNext_0_stall <= out_r_0_stall; // @[Reg.scala 39:30]
    out_r_regNext_1_data <= out_r_1_data; // @[Reg.scala 39:30]
    out_r_regNext_1_load_store <= out_r_1_load_store; // @[Reg.scala 39:30]
    out_r_regNext_1_df_is_ws <= out_r_1_df_is_ws; // @[Reg.scala 39:30]
    out_r_regNext_1_stall <= out_r_1_stall; // @[Reg.scala 39:30]
    out_r_regNext_2_data <= out_r_2_data; // @[Reg.scala 39:30]
    out_r_regNext_2_load_store <= out_r_2_load_store; // @[Reg.scala 39:30]
    out_r_regNext_2_df_is_ws <= out_r_2_df_is_ws; // @[Reg.scala 39:30]
    out_r_regNext_2_stall <= out_r_2_stall; // @[Reg.scala 39:30]
    out_r_regNext_3_data <= out_r_3_data; // @[Reg.scala 39:30]
    out_r_regNext_3_load_store <= out_r_3_load_store; // @[Reg.scala 39:30]
    out_r_regNext_3_df_is_ws <= out_r_3_df_is_ws; // @[Reg.scala 39:30]
    out_r_regNext_3_stall <= out_r_3_stall; // @[Reg.scala 39:30]
    out_c_regNext_0_data <= out_c_0_data; // @[Reg.scala 39:30]
    out_c_regNext_0_is_stationary <= out_c_0_is_stationary; // @[Reg.scala 39:30]
    out_c_regNext_1_data <= out_c_1_data; // @[Reg.scala 39:30]
    out_c_regNext_1_is_stationary <= out_c_1_is_stationary; // @[Reg.scala 39:30]
    out_c_regNext_2_data <= out_c_2_data; // @[Reg.scala 39:30]
    out_c_regNext_2_is_stationary <= out_c_2_is_stationary; // @[Reg.scala 39:30]
    out_c_regNext_3_data <= out_c_3_data; // @[Reg.scala 39:30]
    out_c_regNext_3_is_stationary <= out_c_3_is_stationary; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_0_data <= io_in_r_bypass_0_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_0_load_store <= io_in_r_bypass_0_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_0_df_is_ws <= io_in_r_bypass_0_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_0_stall <= io_in_r_bypass_0_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_1_data <= io_in_r_bypass_0_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_1_load_store <= io_in_r_bypass_0_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_1_df_is_ws <= io_in_r_bypass_0_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_1_stall <= io_in_r_bypass_0_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_2_data <= io_in_r_bypass_0_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_2_load_store <= io_in_r_bypass_0_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_2_df_is_ws <= io_in_r_bypass_0_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_2_stall <= io_in_r_bypass_0_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_3_data <= io_in_r_bypass_0_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_3_load_store <= io_in_r_bypass_0_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_3_df_is_ws <= io_in_r_bypass_0_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_0_3_stall <= io_in_r_bypass_0_3_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_0_data <= io_in_r_bypass_1_0_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_0_load_store <= io_in_r_bypass_1_0_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_0_df_is_ws <= io_in_r_bypass_1_0_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_0_stall <= io_in_r_bypass_1_0_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_1_data <= io_in_r_bypass_1_1_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_1_load_store <= io_in_r_bypass_1_1_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_1_df_is_ws <= io_in_r_bypass_1_1_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_1_stall <= io_in_r_bypass_1_1_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_2_data <= io_in_r_bypass_1_2_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_2_load_store <= io_in_r_bypass_1_2_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_2_df_is_ws <= io_in_r_bypass_1_2_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_2_stall <= io_in_r_bypass_1_2_stall; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_3_data <= io_in_r_bypass_1_3_data; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_3_load_store <= io_in_r_bypass_1_3_load_store; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_3_df_is_ws <= io_in_r_bypass_1_3_df_is_ws; // @[Reg.scala 39:30]
    io_in_r_bypass_regNext_1_3_stall <= io_in_r_bypass_1_3_stall; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_0_data <= io_in_c_bypass_0_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_0_is_stationary <= io_in_c_bypass_0_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_1_data <= io_in_c_bypass_0_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_1_is_stationary <= io_in_c_bypass_0_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_2_data <= io_in_c_bypass_0_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_2_is_stationary <= io_in_c_bypass_0_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_3_data <= io_in_c_bypass_0_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_0_3_is_stationary <= io_in_c_bypass_0_3_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_0_data <= io_in_c_bypass_1_0_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_0_is_stationary <= io_in_c_bypass_1_0_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_1_data <= io_in_c_bypass_1_1_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_1_is_stationary <= io_in_c_bypass_1_1_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_2_data <= io_in_c_bypass_1_2_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_2_is_stationary <= io_in_c_bypass_1_2_is_stationary; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_3_data <= io_in_c_bypass_1_3_data; // @[Reg.scala 39:30]
    io_in_c_bypass_regNext_1_3_is_stationary <= io_in_c_bypass_1_3_is_stationary; // @[Reg.scala 39:30]
    io_in_r_input_from_bypass_regNext_0 <= io_in_r_input_from_bypass_0; // @[Reg.scala 39:30]
    io_in_r_input_from_bypass_regNext_1 <= io_in_r_input_from_bypass_1; // @[Reg.scala 39:30]
    io_in_c_input_from_bypass_regNext_0 <= io_in_c_input_from_bypass_0; // @[Reg.scala 39:30]
    io_in_c_input_from_bypass_regNext_1 <= io_in_c_input_from_bypass_1; // @[Reg.scala 39:30]
  end


endmodule

//PEWSOS_127 replaced by PEWSOS_127

//PEWSOS_127 replaced by PEWSOS_127

//PEWSOS_127 replaced by PEWSOS_127

//PEWSOS_127 replaced by PEWSOS_127

//PEWSOS_127 replaced by PEWSOS_127

//PEWSOS_127 replaced by PEWSOS_127

//PEWSOS_127 replaced by PEWSOS_127

//PEWSOS_127 replaced by PEWSOS_127

//PEWSOS_127 replaced by PEWSOS_127

//PEWSOS_127 replaced by PEWSOS_127

//PEWSOS_127 replaced by PEWSOS_127

//PEWSOS_127 replaced by PEWSOS_127

//PEWSOS_127 replaced by PEWSOS_127

//PEWSOS_127 replaced by PEWSOS_127

//PEWSOS_127 replaced by PEWSOS_127

//PEWSOS_127 replaced by PEWSOS_127

//PEWSOS_127 replaced by PEWSOS_127

//PEWSOS_127 replaced by PEWSOS_127

//PEWSOS_127 replaced by PEWSOS_127

//PEWSOS_127 replaced by PEWSOS_127

//PEWSOS_127 replaced by PEWSOS_127

//PEWSOS_127 replaced by PEWSOS_127

//PEWSOS_127 replaced by PEWSOS_127

//PEWSOS_127 replaced by PEWSOS_127

//PEWSOS_127 replaced by PEWSOS_127

//PEWSOS_127 replaced by PEWSOS_127

//PEWSOS_127 replaced by PEWSOS_127

//PEWSOS_127 replaced by PEWSOS_127

//PEWSOS_127 replaced by PEWSOS_127

//PEWSOS_127 replaced by PEWSOS_127

//PEWSOS_127 replaced by PEWSOS_127

//PEWSOS_127 replaced by PEWSOS_127

//PEWSOS_127 replaced by PEWSOS_127

//PEWSOS_127 replaced by PEWSOS_127

//PEWSOS_127 replaced by PEWSOS_127

//PEWSOS_127 replaced by PEWSOS_127

//PEWSOS_127 replaced by PEWSOS_127

//PEWSOS_127 replaced by PEWSOS_127

//PEWSOS_127 replaced by PEWSOS_127

//PEWSOS_127 replaced by PEWSOS_127

//PEWSOS_127 replaced by PEWSOS_127

//PEWSOS_127 replaced by PEWSOS_127

//PEWSOS_127 replaced by PEWSOS_127

//PEWSOS_127 replaced by PEWSOS_127

//PEWSOS_127 replaced by PEWSOS_127

//PEWSOS_127 replaced by PEWSOS_127

//PEWSOS_127 replaced by PEWSOS_127

//PEWSOS_127 replaced by PEWSOS_127

//PEWSOS_127 replaced by PEWSOS_127

//PEWSOS_127 replaced by PEWSOS_127

//PEWSOS_127 replaced by PEWSOS_127

//PEWSOS_127 replaced by PEWSOS_127

//PEWSOS_127 replaced by PEWSOS_127

//PEWSOS_127 replaced by PEWSOS_127

//PEWSOS_127 replaced by PEWSOS_127

//PEWSOS_127 replaced by PEWSOS_127

//PEWSOS_127 replaced by PEWSOS_127

//PEWSOS_127 replaced by PEWSOS_127

//PEWSOS_127 replaced by PEWSOS_127

//PEWSOS_127 replaced by PEWSOS_127

//PEWSOS_127 replaced by PEWSOS_127

//PEWSOS_127 replaced by PEWSOS_127

//PEWSOS_127 replaced by PEWSOS_127

//PEWSOS_127 replaced by PEWSOS_127

//PEWSOS_127 replaced by PEWSOS_127

//PEWSOS_127 replaced by PEWSOS_127

//PEWSOS_127 replaced by PEWSOS_127

//PEWSOS_127 replaced by PEWSOS_127

//PEWSOS_127 replaced by PEWSOS_127

//PEWSOS_127 replaced by PEWSOS_127

//PEWSOS_127 replaced by PEWSOS_127

//PEWSOS_127 replaced by PEWSOS_127

//PEWSOS_127 replaced by PEWSOS_127

//PEWSOS_127 replaced by PEWSOS_127

//PEWSOS_127 replaced by PEWSOS_127

//PEWSOS_127 replaced by PEWSOS_127

//PEWSOS_127 replaced by PEWSOS_127

//PEWSOS_127 replaced by PEWSOS_127

//PEWSOS_127 replaced by PEWSOS_127

//PEWSOS_127 replaced by PEWSOS_127

//PEWSOS_127 replaced by PEWSOS_127

//PEWSOS_127 replaced by PEWSOS_127

//PEWSOS_127 replaced by PEWSOS_127

//PEWSOS_127 replaced by PEWSOS_127

//PEWSOS_127 replaced by PEWSOS_127

//PEWSOS_127 replaced by PEWSOS_127

//PEWSOS_127 replaced by PEWSOS_127

//PEWSOS_127 replaced by PEWSOS_127

//PEWSOS_127 replaced by PEWSOS_127

//PEWSOS_127 replaced by PEWSOS_127

//PEWSOS_127 replaced by PEWSOS_127

//PEWSOS_127 replaced by PEWSOS_127

//PEWSOS_127 replaced by PEWSOS_127

//PEWSOS_127 replaced by PEWSOS_127

//PEWSOS_127 replaced by PEWSOS_127

//PEWSOS_127 replaced by PEWSOS_127

//PEWSOS_127 replaced by PEWSOS_127

//PEWSOS_127 replaced by PEWSOS_127

//PEWSOS_127 replaced by PEWSOS_127

//PEWSOS_127 replaced by PEWSOS_127

//PEWSOS_127 replaced by PEWSOS_127

//PEWSOS_127 replaced by PEWSOS_127

//PEWSOS_127 replaced by PEWSOS_127

//PEWSOS_127 replaced by PEWSOS_127

//PEWSOS_127 replaced by PEWSOS_127

//PEWSOS_127 replaced by PEWSOS_127

//PEWSOS_127 replaced by PEWSOS_127

//PEWSOS_127 replaced by PEWSOS_127

//PEWSOS_127 replaced by PEWSOS_127

//PEWSOS_127 replaced by PEWSOS_127

//PEWSOS_127 replaced by PEWSOS_127

//PEWSOS_127 replaced by PEWSOS_127

//PEWSOS_127 replaced by PEWSOS_127

//PEWSOS_127 replaced by PEWSOS_127

//PEWSOS_127 replaced by PEWSOS_127

//PEWSOS_127 replaced by PEWSOS_127

//PEWSOS_127 replaced by PEWSOS_127

//PEWSOS_127 replaced by PEWSOS_127

//PEWSOS_127 replaced by PEWSOS_127

//PEWSOS_127 replaced by PEWSOS_127

//PEWSOS_127 replaced by PEWSOS_127

//PEWSOS_127 replaced by PEWSOS_127

//PEWSOS_127 replaced by PEWSOS_127

//PEWSOS_127 replaced by PEWSOS_127

//PEWSOS_127 replaced by PEWSOS_127

//PEWSOS_127 replaced by PEWSOS_127

//PEWSOS_127 replaced by PEWSOS_127

module PEWSOS_127 (
  input      [15:0]   io_in_r_data,
  input               io_in_r_load_store,
  input               io_in_r_df_is_ws,
  input               io_in_r_stall,
  output     [15:0]   io_out_r_data,
  output              io_out_r_load_store,
  output              io_out_r_df_is_ws,
  output              io_out_r_stall,
  input      [15:0]   io_in_c_data,
  input               io_in_c_is_stationary,
  output     [15:0]   io_out_c_data,
  output              io_out_c_is_stationary,
  input               clk,
  input               reset
);

  wire       [15:0]   mac_128_io_psum;
  wire       [15:0]   mac_128_io_weight;
  wire       [15:0]   mac_128_io_result;
  wire                not_stall;
  wire       [15:0]   mac_result;
  reg        [15:0]   stationary;
  reg                 stationary_en;
  wire                when_PEWSOS_l68;
  reg        [15:0]   stationary_reg;
  reg                 io_in_r_stall_regNext;
  reg        [15:0]   io_in_r_data_regNextWhen;
  reg                 io_in_r_load_store_regNextWhen;
  reg                 io_in_r_df_is_ws_regNextWhen;
  reg        [15:0]   out_c_data;
  reg                 out_c_is_stationary;
  wire                when_PEWSOS_l87;
  wire                when_PEWSOS_l95;
  reg        [15:0]   out_c_data_regNextWhen;
  reg                 out_c_is_stationary_regNextWhen;

  Mac_127 mac_128 (
    .io_psum            (mac_128_io_psum[15:0]  ), //i
    .io_weight          (mac_128_io_weight[15:0]), //i
    .io_inputActivation (io_in_r_data[15:0]     ), //i
    .io_result          (mac_128_io_result[15:0])  //o
  );
  assign not_stall = (! io_in_r_stall); // @[BaseType.scala 299:24]
  always @(*) begin
    if(io_in_r_df_is_ws) begin
      stationary = io_in_c_data; // @[PEWSOS.scala 57:16]
    end else begin
      if(io_in_c_is_stationary) begin
        stationary = 16'h0; // @[PEWSOS.scala 61:18]
      end else begin
        stationary = mac_result; // @[PEWSOS.scala 64:18]
      end
    end
  end

  always @(*) begin
    if(io_in_r_df_is_ws) begin
      stationary_en = io_in_r_load_store; // @[PEWSOS.scala 58:19]
    end else begin
      if(io_in_c_is_stationary) begin
        stationary_en = io_in_r_load_store; // @[PEWSOS.scala 62:21]
      end else begin
        stationary_en = 1'b1; // @[PEWSOS.scala 65:21]
      end
    end
  end

  assign when_PEWSOS_l68 = (stationary_en && not_stall); // @[BaseType.scala 305:24]
  assign mac_128_io_psum = (io_in_r_df_is_ws ? io_in_c_data : stationary_reg); // @[PEWSOS.scala 72:15]
  assign mac_128_io_weight = (io_in_r_df_is_ws ? stationary_reg : io_in_c_data); // @[PEWSOS.scala 73:17]
  assign mac_result = mac_128_io_result; // @[PEWSOS.scala 75:14]
  assign io_out_r_stall = io_in_r_stall_regNext; // @[PEWSOS.scala 78:18]
  assign io_out_r_data = io_in_r_data_regNextWhen; // @[PEWSOS.scala 79:17]
  assign io_out_r_load_store = io_in_r_load_store_regNextWhen; // @[PEWSOS.scala 80:23]
  assign io_out_r_df_is_ws = io_in_r_df_is_ws_regNextWhen; // @[PEWSOS.scala 81:21]
  assign when_PEWSOS_l87 = (io_in_c_is_stationary && (! io_in_r_load_store)); // @[BaseType.scala 305:24]
  always @(*) begin
    if(io_in_r_df_is_ws) begin
      if(when_PEWSOS_l87) begin
        out_c_data = io_in_c_data; // @[PEWSOS.scala 88:18]
      end else begin
        out_c_data = mac_result; // @[PEWSOS.scala 91:18]
      end
    end else begin
      if(when_PEWSOS_l95) begin
        out_c_data = io_in_c_data; // @[PEWSOS.scala 96:18]
      end else begin
        if(io_in_r_load_store) begin
          out_c_data = stationary_reg; // @[PEWSOS.scala 99:18]
        end else begin
          out_c_data = io_in_c_data; // @[PEWSOS.scala 102:18]
        end
      end
    end
  end

  always @(*) begin
    if(io_in_r_df_is_ws) begin
      if(when_PEWSOS_l87) begin
        out_c_is_stationary = 1'b1; // @[PEWSOS.scala 89:27]
      end else begin
        out_c_is_stationary = 1'b0; // @[PEWSOS.scala 92:27]
      end
    end else begin
      if(when_PEWSOS_l95) begin
        out_c_is_stationary = 1'b1; // @[PEWSOS.scala 97:27]
      end else begin
        if(io_in_r_load_store) begin
          out_c_is_stationary = 1'b1; // @[PEWSOS.scala 100:27]
        end else begin
          out_c_is_stationary = 1'b0; // @[PEWSOS.scala 103:27]
        end
      end
    end
  end

  assign when_PEWSOS_l95 = (io_in_c_is_stationary && (! io_in_r_load_store)); // @[BaseType.scala 305:24]
  assign io_out_c_data = out_c_data_regNextWhen; // @[PEWSOS.scala 106:17]
  assign io_out_c_is_stationary = out_c_is_stationary_regNextWhen; // @[PEWSOS.scala 107:26]
  always @(posedge clk) begin
    if(when_PEWSOS_l68) begin
      stationary_reg <= stationary; // @[PEWSOS.scala 68:35]
    end
    io_in_r_stall_regNext <= io_in_r_stall; // @[Reg.scala 39:30]
    if(not_stall) begin
      io_in_r_data_regNextWhen <= io_in_r_data; // @[PEWSOS.scala 79:31]
    end
    if(not_stall) begin
      io_in_r_load_store_regNextWhen <= io_in_r_load_store; // @[PEWSOS.scala 80:37]
    end
    if(not_stall) begin
      io_in_r_df_is_ws_regNextWhen <= io_in_r_df_is_ws; // @[PEWSOS.scala 81:35]
    end
    if(not_stall) begin
      out_c_data_regNextWhen <= out_c_data; // @[PEWSOS.scala 106:31]
    end
    if(not_stall) begin
      out_c_is_stationary_regNextWhen <= out_c_is_stationary; // @[PEWSOS.scala 107:40]
    end
  end


endmodule

//Mac_127 replaced by Mac_127

//Mac_127 replaced by Mac_127

//Mac_127 replaced by Mac_127

//Mac_127 replaced by Mac_127

//Mac_127 replaced by Mac_127

//Mac_127 replaced by Mac_127

//Mac_127 replaced by Mac_127

//Mac_127 replaced by Mac_127

//Mac_127 replaced by Mac_127

//Mac_127 replaced by Mac_127

//Mac_127 replaced by Mac_127

//Mac_127 replaced by Mac_127

//Mac_127 replaced by Mac_127

//Mac_127 replaced by Mac_127

//Mac_127 replaced by Mac_127

//Mac_127 replaced by Mac_127

//Mac_127 replaced by Mac_127

//Mac_127 replaced by Mac_127

//Mac_127 replaced by Mac_127

//Mac_127 replaced by Mac_127

//Mac_127 replaced by Mac_127

//Mac_127 replaced by Mac_127

//Mac_127 replaced by Mac_127

//Mac_127 replaced by Mac_127

//Mac_127 replaced by Mac_127

//Mac_127 replaced by Mac_127

//Mac_127 replaced by Mac_127

//Mac_127 replaced by Mac_127

//Mac_127 replaced by Mac_127

//Mac_127 replaced by Mac_127

//Mac_127 replaced by Mac_127

//Mac_127 replaced by Mac_127

//Mac_127 replaced by Mac_127

//Mac_127 replaced by Mac_127

//Mac_127 replaced by Mac_127

//Mac_127 replaced by Mac_127

//Mac_127 replaced by Mac_127

//Mac_127 replaced by Mac_127

//Mac_127 replaced by Mac_127

//Mac_127 replaced by Mac_127

//Mac_127 replaced by Mac_127

//Mac_127 replaced by Mac_127

//Mac_127 replaced by Mac_127

//Mac_127 replaced by Mac_127

//Mac_127 replaced by Mac_127

//Mac_127 replaced by Mac_127

//Mac_127 replaced by Mac_127

//Mac_127 replaced by Mac_127

//Mac_127 replaced by Mac_127

//Mac_127 replaced by Mac_127

//Mac_127 replaced by Mac_127

//Mac_127 replaced by Mac_127

//Mac_127 replaced by Mac_127

//Mac_127 replaced by Mac_127

//Mac_127 replaced by Mac_127

//Mac_127 replaced by Mac_127

//Mac_127 replaced by Mac_127

//Mac_127 replaced by Mac_127

//Mac_127 replaced by Mac_127

//Mac_127 replaced by Mac_127

//Mac_127 replaced by Mac_127

//Mac_127 replaced by Mac_127

//Mac_127 replaced by Mac_127

//Mac_127 replaced by Mac_127

//Mac_127 replaced by Mac_127

//Mac_127 replaced by Mac_127

//Mac_127 replaced by Mac_127

//Mac_127 replaced by Mac_127

//Mac_127 replaced by Mac_127

//Mac_127 replaced by Mac_127

//Mac_127 replaced by Mac_127

//Mac_127 replaced by Mac_127

//Mac_127 replaced by Mac_127

//Mac_127 replaced by Mac_127

//Mac_127 replaced by Mac_127

//Mac_127 replaced by Mac_127

//Mac_127 replaced by Mac_127

//Mac_127 replaced by Mac_127

//Mac_127 replaced by Mac_127

//Mac_127 replaced by Mac_127

//Mac_127 replaced by Mac_127

//Mac_127 replaced by Mac_127

//Mac_127 replaced by Mac_127

//Mac_127 replaced by Mac_127

//Mac_127 replaced by Mac_127

//Mac_127 replaced by Mac_127

//Mac_127 replaced by Mac_127

//Mac_127 replaced by Mac_127

//Mac_127 replaced by Mac_127

//Mac_127 replaced by Mac_127

//Mac_127 replaced by Mac_127

//Mac_127 replaced by Mac_127

//Mac_127 replaced by Mac_127

//Mac_127 replaced by Mac_127

//Mac_127 replaced by Mac_127

//Mac_127 replaced by Mac_127

//Mac_127 replaced by Mac_127

//Mac_127 replaced by Mac_127

//Mac_127 replaced by Mac_127

//Mac_127 replaced by Mac_127

//Mac_127 replaced by Mac_127

//Mac_127 replaced by Mac_127

//Mac_127 replaced by Mac_127

//Mac_127 replaced by Mac_127

//Mac_127 replaced by Mac_127

//Mac_127 replaced by Mac_127

//Mac_127 replaced by Mac_127

//Mac_127 replaced by Mac_127

//Mac_127 replaced by Mac_127

//Mac_127 replaced by Mac_127

//Mac_127 replaced by Mac_127

//Mac_127 replaced by Mac_127

//Mac_127 replaced by Mac_127

//Mac_127 replaced by Mac_127

//Mac_127 replaced by Mac_127

//Mac_127 replaced by Mac_127

//Mac_127 replaced by Mac_127

//Mac_127 replaced by Mac_127

//Mac_127 replaced by Mac_127

//Mac_127 replaced by Mac_127

//Mac_127 replaced by Mac_127

//Mac_127 replaced by Mac_127

//Mac_127 replaced by Mac_127

//Mac_127 replaced by Mac_127

//Mac_127 replaced by Mac_127

//Mac_127 replaced by Mac_127

//Mac_127 replaced by Mac_127

module Mac_127 (
  input      [15:0]   io_psum,
  input      [15:0]   io_weight,
  input      [15:0]   io_inputActivation,
  output     [15:0]   io_result
);

  wire       [31:0]   _zz_io_result;
  wire       [31:0]   _zz_io_result_1;
  wire       [31:0]   _zz_io_result_2;

  assign _zz_io_result = ($signed(_zz_io_result_1) + $signed(_zz_io_result_2));
  assign _zz_io_result_1 = ($signed(io_inputActivation) * $signed(io_weight));
  assign _zz_io_result_2 = {{16{io_psum[15]}}, io_psum};
  assign io_result = _zz_io_result[15:0]; // @[Mac.scala 14:31]

endmodule
